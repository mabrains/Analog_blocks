magic
tech sky130A
magscale 1 2
timestamp 1624884095
<< checkpaint >>
rect -1245 -977 16357 6410
<< nwell >>
rect 415 600 14720 4720
<< pwell >>
rect 133 4857 14966 5109
rect 133 535 355 4857
rect 14780 535 14966 4857
rect 133 283 14966 535
<< mvpmos >>
rect 881 3152 1001 4152
rect 1311 3152 1431 4152
rect 1873 3152 1993 4152
rect 2303 3152 2423 4152
rect 2865 3152 2985 4152
rect 3295 3152 3415 4152
rect 3857 3152 3977 4152
rect 4287 3152 4407 4152
rect 4849 3152 4969 4152
rect 5279 3152 5399 4152
rect 5841 3152 5961 4152
rect 6271 3152 6391 4152
rect 6833 3152 6953 4152
rect 7263 3152 7383 4152
rect 7825 3152 7945 4152
rect 8255 3152 8375 4152
rect 8817 3152 8937 4152
rect 9247 3152 9367 4152
rect 9809 3152 9929 4152
rect 10239 3152 10359 4152
rect 10801 3152 10921 4152
rect 11231 3152 11351 4152
rect 11793 3152 11913 4152
rect 12223 3152 12343 4152
rect 12785 3152 12905 4152
rect 13215 3152 13335 4152
rect 13777 3152 13897 4152
rect 14135 3152 14255 4152
rect 881 1552 1001 2552
rect 1311 1552 1431 2552
rect 1873 1552 1993 2552
rect 2303 1552 2423 2552
rect 2865 1552 2985 2552
rect 3295 1552 3415 2552
rect 3857 1552 3977 2552
rect 4287 1552 4407 2552
rect 4849 1552 4969 2552
rect 5279 1552 5399 2552
rect 5841 1552 5961 2552
rect 6271 1552 6391 2552
rect 6833 1552 6953 2552
rect 7263 1552 7383 2552
rect 7825 1552 7945 2552
rect 8255 1552 8375 2552
rect 8817 1552 8937 2552
rect 9247 1552 9367 2552
rect 9809 1552 9929 2552
rect 10239 1552 10359 2552
rect 10801 1552 10921 2552
rect 11231 1552 11351 2552
rect 11793 1552 11913 2552
rect 12223 1552 12343 2552
rect 12785 1552 12905 2552
rect 13215 1552 13335 2552
rect 13777 1552 13897 2552
rect 14135 1552 14255 2552
<< mvpdiff >>
rect 708 4082 881 4152
rect 708 4048 745 4082
rect 779 4048 881 4082
rect 708 4014 881 4048
rect 708 3980 745 4014
rect 779 3980 881 4014
rect 708 3946 881 3980
rect 708 3912 745 3946
rect 779 3912 881 3946
rect 708 3878 881 3912
rect 708 3844 745 3878
rect 779 3844 881 3878
rect 708 3810 881 3844
rect 708 3776 745 3810
rect 779 3776 881 3810
rect 708 3742 881 3776
rect 708 3708 745 3742
rect 779 3708 881 3742
rect 708 3674 881 3708
rect 708 3640 745 3674
rect 779 3640 881 3674
rect 708 3606 881 3640
rect 708 3572 745 3606
rect 779 3572 881 3606
rect 708 3538 881 3572
rect 708 3504 745 3538
rect 779 3504 881 3538
rect 708 3470 881 3504
rect 708 3436 745 3470
rect 779 3436 881 3470
rect 708 3402 881 3436
rect 708 3368 745 3402
rect 779 3368 881 3402
rect 708 3334 881 3368
rect 708 3300 745 3334
rect 779 3300 881 3334
rect 708 3266 881 3300
rect 708 3232 745 3266
rect 779 3232 881 3266
rect 708 3198 881 3232
rect 708 3164 745 3198
rect 779 3164 881 3198
rect 708 3152 881 3164
rect 1001 4082 1311 4152
rect 1001 4048 1103 4082
rect 1137 4048 1175 4082
rect 1209 4048 1311 4082
rect 1001 4014 1311 4048
rect 1001 3980 1103 4014
rect 1137 3980 1175 4014
rect 1209 3980 1311 4014
rect 1001 3946 1311 3980
rect 1001 3912 1103 3946
rect 1137 3912 1175 3946
rect 1209 3912 1311 3946
rect 1001 3878 1311 3912
rect 1001 3844 1103 3878
rect 1137 3844 1175 3878
rect 1209 3844 1311 3878
rect 1001 3810 1311 3844
rect 1001 3776 1103 3810
rect 1137 3776 1175 3810
rect 1209 3776 1311 3810
rect 1001 3742 1311 3776
rect 1001 3708 1103 3742
rect 1137 3708 1175 3742
rect 1209 3708 1311 3742
rect 1001 3674 1311 3708
rect 1001 3640 1103 3674
rect 1137 3640 1175 3674
rect 1209 3640 1311 3674
rect 1001 3606 1311 3640
rect 1001 3572 1103 3606
rect 1137 3572 1175 3606
rect 1209 3572 1311 3606
rect 1001 3538 1311 3572
rect 1001 3504 1103 3538
rect 1137 3504 1175 3538
rect 1209 3504 1311 3538
rect 1001 3470 1311 3504
rect 1001 3436 1103 3470
rect 1137 3436 1175 3470
rect 1209 3436 1311 3470
rect 1001 3402 1311 3436
rect 1001 3368 1103 3402
rect 1137 3368 1175 3402
rect 1209 3368 1311 3402
rect 1001 3334 1311 3368
rect 1001 3300 1103 3334
rect 1137 3300 1175 3334
rect 1209 3300 1311 3334
rect 1001 3266 1311 3300
rect 1001 3232 1103 3266
rect 1137 3232 1175 3266
rect 1209 3232 1311 3266
rect 1001 3198 1311 3232
rect 1001 3164 1103 3198
rect 1137 3164 1175 3198
rect 1209 3164 1311 3198
rect 1001 3152 1311 3164
rect 1431 4082 1582 4152
rect 1722 4082 1873 4152
rect 1431 4048 1533 4082
rect 1567 4048 1582 4082
rect 1722 4048 1737 4082
rect 1771 4048 1873 4082
rect 1431 4014 1582 4048
rect 1722 4014 1873 4048
rect 1431 3980 1533 4014
rect 1567 3980 1582 4014
rect 1722 3980 1737 4014
rect 1771 3980 1873 4014
rect 1431 3946 1582 3980
rect 1722 3946 1873 3980
rect 1431 3912 1533 3946
rect 1567 3912 1582 3946
rect 1722 3912 1737 3946
rect 1771 3912 1873 3946
rect 1431 3878 1582 3912
rect 1722 3878 1873 3912
rect 1431 3844 1533 3878
rect 1567 3844 1582 3878
rect 1722 3844 1737 3878
rect 1771 3844 1873 3878
rect 1431 3810 1582 3844
rect 1722 3810 1873 3844
rect 1431 3776 1533 3810
rect 1567 3776 1582 3810
rect 1722 3776 1737 3810
rect 1771 3776 1873 3810
rect 1431 3742 1582 3776
rect 1722 3742 1873 3776
rect 1431 3708 1533 3742
rect 1567 3708 1582 3742
rect 1722 3708 1737 3742
rect 1771 3708 1873 3742
rect 1431 3674 1582 3708
rect 1722 3674 1873 3708
rect 1431 3640 1533 3674
rect 1567 3640 1582 3674
rect 1722 3640 1737 3674
rect 1771 3640 1873 3674
rect 1431 3606 1582 3640
rect 1722 3606 1873 3640
rect 1431 3572 1533 3606
rect 1567 3572 1582 3606
rect 1722 3572 1737 3606
rect 1771 3572 1873 3606
rect 1431 3538 1582 3572
rect 1722 3538 1873 3572
rect 1431 3504 1533 3538
rect 1567 3504 1582 3538
rect 1722 3504 1737 3538
rect 1771 3504 1873 3538
rect 1431 3470 1582 3504
rect 1722 3470 1873 3504
rect 1431 3436 1533 3470
rect 1567 3436 1582 3470
rect 1722 3436 1737 3470
rect 1771 3436 1873 3470
rect 1431 3402 1582 3436
rect 1722 3402 1873 3436
rect 1431 3368 1533 3402
rect 1567 3368 1582 3402
rect 1722 3368 1737 3402
rect 1771 3368 1873 3402
rect 1431 3334 1582 3368
rect 1722 3334 1873 3368
rect 1431 3300 1533 3334
rect 1567 3300 1582 3334
rect 1722 3300 1737 3334
rect 1771 3300 1873 3334
rect 1431 3266 1582 3300
rect 1722 3266 1873 3300
rect 1431 3232 1533 3266
rect 1567 3232 1582 3266
rect 1722 3232 1737 3266
rect 1771 3232 1873 3266
rect 1431 3198 1582 3232
rect 1722 3198 1873 3232
rect 1431 3164 1533 3198
rect 1567 3164 1582 3198
rect 1722 3164 1737 3198
rect 1771 3164 1873 3198
rect 1431 3152 1582 3164
rect 1722 3152 1873 3164
rect 1993 4082 2303 4152
rect 1993 4048 2095 4082
rect 2129 4048 2167 4082
rect 2201 4048 2303 4082
rect 1993 4014 2303 4048
rect 1993 3980 2095 4014
rect 2129 3980 2167 4014
rect 2201 3980 2303 4014
rect 1993 3946 2303 3980
rect 1993 3912 2095 3946
rect 2129 3912 2167 3946
rect 2201 3912 2303 3946
rect 1993 3878 2303 3912
rect 1993 3844 2095 3878
rect 2129 3844 2167 3878
rect 2201 3844 2303 3878
rect 1993 3810 2303 3844
rect 1993 3776 2095 3810
rect 2129 3776 2167 3810
rect 2201 3776 2303 3810
rect 1993 3742 2303 3776
rect 1993 3708 2095 3742
rect 2129 3708 2167 3742
rect 2201 3708 2303 3742
rect 1993 3674 2303 3708
rect 1993 3640 2095 3674
rect 2129 3640 2167 3674
rect 2201 3640 2303 3674
rect 1993 3606 2303 3640
rect 1993 3572 2095 3606
rect 2129 3572 2167 3606
rect 2201 3572 2303 3606
rect 1993 3538 2303 3572
rect 1993 3504 2095 3538
rect 2129 3504 2167 3538
rect 2201 3504 2303 3538
rect 1993 3470 2303 3504
rect 1993 3436 2095 3470
rect 2129 3436 2167 3470
rect 2201 3436 2303 3470
rect 1993 3402 2303 3436
rect 1993 3368 2095 3402
rect 2129 3368 2167 3402
rect 2201 3368 2303 3402
rect 1993 3334 2303 3368
rect 1993 3300 2095 3334
rect 2129 3300 2167 3334
rect 2201 3300 2303 3334
rect 1993 3266 2303 3300
rect 1993 3232 2095 3266
rect 2129 3232 2167 3266
rect 2201 3232 2303 3266
rect 1993 3198 2303 3232
rect 1993 3164 2095 3198
rect 2129 3164 2167 3198
rect 2201 3164 2303 3198
rect 1993 3152 2303 3164
rect 2423 4082 2574 4152
rect 2714 4082 2865 4152
rect 2423 4048 2525 4082
rect 2559 4048 2574 4082
rect 2714 4048 2729 4082
rect 2763 4048 2865 4082
rect 2423 4014 2574 4048
rect 2714 4014 2865 4048
rect 2423 3980 2525 4014
rect 2559 3980 2574 4014
rect 2714 3980 2729 4014
rect 2763 3980 2865 4014
rect 2423 3946 2574 3980
rect 2714 3946 2865 3980
rect 2423 3912 2525 3946
rect 2559 3912 2574 3946
rect 2714 3912 2729 3946
rect 2763 3912 2865 3946
rect 2423 3878 2574 3912
rect 2714 3878 2865 3912
rect 2423 3844 2525 3878
rect 2559 3844 2574 3878
rect 2714 3844 2729 3878
rect 2763 3844 2865 3878
rect 2423 3810 2574 3844
rect 2714 3810 2865 3844
rect 2423 3776 2525 3810
rect 2559 3776 2574 3810
rect 2714 3776 2729 3810
rect 2763 3776 2865 3810
rect 2423 3742 2574 3776
rect 2714 3742 2865 3776
rect 2423 3708 2525 3742
rect 2559 3708 2574 3742
rect 2714 3708 2729 3742
rect 2763 3708 2865 3742
rect 2423 3674 2574 3708
rect 2714 3674 2865 3708
rect 2423 3640 2525 3674
rect 2559 3640 2574 3674
rect 2714 3640 2729 3674
rect 2763 3640 2865 3674
rect 2423 3606 2574 3640
rect 2714 3606 2865 3640
rect 2423 3572 2525 3606
rect 2559 3572 2574 3606
rect 2714 3572 2729 3606
rect 2763 3572 2865 3606
rect 2423 3538 2574 3572
rect 2714 3538 2865 3572
rect 2423 3504 2525 3538
rect 2559 3504 2574 3538
rect 2714 3504 2729 3538
rect 2763 3504 2865 3538
rect 2423 3470 2574 3504
rect 2714 3470 2865 3504
rect 2423 3436 2525 3470
rect 2559 3436 2574 3470
rect 2714 3436 2729 3470
rect 2763 3436 2865 3470
rect 2423 3402 2574 3436
rect 2714 3402 2865 3436
rect 2423 3368 2525 3402
rect 2559 3368 2574 3402
rect 2714 3368 2729 3402
rect 2763 3368 2865 3402
rect 2423 3334 2574 3368
rect 2714 3334 2865 3368
rect 2423 3300 2525 3334
rect 2559 3300 2574 3334
rect 2714 3300 2729 3334
rect 2763 3300 2865 3334
rect 2423 3266 2574 3300
rect 2714 3266 2865 3300
rect 2423 3232 2525 3266
rect 2559 3232 2574 3266
rect 2714 3232 2729 3266
rect 2763 3232 2865 3266
rect 2423 3198 2574 3232
rect 2714 3198 2865 3232
rect 2423 3164 2525 3198
rect 2559 3164 2574 3198
rect 2714 3164 2729 3198
rect 2763 3164 2865 3198
rect 2423 3152 2574 3164
rect 2714 3152 2865 3164
rect 2985 4082 3295 4152
rect 2985 4048 3087 4082
rect 3121 4048 3159 4082
rect 3193 4048 3295 4082
rect 2985 4014 3295 4048
rect 2985 3980 3087 4014
rect 3121 3980 3159 4014
rect 3193 3980 3295 4014
rect 2985 3946 3295 3980
rect 2985 3912 3087 3946
rect 3121 3912 3159 3946
rect 3193 3912 3295 3946
rect 2985 3878 3295 3912
rect 2985 3844 3087 3878
rect 3121 3844 3159 3878
rect 3193 3844 3295 3878
rect 2985 3810 3295 3844
rect 2985 3776 3087 3810
rect 3121 3776 3159 3810
rect 3193 3776 3295 3810
rect 2985 3742 3295 3776
rect 2985 3708 3087 3742
rect 3121 3708 3159 3742
rect 3193 3708 3295 3742
rect 2985 3674 3295 3708
rect 2985 3640 3087 3674
rect 3121 3640 3159 3674
rect 3193 3640 3295 3674
rect 2985 3606 3295 3640
rect 2985 3572 3087 3606
rect 3121 3572 3159 3606
rect 3193 3572 3295 3606
rect 2985 3538 3295 3572
rect 2985 3504 3087 3538
rect 3121 3504 3159 3538
rect 3193 3504 3295 3538
rect 2985 3470 3295 3504
rect 2985 3436 3087 3470
rect 3121 3436 3159 3470
rect 3193 3436 3295 3470
rect 2985 3402 3295 3436
rect 2985 3368 3087 3402
rect 3121 3368 3159 3402
rect 3193 3368 3295 3402
rect 2985 3334 3295 3368
rect 2985 3300 3087 3334
rect 3121 3300 3159 3334
rect 3193 3300 3295 3334
rect 2985 3266 3295 3300
rect 2985 3232 3087 3266
rect 3121 3232 3159 3266
rect 3193 3232 3295 3266
rect 2985 3198 3295 3232
rect 2985 3164 3087 3198
rect 3121 3164 3159 3198
rect 3193 3164 3295 3198
rect 2985 3152 3295 3164
rect 3415 4082 3566 4152
rect 3706 4082 3857 4152
rect 3415 4048 3517 4082
rect 3551 4048 3566 4082
rect 3706 4048 3721 4082
rect 3755 4048 3857 4082
rect 3415 4014 3566 4048
rect 3706 4014 3857 4048
rect 3415 3980 3517 4014
rect 3551 3980 3566 4014
rect 3706 3980 3721 4014
rect 3755 3980 3857 4014
rect 3415 3946 3566 3980
rect 3706 3946 3857 3980
rect 3415 3912 3517 3946
rect 3551 3912 3566 3946
rect 3706 3912 3721 3946
rect 3755 3912 3857 3946
rect 3415 3878 3566 3912
rect 3706 3878 3857 3912
rect 3415 3844 3517 3878
rect 3551 3844 3566 3878
rect 3706 3844 3721 3878
rect 3755 3844 3857 3878
rect 3415 3810 3566 3844
rect 3706 3810 3857 3844
rect 3415 3776 3517 3810
rect 3551 3776 3566 3810
rect 3706 3776 3721 3810
rect 3755 3776 3857 3810
rect 3415 3742 3566 3776
rect 3706 3742 3857 3776
rect 3415 3708 3517 3742
rect 3551 3708 3566 3742
rect 3706 3708 3721 3742
rect 3755 3708 3857 3742
rect 3415 3674 3566 3708
rect 3706 3674 3857 3708
rect 3415 3640 3517 3674
rect 3551 3640 3566 3674
rect 3706 3640 3721 3674
rect 3755 3640 3857 3674
rect 3415 3606 3566 3640
rect 3706 3606 3857 3640
rect 3415 3572 3517 3606
rect 3551 3572 3566 3606
rect 3706 3572 3721 3606
rect 3755 3572 3857 3606
rect 3415 3538 3566 3572
rect 3706 3538 3857 3572
rect 3415 3504 3517 3538
rect 3551 3504 3566 3538
rect 3706 3504 3721 3538
rect 3755 3504 3857 3538
rect 3415 3470 3566 3504
rect 3706 3470 3857 3504
rect 3415 3436 3517 3470
rect 3551 3436 3566 3470
rect 3706 3436 3721 3470
rect 3755 3436 3857 3470
rect 3415 3402 3566 3436
rect 3706 3402 3857 3436
rect 3415 3368 3517 3402
rect 3551 3368 3566 3402
rect 3706 3368 3721 3402
rect 3755 3368 3857 3402
rect 3415 3334 3566 3368
rect 3706 3334 3857 3368
rect 3415 3300 3517 3334
rect 3551 3300 3566 3334
rect 3706 3300 3721 3334
rect 3755 3300 3857 3334
rect 3415 3266 3566 3300
rect 3706 3266 3857 3300
rect 3415 3232 3517 3266
rect 3551 3232 3566 3266
rect 3706 3232 3721 3266
rect 3755 3232 3857 3266
rect 3415 3198 3566 3232
rect 3706 3198 3857 3232
rect 3415 3164 3517 3198
rect 3551 3164 3566 3198
rect 3706 3164 3721 3198
rect 3755 3164 3857 3198
rect 3415 3152 3566 3164
rect 3706 3152 3857 3164
rect 3977 4082 4287 4152
rect 3977 4048 4079 4082
rect 4113 4048 4151 4082
rect 4185 4048 4287 4082
rect 3977 4014 4287 4048
rect 3977 3980 4079 4014
rect 4113 3980 4151 4014
rect 4185 3980 4287 4014
rect 3977 3946 4287 3980
rect 3977 3912 4079 3946
rect 4113 3912 4151 3946
rect 4185 3912 4287 3946
rect 3977 3878 4287 3912
rect 3977 3844 4079 3878
rect 4113 3844 4151 3878
rect 4185 3844 4287 3878
rect 3977 3810 4287 3844
rect 3977 3776 4079 3810
rect 4113 3776 4151 3810
rect 4185 3776 4287 3810
rect 3977 3742 4287 3776
rect 3977 3708 4079 3742
rect 4113 3708 4151 3742
rect 4185 3708 4287 3742
rect 3977 3674 4287 3708
rect 3977 3640 4079 3674
rect 4113 3640 4151 3674
rect 4185 3640 4287 3674
rect 3977 3606 4287 3640
rect 3977 3572 4079 3606
rect 4113 3572 4151 3606
rect 4185 3572 4287 3606
rect 3977 3538 4287 3572
rect 3977 3504 4079 3538
rect 4113 3504 4151 3538
rect 4185 3504 4287 3538
rect 3977 3470 4287 3504
rect 3977 3436 4079 3470
rect 4113 3436 4151 3470
rect 4185 3436 4287 3470
rect 3977 3402 4287 3436
rect 3977 3368 4079 3402
rect 4113 3368 4151 3402
rect 4185 3368 4287 3402
rect 3977 3334 4287 3368
rect 3977 3300 4079 3334
rect 4113 3300 4151 3334
rect 4185 3300 4287 3334
rect 3977 3266 4287 3300
rect 3977 3232 4079 3266
rect 4113 3232 4151 3266
rect 4185 3232 4287 3266
rect 3977 3198 4287 3232
rect 3977 3164 4079 3198
rect 4113 3164 4151 3198
rect 4185 3164 4287 3198
rect 3977 3152 4287 3164
rect 4407 4082 4558 4152
rect 4698 4082 4849 4152
rect 4407 4048 4509 4082
rect 4543 4048 4558 4082
rect 4698 4048 4713 4082
rect 4747 4048 4849 4082
rect 4407 4014 4558 4048
rect 4698 4014 4849 4048
rect 4407 3980 4509 4014
rect 4543 3980 4558 4014
rect 4698 3980 4713 4014
rect 4747 3980 4849 4014
rect 4407 3946 4558 3980
rect 4698 3946 4849 3980
rect 4407 3912 4509 3946
rect 4543 3912 4558 3946
rect 4698 3912 4713 3946
rect 4747 3912 4849 3946
rect 4407 3878 4558 3912
rect 4698 3878 4849 3912
rect 4407 3844 4509 3878
rect 4543 3844 4558 3878
rect 4698 3844 4713 3878
rect 4747 3844 4849 3878
rect 4407 3810 4558 3844
rect 4698 3810 4849 3844
rect 4407 3776 4509 3810
rect 4543 3776 4558 3810
rect 4698 3776 4713 3810
rect 4747 3776 4849 3810
rect 4407 3742 4558 3776
rect 4698 3742 4849 3776
rect 4407 3708 4509 3742
rect 4543 3708 4558 3742
rect 4698 3708 4713 3742
rect 4747 3708 4849 3742
rect 4407 3674 4558 3708
rect 4698 3674 4849 3708
rect 4407 3640 4509 3674
rect 4543 3640 4558 3674
rect 4698 3640 4713 3674
rect 4747 3640 4849 3674
rect 4407 3606 4558 3640
rect 4698 3606 4849 3640
rect 4407 3572 4509 3606
rect 4543 3572 4558 3606
rect 4698 3572 4713 3606
rect 4747 3572 4849 3606
rect 4407 3538 4558 3572
rect 4698 3538 4849 3572
rect 4407 3504 4509 3538
rect 4543 3504 4558 3538
rect 4698 3504 4713 3538
rect 4747 3504 4849 3538
rect 4407 3470 4558 3504
rect 4698 3470 4849 3504
rect 4407 3436 4509 3470
rect 4543 3436 4558 3470
rect 4698 3436 4713 3470
rect 4747 3436 4849 3470
rect 4407 3402 4558 3436
rect 4698 3402 4849 3436
rect 4407 3368 4509 3402
rect 4543 3368 4558 3402
rect 4698 3368 4713 3402
rect 4747 3368 4849 3402
rect 4407 3334 4558 3368
rect 4698 3334 4849 3368
rect 4407 3300 4509 3334
rect 4543 3300 4558 3334
rect 4698 3300 4713 3334
rect 4747 3300 4849 3334
rect 4407 3266 4558 3300
rect 4698 3266 4849 3300
rect 4407 3232 4509 3266
rect 4543 3232 4558 3266
rect 4698 3232 4713 3266
rect 4747 3232 4849 3266
rect 4407 3198 4558 3232
rect 4698 3198 4849 3232
rect 4407 3164 4509 3198
rect 4543 3164 4558 3198
rect 4698 3164 4713 3198
rect 4747 3164 4849 3198
rect 4407 3152 4558 3164
rect 4698 3152 4849 3164
rect 4969 4082 5279 4152
rect 4969 4048 5071 4082
rect 5105 4048 5143 4082
rect 5177 4048 5279 4082
rect 4969 4014 5279 4048
rect 4969 3980 5071 4014
rect 5105 3980 5143 4014
rect 5177 3980 5279 4014
rect 4969 3946 5279 3980
rect 4969 3912 5071 3946
rect 5105 3912 5143 3946
rect 5177 3912 5279 3946
rect 4969 3878 5279 3912
rect 4969 3844 5071 3878
rect 5105 3844 5143 3878
rect 5177 3844 5279 3878
rect 4969 3810 5279 3844
rect 4969 3776 5071 3810
rect 5105 3776 5143 3810
rect 5177 3776 5279 3810
rect 4969 3742 5279 3776
rect 4969 3708 5071 3742
rect 5105 3708 5143 3742
rect 5177 3708 5279 3742
rect 4969 3674 5279 3708
rect 4969 3640 5071 3674
rect 5105 3640 5143 3674
rect 5177 3640 5279 3674
rect 4969 3606 5279 3640
rect 4969 3572 5071 3606
rect 5105 3572 5143 3606
rect 5177 3572 5279 3606
rect 4969 3538 5279 3572
rect 4969 3504 5071 3538
rect 5105 3504 5143 3538
rect 5177 3504 5279 3538
rect 4969 3470 5279 3504
rect 4969 3436 5071 3470
rect 5105 3436 5143 3470
rect 5177 3436 5279 3470
rect 4969 3402 5279 3436
rect 4969 3368 5071 3402
rect 5105 3368 5143 3402
rect 5177 3368 5279 3402
rect 4969 3334 5279 3368
rect 4969 3300 5071 3334
rect 5105 3300 5143 3334
rect 5177 3300 5279 3334
rect 4969 3266 5279 3300
rect 4969 3232 5071 3266
rect 5105 3232 5143 3266
rect 5177 3232 5279 3266
rect 4969 3198 5279 3232
rect 4969 3164 5071 3198
rect 5105 3164 5143 3198
rect 5177 3164 5279 3198
rect 4969 3152 5279 3164
rect 5399 4082 5550 4152
rect 5690 4082 5841 4152
rect 5399 4048 5501 4082
rect 5535 4048 5550 4082
rect 5690 4048 5705 4082
rect 5739 4048 5841 4082
rect 5399 4014 5550 4048
rect 5690 4014 5841 4048
rect 5399 3980 5501 4014
rect 5535 3980 5550 4014
rect 5690 3980 5705 4014
rect 5739 3980 5841 4014
rect 5399 3946 5550 3980
rect 5690 3946 5841 3980
rect 5399 3912 5501 3946
rect 5535 3912 5550 3946
rect 5690 3912 5705 3946
rect 5739 3912 5841 3946
rect 5399 3878 5550 3912
rect 5690 3878 5841 3912
rect 5399 3844 5501 3878
rect 5535 3844 5550 3878
rect 5690 3844 5705 3878
rect 5739 3844 5841 3878
rect 5399 3810 5550 3844
rect 5690 3810 5841 3844
rect 5399 3776 5501 3810
rect 5535 3776 5550 3810
rect 5690 3776 5705 3810
rect 5739 3776 5841 3810
rect 5399 3742 5550 3776
rect 5690 3742 5841 3776
rect 5399 3708 5501 3742
rect 5535 3708 5550 3742
rect 5690 3708 5705 3742
rect 5739 3708 5841 3742
rect 5399 3674 5550 3708
rect 5690 3674 5841 3708
rect 5399 3640 5501 3674
rect 5535 3640 5550 3674
rect 5690 3640 5705 3674
rect 5739 3640 5841 3674
rect 5399 3606 5550 3640
rect 5690 3606 5841 3640
rect 5399 3572 5501 3606
rect 5535 3572 5550 3606
rect 5690 3572 5705 3606
rect 5739 3572 5841 3606
rect 5399 3538 5550 3572
rect 5690 3538 5841 3572
rect 5399 3504 5501 3538
rect 5535 3504 5550 3538
rect 5690 3504 5705 3538
rect 5739 3504 5841 3538
rect 5399 3470 5550 3504
rect 5690 3470 5841 3504
rect 5399 3436 5501 3470
rect 5535 3436 5550 3470
rect 5690 3436 5705 3470
rect 5739 3436 5841 3470
rect 5399 3402 5550 3436
rect 5690 3402 5841 3436
rect 5399 3368 5501 3402
rect 5535 3368 5550 3402
rect 5690 3368 5705 3402
rect 5739 3368 5841 3402
rect 5399 3334 5550 3368
rect 5690 3334 5841 3368
rect 5399 3300 5501 3334
rect 5535 3300 5550 3334
rect 5690 3300 5705 3334
rect 5739 3300 5841 3334
rect 5399 3266 5550 3300
rect 5690 3266 5841 3300
rect 5399 3232 5501 3266
rect 5535 3232 5550 3266
rect 5690 3232 5705 3266
rect 5739 3232 5841 3266
rect 5399 3198 5550 3232
rect 5690 3198 5841 3232
rect 5399 3164 5501 3198
rect 5535 3164 5550 3198
rect 5690 3164 5705 3198
rect 5739 3164 5841 3198
rect 5399 3152 5550 3164
rect 5690 3152 5841 3164
rect 5961 4082 6271 4152
rect 5961 4048 6063 4082
rect 6097 4048 6135 4082
rect 6169 4048 6271 4082
rect 5961 4014 6271 4048
rect 5961 3980 6063 4014
rect 6097 3980 6135 4014
rect 6169 3980 6271 4014
rect 5961 3946 6271 3980
rect 5961 3912 6063 3946
rect 6097 3912 6135 3946
rect 6169 3912 6271 3946
rect 5961 3878 6271 3912
rect 5961 3844 6063 3878
rect 6097 3844 6135 3878
rect 6169 3844 6271 3878
rect 5961 3810 6271 3844
rect 5961 3776 6063 3810
rect 6097 3776 6135 3810
rect 6169 3776 6271 3810
rect 5961 3742 6271 3776
rect 5961 3708 6063 3742
rect 6097 3708 6135 3742
rect 6169 3708 6271 3742
rect 5961 3674 6271 3708
rect 5961 3640 6063 3674
rect 6097 3640 6135 3674
rect 6169 3640 6271 3674
rect 5961 3606 6271 3640
rect 5961 3572 6063 3606
rect 6097 3572 6135 3606
rect 6169 3572 6271 3606
rect 5961 3538 6271 3572
rect 5961 3504 6063 3538
rect 6097 3504 6135 3538
rect 6169 3504 6271 3538
rect 5961 3470 6271 3504
rect 5961 3436 6063 3470
rect 6097 3436 6135 3470
rect 6169 3436 6271 3470
rect 5961 3402 6271 3436
rect 5961 3368 6063 3402
rect 6097 3368 6135 3402
rect 6169 3368 6271 3402
rect 5961 3334 6271 3368
rect 5961 3300 6063 3334
rect 6097 3300 6135 3334
rect 6169 3300 6271 3334
rect 5961 3266 6271 3300
rect 5961 3232 6063 3266
rect 6097 3232 6135 3266
rect 6169 3232 6271 3266
rect 5961 3198 6271 3232
rect 5961 3164 6063 3198
rect 6097 3164 6135 3198
rect 6169 3164 6271 3198
rect 5961 3152 6271 3164
rect 6391 4082 6542 4152
rect 6682 4082 6833 4152
rect 6391 4048 6493 4082
rect 6527 4048 6542 4082
rect 6682 4048 6697 4082
rect 6731 4048 6833 4082
rect 6391 4014 6542 4048
rect 6682 4014 6833 4048
rect 6391 3980 6493 4014
rect 6527 3980 6542 4014
rect 6682 3980 6697 4014
rect 6731 3980 6833 4014
rect 6391 3946 6542 3980
rect 6682 3946 6833 3980
rect 6391 3912 6493 3946
rect 6527 3912 6542 3946
rect 6682 3912 6697 3946
rect 6731 3912 6833 3946
rect 6391 3878 6542 3912
rect 6682 3878 6833 3912
rect 6391 3844 6493 3878
rect 6527 3844 6542 3878
rect 6682 3844 6697 3878
rect 6731 3844 6833 3878
rect 6391 3810 6542 3844
rect 6682 3810 6833 3844
rect 6391 3776 6493 3810
rect 6527 3776 6542 3810
rect 6682 3776 6697 3810
rect 6731 3776 6833 3810
rect 6391 3742 6542 3776
rect 6682 3742 6833 3776
rect 6391 3708 6493 3742
rect 6527 3708 6542 3742
rect 6682 3708 6697 3742
rect 6731 3708 6833 3742
rect 6391 3674 6542 3708
rect 6682 3674 6833 3708
rect 6391 3640 6493 3674
rect 6527 3640 6542 3674
rect 6682 3640 6697 3674
rect 6731 3640 6833 3674
rect 6391 3606 6542 3640
rect 6682 3606 6833 3640
rect 6391 3572 6493 3606
rect 6527 3572 6542 3606
rect 6682 3572 6697 3606
rect 6731 3572 6833 3606
rect 6391 3538 6542 3572
rect 6682 3538 6833 3572
rect 6391 3504 6493 3538
rect 6527 3504 6542 3538
rect 6682 3504 6697 3538
rect 6731 3504 6833 3538
rect 6391 3470 6542 3504
rect 6682 3470 6833 3504
rect 6391 3436 6493 3470
rect 6527 3436 6542 3470
rect 6682 3436 6697 3470
rect 6731 3436 6833 3470
rect 6391 3402 6542 3436
rect 6682 3402 6833 3436
rect 6391 3368 6493 3402
rect 6527 3368 6542 3402
rect 6682 3368 6697 3402
rect 6731 3368 6833 3402
rect 6391 3334 6542 3368
rect 6682 3334 6833 3368
rect 6391 3300 6493 3334
rect 6527 3300 6542 3334
rect 6682 3300 6697 3334
rect 6731 3300 6833 3334
rect 6391 3266 6542 3300
rect 6682 3266 6833 3300
rect 6391 3232 6493 3266
rect 6527 3232 6542 3266
rect 6682 3232 6697 3266
rect 6731 3232 6833 3266
rect 6391 3198 6542 3232
rect 6682 3198 6833 3232
rect 6391 3164 6493 3198
rect 6527 3164 6542 3198
rect 6682 3164 6697 3198
rect 6731 3164 6833 3198
rect 6391 3152 6542 3164
rect 6682 3152 6833 3164
rect 6953 4082 7263 4152
rect 6953 4048 7055 4082
rect 7089 4048 7127 4082
rect 7161 4048 7263 4082
rect 6953 4014 7263 4048
rect 6953 3980 7055 4014
rect 7089 3980 7127 4014
rect 7161 3980 7263 4014
rect 6953 3946 7263 3980
rect 6953 3912 7055 3946
rect 7089 3912 7127 3946
rect 7161 3912 7263 3946
rect 6953 3878 7263 3912
rect 6953 3844 7055 3878
rect 7089 3844 7127 3878
rect 7161 3844 7263 3878
rect 6953 3810 7263 3844
rect 6953 3776 7055 3810
rect 7089 3776 7127 3810
rect 7161 3776 7263 3810
rect 6953 3742 7263 3776
rect 6953 3708 7055 3742
rect 7089 3708 7127 3742
rect 7161 3708 7263 3742
rect 6953 3674 7263 3708
rect 6953 3640 7055 3674
rect 7089 3640 7127 3674
rect 7161 3640 7263 3674
rect 6953 3606 7263 3640
rect 6953 3572 7055 3606
rect 7089 3572 7127 3606
rect 7161 3572 7263 3606
rect 6953 3538 7263 3572
rect 6953 3504 7055 3538
rect 7089 3504 7127 3538
rect 7161 3504 7263 3538
rect 6953 3470 7263 3504
rect 6953 3436 7055 3470
rect 7089 3436 7127 3470
rect 7161 3436 7263 3470
rect 6953 3402 7263 3436
rect 6953 3368 7055 3402
rect 7089 3368 7127 3402
rect 7161 3368 7263 3402
rect 6953 3334 7263 3368
rect 6953 3300 7055 3334
rect 7089 3300 7127 3334
rect 7161 3300 7263 3334
rect 6953 3266 7263 3300
rect 6953 3232 7055 3266
rect 7089 3232 7127 3266
rect 7161 3232 7263 3266
rect 6953 3198 7263 3232
rect 6953 3164 7055 3198
rect 7089 3164 7127 3198
rect 7161 3164 7263 3198
rect 6953 3152 7263 3164
rect 7383 4082 7534 4152
rect 7674 4082 7825 4152
rect 7383 4048 7485 4082
rect 7519 4048 7534 4082
rect 7674 4048 7689 4082
rect 7723 4048 7825 4082
rect 7383 4014 7534 4048
rect 7674 4014 7825 4048
rect 7383 3980 7485 4014
rect 7519 3980 7534 4014
rect 7674 3980 7689 4014
rect 7723 3980 7825 4014
rect 7383 3946 7534 3980
rect 7674 3946 7825 3980
rect 7383 3912 7485 3946
rect 7519 3912 7534 3946
rect 7674 3912 7689 3946
rect 7723 3912 7825 3946
rect 7383 3878 7534 3912
rect 7674 3878 7825 3912
rect 7383 3844 7485 3878
rect 7519 3844 7534 3878
rect 7674 3844 7689 3878
rect 7723 3844 7825 3878
rect 7383 3810 7534 3844
rect 7674 3810 7825 3844
rect 7383 3776 7485 3810
rect 7519 3776 7534 3810
rect 7674 3776 7689 3810
rect 7723 3776 7825 3810
rect 7383 3742 7534 3776
rect 7674 3742 7825 3776
rect 7383 3708 7485 3742
rect 7519 3708 7534 3742
rect 7674 3708 7689 3742
rect 7723 3708 7825 3742
rect 7383 3674 7534 3708
rect 7674 3674 7825 3708
rect 7383 3640 7485 3674
rect 7519 3640 7534 3674
rect 7674 3640 7689 3674
rect 7723 3640 7825 3674
rect 7383 3606 7534 3640
rect 7674 3606 7825 3640
rect 7383 3572 7485 3606
rect 7519 3572 7534 3606
rect 7674 3572 7689 3606
rect 7723 3572 7825 3606
rect 7383 3538 7534 3572
rect 7674 3538 7825 3572
rect 7383 3504 7485 3538
rect 7519 3504 7534 3538
rect 7674 3504 7689 3538
rect 7723 3504 7825 3538
rect 7383 3470 7534 3504
rect 7674 3470 7825 3504
rect 7383 3436 7485 3470
rect 7519 3436 7534 3470
rect 7674 3436 7689 3470
rect 7723 3436 7825 3470
rect 7383 3402 7534 3436
rect 7674 3402 7825 3436
rect 7383 3368 7485 3402
rect 7519 3368 7534 3402
rect 7674 3368 7689 3402
rect 7723 3368 7825 3402
rect 7383 3334 7534 3368
rect 7674 3334 7825 3368
rect 7383 3300 7485 3334
rect 7519 3300 7534 3334
rect 7674 3300 7689 3334
rect 7723 3300 7825 3334
rect 7383 3266 7534 3300
rect 7674 3266 7825 3300
rect 7383 3232 7485 3266
rect 7519 3232 7534 3266
rect 7674 3232 7689 3266
rect 7723 3232 7825 3266
rect 7383 3198 7534 3232
rect 7674 3198 7825 3232
rect 7383 3164 7485 3198
rect 7519 3164 7534 3198
rect 7674 3164 7689 3198
rect 7723 3164 7825 3198
rect 7383 3152 7534 3164
rect 7674 3152 7825 3164
rect 7945 4082 8255 4152
rect 7945 4048 8047 4082
rect 8081 4048 8119 4082
rect 8153 4048 8255 4082
rect 7945 4014 8255 4048
rect 7945 3980 8047 4014
rect 8081 3980 8119 4014
rect 8153 3980 8255 4014
rect 7945 3946 8255 3980
rect 7945 3912 8047 3946
rect 8081 3912 8119 3946
rect 8153 3912 8255 3946
rect 7945 3878 8255 3912
rect 7945 3844 8047 3878
rect 8081 3844 8119 3878
rect 8153 3844 8255 3878
rect 7945 3810 8255 3844
rect 7945 3776 8047 3810
rect 8081 3776 8119 3810
rect 8153 3776 8255 3810
rect 7945 3742 8255 3776
rect 7945 3708 8047 3742
rect 8081 3708 8119 3742
rect 8153 3708 8255 3742
rect 7945 3674 8255 3708
rect 7945 3640 8047 3674
rect 8081 3640 8119 3674
rect 8153 3640 8255 3674
rect 7945 3606 8255 3640
rect 7945 3572 8047 3606
rect 8081 3572 8119 3606
rect 8153 3572 8255 3606
rect 7945 3538 8255 3572
rect 7945 3504 8047 3538
rect 8081 3504 8119 3538
rect 8153 3504 8255 3538
rect 7945 3470 8255 3504
rect 7945 3436 8047 3470
rect 8081 3436 8119 3470
rect 8153 3436 8255 3470
rect 7945 3402 8255 3436
rect 7945 3368 8047 3402
rect 8081 3368 8119 3402
rect 8153 3368 8255 3402
rect 7945 3334 8255 3368
rect 7945 3300 8047 3334
rect 8081 3300 8119 3334
rect 8153 3300 8255 3334
rect 7945 3266 8255 3300
rect 7945 3232 8047 3266
rect 8081 3232 8119 3266
rect 8153 3232 8255 3266
rect 7945 3198 8255 3232
rect 7945 3164 8047 3198
rect 8081 3164 8119 3198
rect 8153 3164 8255 3198
rect 7945 3152 8255 3164
rect 8375 4082 8526 4152
rect 8666 4082 8817 4152
rect 8375 4048 8477 4082
rect 8511 4048 8526 4082
rect 8666 4048 8681 4082
rect 8715 4048 8817 4082
rect 8375 4014 8526 4048
rect 8666 4014 8817 4048
rect 8375 3980 8477 4014
rect 8511 3980 8526 4014
rect 8666 3980 8681 4014
rect 8715 3980 8817 4014
rect 8375 3946 8526 3980
rect 8666 3946 8817 3980
rect 8375 3912 8477 3946
rect 8511 3912 8526 3946
rect 8666 3912 8681 3946
rect 8715 3912 8817 3946
rect 8375 3878 8526 3912
rect 8666 3878 8817 3912
rect 8375 3844 8477 3878
rect 8511 3844 8526 3878
rect 8666 3844 8681 3878
rect 8715 3844 8817 3878
rect 8375 3810 8526 3844
rect 8666 3810 8817 3844
rect 8375 3776 8477 3810
rect 8511 3776 8526 3810
rect 8666 3776 8681 3810
rect 8715 3776 8817 3810
rect 8375 3742 8526 3776
rect 8666 3742 8817 3776
rect 8375 3708 8477 3742
rect 8511 3708 8526 3742
rect 8666 3708 8681 3742
rect 8715 3708 8817 3742
rect 8375 3674 8526 3708
rect 8666 3674 8817 3708
rect 8375 3640 8477 3674
rect 8511 3640 8526 3674
rect 8666 3640 8681 3674
rect 8715 3640 8817 3674
rect 8375 3606 8526 3640
rect 8666 3606 8817 3640
rect 8375 3572 8477 3606
rect 8511 3572 8526 3606
rect 8666 3572 8681 3606
rect 8715 3572 8817 3606
rect 8375 3538 8526 3572
rect 8666 3538 8817 3572
rect 8375 3504 8477 3538
rect 8511 3504 8526 3538
rect 8666 3504 8681 3538
rect 8715 3504 8817 3538
rect 8375 3470 8526 3504
rect 8666 3470 8817 3504
rect 8375 3436 8477 3470
rect 8511 3436 8526 3470
rect 8666 3436 8681 3470
rect 8715 3436 8817 3470
rect 8375 3402 8526 3436
rect 8666 3402 8817 3436
rect 8375 3368 8477 3402
rect 8511 3368 8526 3402
rect 8666 3368 8681 3402
rect 8715 3368 8817 3402
rect 8375 3334 8526 3368
rect 8666 3334 8817 3368
rect 8375 3300 8477 3334
rect 8511 3300 8526 3334
rect 8666 3300 8681 3334
rect 8715 3300 8817 3334
rect 8375 3266 8526 3300
rect 8666 3266 8817 3300
rect 8375 3232 8477 3266
rect 8511 3232 8526 3266
rect 8666 3232 8681 3266
rect 8715 3232 8817 3266
rect 8375 3198 8526 3232
rect 8666 3198 8817 3232
rect 8375 3164 8477 3198
rect 8511 3164 8526 3198
rect 8666 3164 8681 3198
rect 8715 3164 8817 3198
rect 8375 3152 8526 3164
rect 8666 3152 8817 3164
rect 8937 4082 9247 4152
rect 8937 4048 9039 4082
rect 9073 4048 9111 4082
rect 9145 4048 9247 4082
rect 8937 4014 9247 4048
rect 8937 3980 9039 4014
rect 9073 3980 9111 4014
rect 9145 3980 9247 4014
rect 8937 3946 9247 3980
rect 8937 3912 9039 3946
rect 9073 3912 9111 3946
rect 9145 3912 9247 3946
rect 8937 3878 9247 3912
rect 8937 3844 9039 3878
rect 9073 3844 9111 3878
rect 9145 3844 9247 3878
rect 8937 3810 9247 3844
rect 8937 3776 9039 3810
rect 9073 3776 9111 3810
rect 9145 3776 9247 3810
rect 8937 3742 9247 3776
rect 8937 3708 9039 3742
rect 9073 3708 9111 3742
rect 9145 3708 9247 3742
rect 8937 3674 9247 3708
rect 8937 3640 9039 3674
rect 9073 3640 9111 3674
rect 9145 3640 9247 3674
rect 8937 3606 9247 3640
rect 8937 3572 9039 3606
rect 9073 3572 9111 3606
rect 9145 3572 9247 3606
rect 8937 3538 9247 3572
rect 8937 3504 9039 3538
rect 9073 3504 9111 3538
rect 9145 3504 9247 3538
rect 8937 3470 9247 3504
rect 8937 3436 9039 3470
rect 9073 3436 9111 3470
rect 9145 3436 9247 3470
rect 8937 3402 9247 3436
rect 8937 3368 9039 3402
rect 9073 3368 9111 3402
rect 9145 3368 9247 3402
rect 8937 3334 9247 3368
rect 8937 3300 9039 3334
rect 9073 3300 9111 3334
rect 9145 3300 9247 3334
rect 8937 3266 9247 3300
rect 8937 3232 9039 3266
rect 9073 3232 9111 3266
rect 9145 3232 9247 3266
rect 8937 3198 9247 3232
rect 8937 3164 9039 3198
rect 9073 3164 9111 3198
rect 9145 3164 9247 3198
rect 8937 3152 9247 3164
rect 9367 4082 9518 4152
rect 9658 4082 9809 4152
rect 9367 4048 9469 4082
rect 9503 4048 9518 4082
rect 9658 4048 9673 4082
rect 9707 4048 9809 4082
rect 9367 4014 9518 4048
rect 9658 4014 9809 4048
rect 9367 3980 9469 4014
rect 9503 3980 9518 4014
rect 9658 3980 9673 4014
rect 9707 3980 9809 4014
rect 9367 3946 9518 3980
rect 9658 3946 9809 3980
rect 9367 3912 9469 3946
rect 9503 3912 9518 3946
rect 9658 3912 9673 3946
rect 9707 3912 9809 3946
rect 9367 3878 9518 3912
rect 9658 3878 9809 3912
rect 9367 3844 9469 3878
rect 9503 3844 9518 3878
rect 9658 3844 9673 3878
rect 9707 3844 9809 3878
rect 9367 3810 9518 3844
rect 9658 3810 9809 3844
rect 9367 3776 9469 3810
rect 9503 3776 9518 3810
rect 9658 3776 9673 3810
rect 9707 3776 9809 3810
rect 9367 3742 9518 3776
rect 9658 3742 9809 3776
rect 9367 3708 9469 3742
rect 9503 3708 9518 3742
rect 9658 3708 9673 3742
rect 9707 3708 9809 3742
rect 9367 3674 9518 3708
rect 9658 3674 9809 3708
rect 9367 3640 9469 3674
rect 9503 3640 9518 3674
rect 9658 3640 9673 3674
rect 9707 3640 9809 3674
rect 9367 3606 9518 3640
rect 9658 3606 9809 3640
rect 9367 3572 9469 3606
rect 9503 3572 9518 3606
rect 9658 3572 9673 3606
rect 9707 3572 9809 3606
rect 9367 3538 9518 3572
rect 9658 3538 9809 3572
rect 9367 3504 9469 3538
rect 9503 3504 9518 3538
rect 9658 3504 9673 3538
rect 9707 3504 9809 3538
rect 9367 3470 9518 3504
rect 9658 3470 9809 3504
rect 9367 3436 9469 3470
rect 9503 3436 9518 3470
rect 9658 3436 9673 3470
rect 9707 3436 9809 3470
rect 9367 3402 9518 3436
rect 9658 3402 9809 3436
rect 9367 3368 9469 3402
rect 9503 3368 9518 3402
rect 9658 3368 9673 3402
rect 9707 3368 9809 3402
rect 9367 3334 9518 3368
rect 9658 3334 9809 3368
rect 9367 3300 9469 3334
rect 9503 3300 9518 3334
rect 9658 3300 9673 3334
rect 9707 3300 9809 3334
rect 9367 3266 9518 3300
rect 9658 3266 9809 3300
rect 9367 3232 9469 3266
rect 9503 3232 9518 3266
rect 9658 3232 9673 3266
rect 9707 3232 9809 3266
rect 9367 3198 9518 3232
rect 9658 3198 9809 3232
rect 9367 3164 9469 3198
rect 9503 3164 9518 3198
rect 9658 3164 9673 3198
rect 9707 3164 9809 3198
rect 9367 3152 9518 3164
rect 9658 3152 9809 3164
rect 9929 4082 10239 4152
rect 9929 4048 10031 4082
rect 10065 4048 10103 4082
rect 10137 4048 10239 4082
rect 9929 4014 10239 4048
rect 9929 3980 10031 4014
rect 10065 3980 10103 4014
rect 10137 3980 10239 4014
rect 9929 3946 10239 3980
rect 9929 3912 10031 3946
rect 10065 3912 10103 3946
rect 10137 3912 10239 3946
rect 9929 3878 10239 3912
rect 9929 3844 10031 3878
rect 10065 3844 10103 3878
rect 10137 3844 10239 3878
rect 9929 3810 10239 3844
rect 9929 3776 10031 3810
rect 10065 3776 10103 3810
rect 10137 3776 10239 3810
rect 9929 3742 10239 3776
rect 9929 3708 10031 3742
rect 10065 3708 10103 3742
rect 10137 3708 10239 3742
rect 9929 3674 10239 3708
rect 9929 3640 10031 3674
rect 10065 3640 10103 3674
rect 10137 3640 10239 3674
rect 9929 3606 10239 3640
rect 9929 3572 10031 3606
rect 10065 3572 10103 3606
rect 10137 3572 10239 3606
rect 9929 3538 10239 3572
rect 9929 3504 10031 3538
rect 10065 3504 10103 3538
rect 10137 3504 10239 3538
rect 9929 3470 10239 3504
rect 9929 3436 10031 3470
rect 10065 3436 10103 3470
rect 10137 3436 10239 3470
rect 9929 3402 10239 3436
rect 9929 3368 10031 3402
rect 10065 3368 10103 3402
rect 10137 3368 10239 3402
rect 9929 3334 10239 3368
rect 9929 3300 10031 3334
rect 10065 3300 10103 3334
rect 10137 3300 10239 3334
rect 9929 3266 10239 3300
rect 9929 3232 10031 3266
rect 10065 3232 10103 3266
rect 10137 3232 10239 3266
rect 9929 3198 10239 3232
rect 9929 3164 10031 3198
rect 10065 3164 10103 3198
rect 10137 3164 10239 3198
rect 9929 3152 10239 3164
rect 10359 4082 10510 4152
rect 10650 4082 10801 4152
rect 10359 4048 10461 4082
rect 10495 4048 10510 4082
rect 10650 4048 10665 4082
rect 10699 4048 10801 4082
rect 10359 4014 10510 4048
rect 10650 4014 10801 4048
rect 10359 3980 10461 4014
rect 10495 3980 10510 4014
rect 10650 3980 10665 4014
rect 10699 3980 10801 4014
rect 10359 3946 10510 3980
rect 10650 3946 10801 3980
rect 10359 3912 10461 3946
rect 10495 3912 10510 3946
rect 10650 3912 10665 3946
rect 10699 3912 10801 3946
rect 10359 3878 10510 3912
rect 10650 3878 10801 3912
rect 10359 3844 10461 3878
rect 10495 3844 10510 3878
rect 10650 3844 10665 3878
rect 10699 3844 10801 3878
rect 10359 3810 10510 3844
rect 10650 3810 10801 3844
rect 10359 3776 10461 3810
rect 10495 3776 10510 3810
rect 10650 3776 10665 3810
rect 10699 3776 10801 3810
rect 10359 3742 10510 3776
rect 10650 3742 10801 3776
rect 10359 3708 10461 3742
rect 10495 3708 10510 3742
rect 10650 3708 10665 3742
rect 10699 3708 10801 3742
rect 10359 3674 10510 3708
rect 10650 3674 10801 3708
rect 10359 3640 10461 3674
rect 10495 3640 10510 3674
rect 10650 3640 10665 3674
rect 10699 3640 10801 3674
rect 10359 3606 10510 3640
rect 10650 3606 10801 3640
rect 10359 3572 10461 3606
rect 10495 3572 10510 3606
rect 10650 3572 10665 3606
rect 10699 3572 10801 3606
rect 10359 3538 10510 3572
rect 10650 3538 10801 3572
rect 10359 3504 10461 3538
rect 10495 3504 10510 3538
rect 10650 3504 10665 3538
rect 10699 3504 10801 3538
rect 10359 3470 10510 3504
rect 10650 3470 10801 3504
rect 10359 3436 10461 3470
rect 10495 3436 10510 3470
rect 10650 3436 10665 3470
rect 10699 3436 10801 3470
rect 10359 3402 10510 3436
rect 10650 3402 10801 3436
rect 10359 3368 10461 3402
rect 10495 3368 10510 3402
rect 10650 3368 10665 3402
rect 10699 3368 10801 3402
rect 10359 3334 10510 3368
rect 10650 3334 10801 3368
rect 10359 3300 10461 3334
rect 10495 3300 10510 3334
rect 10650 3300 10665 3334
rect 10699 3300 10801 3334
rect 10359 3266 10510 3300
rect 10650 3266 10801 3300
rect 10359 3232 10461 3266
rect 10495 3232 10510 3266
rect 10650 3232 10665 3266
rect 10699 3232 10801 3266
rect 10359 3198 10510 3232
rect 10650 3198 10801 3232
rect 10359 3164 10461 3198
rect 10495 3164 10510 3198
rect 10650 3164 10665 3198
rect 10699 3164 10801 3198
rect 10359 3152 10510 3164
rect 10650 3152 10801 3164
rect 10921 4082 11231 4152
rect 10921 4048 11023 4082
rect 11057 4048 11095 4082
rect 11129 4048 11231 4082
rect 10921 4014 11231 4048
rect 10921 3980 11023 4014
rect 11057 3980 11095 4014
rect 11129 3980 11231 4014
rect 10921 3946 11231 3980
rect 10921 3912 11023 3946
rect 11057 3912 11095 3946
rect 11129 3912 11231 3946
rect 10921 3878 11231 3912
rect 10921 3844 11023 3878
rect 11057 3844 11095 3878
rect 11129 3844 11231 3878
rect 10921 3810 11231 3844
rect 10921 3776 11023 3810
rect 11057 3776 11095 3810
rect 11129 3776 11231 3810
rect 10921 3742 11231 3776
rect 10921 3708 11023 3742
rect 11057 3708 11095 3742
rect 11129 3708 11231 3742
rect 10921 3674 11231 3708
rect 10921 3640 11023 3674
rect 11057 3640 11095 3674
rect 11129 3640 11231 3674
rect 10921 3606 11231 3640
rect 10921 3572 11023 3606
rect 11057 3572 11095 3606
rect 11129 3572 11231 3606
rect 10921 3538 11231 3572
rect 10921 3504 11023 3538
rect 11057 3504 11095 3538
rect 11129 3504 11231 3538
rect 10921 3470 11231 3504
rect 10921 3436 11023 3470
rect 11057 3436 11095 3470
rect 11129 3436 11231 3470
rect 10921 3402 11231 3436
rect 10921 3368 11023 3402
rect 11057 3368 11095 3402
rect 11129 3368 11231 3402
rect 10921 3334 11231 3368
rect 10921 3300 11023 3334
rect 11057 3300 11095 3334
rect 11129 3300 11231 3334
rect 10921 3266 11231 3300
rect 10921 3232 11023 3266
rect 11057 3232 11095 3266
rect 11129 3232 11231 3266
rect 10921 3198 11231 3232
rect 10921 3164 11023 3198
rect 11057 3164 11095 3198
rect 11129 3164 11231 3198
rect 10921 3152 11231 3164
rect 11351 4082 11502 4152
rect 11642 4082 11793 4152
rect 11351 4048 11453 4082
rect 11487 4048 11502 4082
rect 11642 4048 11657 4082
rect 11691 4048 11793 4082
rect 11351 4014 11502 4048
rect 11642 4014 11793 4048
rect 11351 3980 11453 4014
rect 11487 3980 11502 4014
rect 11642 3980 11657 4014
rect 11691 3980 11793 4014
rect 11351 3946 11502 3980
rect 11642 3946 11793 3980
rect 11351 3912 11453 3946
rect 11487 3912 11502 3946
rect 11642 3912 11657 3946
rect 11691 3912 11793 3946
rect 11351 3878 11502 3912
rect 11642 3878 11793 3912
rect 11351 3844 11453 3878
rect 11487 3844 11502 3878
rect 11642 3844 11657 3878
rect 11691 3844 11793 3878
rect 11351 3810 11502 3844
rect 11642 3810 11793 3844
rect 11351 3776 11453 3810
rect 11487 3776 11502 3810
rect 11642 3776 11657 3810
rect 11691 3776 11793 3810
rect 11351 3742 11502 3776
rect 11642 3742 11793 3776
rect 11351 3708 11453 3742
rect 11487 3708 11502 3742
rect 11642 3708 11657 3742
rect 11691 3708 11793 3742
rect 11351 3674 11502 3708
rect 11642 3674 11793 3708
rect 11351 3640 11453 3674
rect 11487 3640 11502 3674
rect 11642 3640 11657 3674
rect 11691 3640 11793 3674
rect 11351 3606 11502 3640
rect 11642 3606 11793 3640
rect 11351 3572 11453 3606
rect 11487 3572 11502 3606
rect 11642 3572 11657 3606
rect 11691 3572 11793 3606
rect 11351 3538 11502 3572
rect 11642 3538 11793 3572
rect 11351 3504 11453 3538
rect 11487 3504 11502 3538
rect 11642 3504 11657 3538
rect 11691 3504 11793 3538
rect 11351 3470 11502 3504
rect 11642 3470 11793 3504
rect 11351 3436 11453 3470
rect 11487 3436 11502 3470
rect 11642 3436 11657 3470
rect 11691 3436 11793 3470
rect 11351 3402 11502 3436
rect 11642 3402 11793 3436
rect 11351 3368 11453 3402
rect 11487 3368 11502 3402
rect 11642 3368 11657 3402
rect 11691 3368 11793 3402
rect 11351 3334 11502 3368
rect 11642 3334 11793 3368
rect 11351 3300 11453 3334
rect 11487 3300 11502 3334
rect 11642 3300 11657 3334
rect 11691 3300 11793 3334
rect 11351 3266 11502 3300
rect 11642 3266 11793 3300
rect 11351 3232 11453 3266
rect 11487 3232 11502 3266
rect 11642 3232 11657 3266
rect 11691 3232 11793 3266
rect 11351 3198 11502 3232
rect 11642 3198 11793 3232
rect 11351 3164 11453 3198
rect 11487 3164 11502 3198
rect 11642 3164 11657 3198
rect 11691 3164 11793 3198
rect 11351 3152 11502 3164
rect 11642 3152 11793 3164
rect 11913 4082 12223 4152
rect 11913 4048 12015 4082
rect 12049 4048 12087 4082
rect 12121 4048 12223 4082
rect 11913 4014 12223 4048
rect 11913 3980 12015 4014
rect 12049 3980 12087 4014
rect 12121 3980 12223 4014
rect 11913 3946 12223 3980
rect 11913 3912 12015 3946
rect 12049 3912 12087 3946
rect 12121 3912 12223 3946
rect 11913 3878 12223 3912
rect 11913 3844 12015 3878
rect 12049 3844 12087 3878
rect 12121 3844 12223 3878
rect 11913 3810 12223 3844
rect 11913 3776 12015 3810
rect 12049 3776 12087 3810
rect 12121 3776 12223 3810
rect 11913 3742 12223 3776
rect 11913 3708 12015 3742
rect 12049 3708 12087 3742
rect 12121 3708 12223 3742
rect 11913 3674 12223 3708
rect 11913 3640 12015 3674
rect 12049 3640 12087 3674
rect 12121 3640 12223 3674
rect 11913 3606 12223 3640
rect 11913 3572 12015 3606
rect 12049 3572 12087 3606
rect 12121 3572 12223 3606
rect 11913 3538 12223 3572
rect 11913 3504 12015 3538
rect 12049 3504 12087 3538
rect 12121 3504 12223 3538
rect 11913 3470 12223 3504
rect 11913 3436 12015 3470
rect 12049 3436 12087 3470
rect 12121 3436 12223 3470
rect 11913 3402 12223 3436
rect 11913 3368 12015 3402
rect 12049 3368 12087 3402
rect 12121 3368 12223 3402
rect 11913 3334 12223 3368
rect 11913 3300 12015 3334
rect 12049 3300 12087 3334
rect 12121 3300 12223 3334
rect 11913 3266 12223 3300
rect 11913 3232 12015 3266
rect 12049 3232 12087 3266
rect 12121 3232 12223 3266
rect 11913 3198 12223 3232
rect 11913 3164 12015 3198
rect 12049 3164 12087 3198
rect 12121 3164 12223 3198
rect 11913 3152 12223 3164
rect 12343 4082 12494 4152
rect 12634 4082 12785 4152
rect 12343 4048 12445 4082
rect 12479 4048 12494 4082
rect 12634 4048 12649 4082
rect 12683 4048 12785 4082
rect 12343 4014 12494 4048
rect 12634 4014 12785 4048
rect 12343 3980 12445 4014
rect 12479 3980 12494 4014
rect 12634 3980 12649 4014
rect 12683 3980 12785 4014
rect 12343 3946 12494 3980
rect 12634 3946 12785 3980
rect 12343 3912 12445 3946
rect 12479 3912 12494 3946
rect 12634 3912 12649 3946
rect 12683 3912 12785 3946
rect 12343 3878 12494 3912
rect 12634 3878 12785 3912
rect 12343 3844 12445 3878
rect 12479 3844 12494 3878
rect 12634 3844 12649 3878
rect 12683 3844 12785 3878
rect 12343 3810 12494 3844
rect 12634 3810 12785 3844
rect 12343 3776 12445 3810
rect 12479 3776 12494 3810
rect 12634 3776 12649 3810
rect 12683 3776 12785 3810
rect 12343 3742 12494 3776
rect 12634 3742 12785 3776
rect 12343 3708 12445 3742
rect 12479 3708 12494 3742
rect 12634 3708 12649 3742
rect 12683 3708 12785 3742
rect 12343 3674 12494 3708
rect 12634 3674 12785 3708
rect 12343 3640 12445 3674
rect 12479 3640 12494 3674
rect 12634 3640 12649 3674
rect 12683 3640 12785 3674
rect 12343 3606 12494 3640
rect 12634 3606 12785 3640
rect 12343 3572 12445 3606
rect 12479 3572 12494 3606
rect 12634 3572 12649 3606
rect 12683 3572 12785 3606
rect 12343 3538 12494 3572
rect 12634 3538 12785 3572
rect 12343 3504 12445 3538
rect 12479 3504 12494 3538
rect 12634 3504 12649 3538
rect 12683 3504 12785 3538
rect 12343 3470 12494 3504
rect 12634 3470 12785 3504
rect 12343 3436 12445 3470
rect 12479 3436 12494 3470
rect 12634 3436 12649 3470
rect 12683 3436 12785 3470
rect 12343 3402 12494 3436
rect 12634 3402 12785 3436
rect 12343 3368 12445 3402
rect 12479 3368 12494 3402
rect 12634 3368 12649 3402
rect 12683 3368 12785 3402
rect 12343 3334 12494 3368
rect 12634 3334 12785 3368
rect 12343 3300 12445 3334
rect 12479 3300 12494 3334
rect 12634 3300 12649 3334
rect 12683 3300 12785 3334
rect 12343 3266 12494 3300
rect 12634 3266 12785 3300
rect 12343 3232 12445 3266
rect 12479 3232 12494 3266
rect 12634 3232 12649 3266
rect 12683 3232 12785 3266
rect 12343 3198 12494 3232
rect 12634 3198 12785 3232
rect 12343 3164 12445 3198
rect 12479 3164 12494 3198
rect 12634 3164 12649 3198
rect 12683 3164 12785 3198
rect 12343 3152 12494 3164
rect 12634 3152 12785 3164
rect 12905 4082 13215 4152
rect 12905 4048 13007 4082
rect 13041 4048 13079 4082
rect 13113 4048 13215 4082
rect 12905 4014 13215 4048
rect 12905 3980 13007 4014
rect 13041 3980 13079 4014
rect 13113 3980 13215 4014
rect 12905 3946 13215 3980
rect 12905 3912 13007 3946
rect 13041 3912 13079 3946
rect 13113 3912 13215 3946
rect 12905 3878 13215 3912
rect 12905 3844 13007 3878
rect 13041 3844 13079 3878
rect 13113 3844 13215 3878
rect 12905 3810 13215 3844
rect 12905 3776 13007 3810
rect 13041 3776 13079 3810
rect 13113 3776 13215 3810
rect 12905 3742 13215 3776
rect 12905 3708 13007 3742
rect 13041 3708 13079 3742
rect 13113 3708 13215 3742
rect 12905 3674 13215 3708
rect 12905 3640 13007 3674
rect 13041 3640 13079 3674
rect 13113 3640 13215 3674
rect 12905 3606 13215 3640
rect 12905 3572 13007 3606
rect 13041 3572 13079 3606
rect 13113 3572 13215 3606
rect 12905 3538 13215 3572
rect 12905 3504 13007 3538
rect 13041 3504 13079 3538
rect 13113 3504 13215 3538
rect 12905 3470 13215 3504
rect 12905 3436 13007 3470
rect 13041 3436 13079 3470
rect 13113 3436 13215 3470
rect 12905 3402 13215 3436
rect 12905 3368 13007 3402
rect 13041 3368 13079 3402
rect 13113 3368 13215 3402
rect 12905 3334 13215 3368
rect 12905 3300 13007 3334
rect 13041 3300 13079 3334
rect 13113 3300 13215 3334
rect 12905 3266 13215 3300
rect 12905 3232 13007 3266
rect 13041 3232 13079 3266
rect 13113 3232 13215 3266
rect 12905 3198 13215 3232
rect 12905 3164 13007 3198
rect 13041 3164 13079 3198
rect 13113 3164 13215 3198
rect 12905 3152 13215 3164
rect 13335 4082 13486 4152
rect 13626 4082 13777 4152
rect 13335 4048 13437 4082
rect 13471 4048 13486 4082
rect 13626 4048 13641 4082
rect 13675 4048 13777 4082
rect 13335 4014 13486 4048
rect 13626 4014 13777 4048
rect 13335 3980 13437 4014
rect 13471 3980 13486 4014
rect 13626 3980 13641 4014
rect 13675 3980 13777 4014
rect 13335 3946 13486 3980
rect 13626 3946 13777 3980
rect 13335 3912 13437 3946
rect 13471 3912 13486 3946
rect 13626 3912 13641 3946
rect 13675 3912 13777 3946
rect 13335 3878 13486 3912
rect 13626 3878 13777 3912
rect 13335 3844 13437 3878
rect 13471 3844 13486 3878
rect 13626 3844 13641 3878
rect 13675 3844 13777 3878
rect 13335 3810 13486 3844
rect 13626 3810 13777 3844
rect 13335 3776 13437 3810
rect 13471 3776 13486 3810
rect 13626 3776 13641 3810
rect 13675 3776 13777 3810
rect 13335 3742 13486 3776
rect 13626 3742 13777 3776
rect 13335 3708 13437 3742
rect 13471 3708 13486 3742
rect 13626 3708 13641 3742
rect 13675 3708 13777 3742
rect 13335 3674 13486 3708
rect 13626 3674 13777 3708
rect 13335 3640 13437 3674
rect 13471 3640 13486 3674
rect 13626 3640 13641 3674
rect 13675 3640 13777 3674
rect 13335 3606 13486 3640
rect 13626 3606 13777 3640
rect 13335 3572 13437 3606
rect 13471 3572 13486 3606
rect 13626 3572 13641 3606
rect 13675 3572 13777 3606
rect 13335 3538 13486 3572
rect 13626 3538 13777 3572
rect 13335 3504 13437 3538
rect 13471 3504 13486 3538
rect 13626 3504 13641 3538
rect 13675 3504 13777 3538
rect 13335 3470 13486 3504
rect 13626 3470 13777 3504
rect 13335 3436 13437 3470
rect 13471 3436 13486 3470
rect 13626 3436 13641 3470
rect 13675 3436 13777 3470
rect 13335 3402 13486 3436
rect 13626 3402 13777 3436
rect 13335 3368 13437 3402
rect 13471 3368 13486 3402
rect 13626 3368 13641 3402
rect 13675 3368 13777 3402
rect 13335 3334 13486 3368
rect 13626 3334 13777 3368
rect 13335 3300 13437 3334
rect 13471 3300 13486 3334
rect 13626 3300 13641 3334
rect 13675 3300 13777 3334
rect 13335 3266 13486 3300
rect 13626 3266 13777 3300
rect 13335 3232 13437 3266
rect 13471 3232 13486 3266
rect 13626 3232 13641 3266
rect 13675 3232 13777 3266
rect 13335 3198 13486 3232
rect 13626 3198 13777 3232
rect 13335 3164 13437 3198
rect 13471 3164 13486 3198
rect 13626 3164 13641 3198
rect 13675 3164 13777 3198
rect 13335 3152 13486 3164
rect 13626 3152 13777 3164
rect 13897 4082 14135 4152
rect 13897 4048 13999 4082
rect 14033 4048 14135 4082
rect 13897 4014 14135 4048
rect 13897 3980 13999 4014
rect 14033 3980 14135 4014
rect 13897 3946 14135 3980
rect 13897 3912 13999 3946
rect 14033 3912 14135 3946
rect 13897 3878 14135 3912
rect 13897 3844 13999 3878
rect 14033 3844 14135 3878
rect 13897 3810 14135 3844
rect 13897 3776 13999 3810
rect 14033 3776 14135 3810
rect 13897 3742 14135 3776
rect 13897 3708 13999 3742
rect 14033 3708 14135 3742
rect 13897 3674 14135 3708
rect 13897 3640 13999 3674
rect 14033 3640 14135 3674
rect 13897 3606 14135 3640
rect 13897 3572 13999 3606
rect 14033 3572 14135 3606
rect 13897 3538 14135 3572
rect 13897 3504 13999 3538
rect 14033 3504 14135 3538
rect 13897 3470 14135 3504
rect 13897 3436 13999 3470
rect 14033 3436 14135 3470
rect 13897 3402 14135 3436
rect 13897 3368 13999 3402
rect 14033 3368 14135 3402
rect 13897 3334 14135 3368
rect 13897 3300 13999 3334
rect 14033 3300 14135 3334
rect 13897 3266 14135 3300
rect 13897 3232 13999 3266
rect 14033 3232 14135 3266
rect 13897 3198 14135 3232
rect 13897 3164 13999 3198
rect 14033 3164 14135 3198
rect 13897 3152 14135 3164
rect 14255 4082 14427 4152
rect 14255 4048 14356 4082
rect 14390 4048 14427 4082
rect 14255 4014 14427 4048
rect 14255 3980 14356 4014
rect 14390 3980 14427 4014
rect 14255 3946 14427 3980
rect 14255 3912 14356 3946
rect 14390 3912 14427 3946
rect 14255 3878 14427 3912
rect 14255 3844 14356 3878
rect 14390 3844 14427 3878
rect 14255 3810 14427 3844
rect 14255 3776 14356 3810
rect 14390 3776 14427 3810
rect 14255 3742 14427 3776
rect 14255 3708 14356 3742
rect 14390 3708 14427 3742
rect 14255 3674 14427 3708
rect 14255 3640 14356 3674
rect 14390 3640 14427 3674
rect 14255 3606 14427 3640
rect 14255 3572 14356 3606
rect 14390 3572 14427 3606
rect 14255 3538 14427 3572
rect 14255 3504 14356 3538
rect 14390 3504 14427 3538
rect 14255 3470 14427 3504
rect 14255 3436 14356 3470
rect 14390 3436 14427 3470
rect 14255 3402 14427 3436
rect 14255 3368 14356 3402
rect 14390 3368 14427 3402
rect 14255 3334 14427 3368
rect 14255 3300 14356 3334
rect 14390 3300 14427 3334
rect 14255 3266 14427 3300
rect 14255 3232 14356 3266
rect 14390 3232 14427 3266
rect 14255 3198 14427 3232
rect 14255 3164 14356 3198
rect 14390 3164 14427 3198
rect 14255 3152 14427 3164
rect 708 2482 881 2552
rect 708 2448 745 2482
rect 779 2448 881 2482
rect 708 2414 881 2448
rect 708 2380 745 2414
rect 779 2380 881 2414
rect 708 2346 881 2380
rect 708 2312 745 2346
rect 779 2312 881 2346
rect 708 2278 881 2312
rect 708 2244 745 2278
rect 779 2244 881 2278
rect 708 2210 881 2244
rect 708 2176 745 2210
rect 779 2176 881 2210
rect 708 2142 881 2176
rect 708 2108 745 2142
rect 779 2108 881 2142
rect 708 2074 881 2108
rect 708 2040 745 2074
rect 779 2040 881 2074
rect 708 2006 881 2040
rect 708 1972 745 2006
rect 779 1972 881 2006
rect 708 1938 881 1972
rect 708 1904 745 1938
rect 779 1904 881 1938
rect 708 1870 881 1904
rect 708 1836 745 1870
rect 779 1836 881 1870
rect 708 1802 881 1836
rect 708 1768 745 1802
rect 779 1768 881 1802
rect 708 1734 881 1768
rect 708 1700 745 1734
rect 779 1700 881 1734
rect 708 1666 881 1700
rect 708 1632 745 1666
rect 779 1632 881 1666
rect 708 1598 881 1632
rect 708 1564 745 1598
rect 779 1564 881 1598
rect 708 1552 881 1564
rect 1001 2482 1311 2552
rect 1001 2448 1103 2482
rect 1137 2448 1175 2482
rect 1209 2448 1311 2482
rect 1001 2414 1311 2448
rect 1001 2380 1103 2414
rect 1137 2380 1175 2414
rect 1209 2380 1311 2414
rect 1001 2346 1311 2380
rect 1001 2312 1103 2346
rect 1137 2312 1175 2346
rect 1209 2312 1311 2346
rect 1001 2278 1311 2312
rect 1001 2244 1103 2278
rect 1137 2244 1175 2278
rect 1209 2244 1311 2278
rect 1001 2210 1311 2244
rect 1001 2176 1103 2210
rect 1137 2176 1175 2210
rect 1209 2176 1311 2210
rect 1001 2142 1311 2176
rect 1001 2108 1103 2142
rect 1137 2108 1175 2142
rect 1209 2108 1311 2142
rect 1001 2074 1311 2108
rect 1001 2040 1103 2074
rect 1137 2040 1175 2074
rect 1209 2040 1311 2074
rect 1001 2006 1311 2040
rect 1001 1972 1103 2006
rect 1137 1972 1175 2006
rect 1209 1972 1311 2006
rect 1001 1938 1311 1972
rect 1001 1904 1103 1938
rect 1137 1904 1175 1938
rect 1209 1904 1311 1938
rect 1001 1870 1311 1904
rect 1001 1836 1103 1870
rect 1137 1836 1175 1870
rect 1209 1836 1311 1870
rect 1001 1802 1311 1836
rect 1001 1768 1103 1802
rect 1137 1768 1175 1802
rect 1209 1768 1311 1802
rect 1001 1734 1311 1768
rect 1001 1700 1103 1734
rect 1137 1700 1175 1734
rect 1209 1700 1311 1734
rect 1001 1666 1311 1700
rect 1001 1632 1103 1666
rect 1137 1632 1175 1666
rect 1209 1632 1311 1666
rect 1001 1598 1311 1632
rect 1001 1564 1103 1598
rect 1137 1564 1175 1598
rect 1209 1564 1311 1598
rect 1001 1552 1311 1564
rect 1431 2540 1582 2552
rect 1722 2540 1873 2552
rect 1431 2506 1533 2540
rect 1567 2506 1582 2540
rect 1722 2506 1737 2540
rect 1771 2506 1873 2540
rect 1431 2472 1582 2506
rect 1722 2472 1873 2506
rect 1431 2438 1533 2472
rect 1567 2438 1582 2472
rect 1722 2438 1737 2472
rect 1771 2438 1873 2472
rect 1431 2404 1582 2438
rect 1722 2404 1873 2438
rect 1431 2370 1533 2404
rect 1567 2370 1582 2404
rect 1722 2370 1737 2404
rect 1771 2370 1873 2404
rect 1431 2336 1582 2370
rect 1722 2336 1873 2370
rect 1431 2302 1533 2336
rect 1567 2302 1582 2336
rect 1722 2302 1737 2336
rect 1771 2302 1873 2336
rect 1431 2268 1582 2302
rect 1722 2268 1873 2302
rect 1431 2234 1533 2268
rect 1567 2234 1582 2268
rect 1722 2234 1737 2268
rect 1771 2234 1873 2268
rect 1431 2200 1582 2234
rect 1722 2200 1873 2234
rect 1431 2166 1533 2200
rect 1567 2166 1582 2200
rect 1722 2166 1737 2200
rect 1771 2166 1873 2200
rect 1431 2132 1582 2166
rect 1722 2132 1873 2166
rect 1431 2098 1533 2132
rect 1567 2098 1582 2132
rect 1722 2098 1737 2132
rect 1771 2098 1873 2132
rect 1431 2064 1582 2098
rect 1722 2064 1873 2098
rect 1431 2030 1533 2064
rect 1567 2030 1582 2064
rect 1722 2030 1737 2064
rect 1771 2030 1873 2064
rect 1431 1996 1582 2030
rect 1722 1996 1873 2030
rect 1431 1962 1533 1996
rect 1567 1962 1582 1996
rect 1722 1962 1737 1996
rect 1771 1962 1873 1996
rect 1431 1928 1582 1962
rect 1722 1928 1873 1962
rect 1431 1894 1533 1928
rect 1567 1894 1582 1928
rect 1722 1894 1737 1928
rect 1771 1894 1873 1928
rect 1431 1860 1582 1894
rect 1722 1860 1873 1894
rect 1431 1826 1533 1860
rect 1567 1826 1582 1860
rect 1722 1826 1737 1860
rect 1771 1826 1873 1860
rect 1431 1792 1582 1826
rect 1722 1792 1873 1826
rect 1431 1758 1533 1792
rect 1567 1758 1582 1792
rect 1722 1758 1737 1792
rect 1771 1758 1873 1792
rect 1431 1724 1582 1758
rect 1722 1724 1873 1758
rect 1431 1690 1533 1724
rect 1567 1690 1582 1724
rect 1722 1690 1737 1724
rect 1771 1690 1873 1724
rect 1431 1656 1582 1690
rect 1722 1656 1873 1690
rect 1431 1622 1533 1656
rect 1567 1622 1582 1656
rect 1722 1622 1737 1656
rect 1771 1622 1873 1656
rect 1431 1552 1582 1622
rect 1722 1552 1873 1622
rect 1993 2482 2303 2552
rect 1993 2448 2095 2482
rect 2129 2448 2167 2482
rect 2201 2448 2303 2482
rect 1993 2414 2303 2448
rect 1993 2380 2095 2414
rect 2129 2380 2167 2414
rect 2201 2380 2303 2414
rect 1993 2346 2303 2380
rect 1993 2312 2095 2346
rect 2129 2312 2167 2346
rect 2201 2312 2303 2346
rect 1993 2278 2303 2312
rect 1993 2244 2095 2278
rect 2129 2244 2167 2278
rect 2201 2244 2303 2278
rect 1993 2210 2303 2244
rect 1993 2176 2095 2210
rect 2129 2176 2167 2210
rect 2201 2176 2303 2210
rect 1993 2142 2303 2176
rect 1993 2108 2095 2142
rect 2129 2108 2167 2142
rect 2201 2108 2303 2142
rect 1993 2074 2303 2108
rect 1993 2040 2095 2074
rect 2129 2040 2167 2074
rect 2201 2040 2303 2074
rect 1993 2006 2303 2040
rect 1993 1972 2095 2006
rect 2129 1972 2167 2006
rect 2201 1972 2303 2006
rect 1993 1938 2303 1972
rect 1993 1904 2095 1938
rect 2129 1904 2167 1938
rect 2201 1904 2303 1938
rect 1993 1870 2303 1904
rect 1993 1836 2095 1870
rect 2129 1836 2167 1870
rect 2201 1836 2303 1870
rect 1993 1802 2303 1836
rect 1993 1768 2095 1802
rect 2129 1768 2167 1802
rect 2201 1768 2303 1802
rect 1993 1734 2303 1768
rect 1993 1700 2095 1734
rect 2129 1700 2167 1734
rect 2201 1700 2303 1734
rect 1993 1666 2303 1700
rect 1993 1632 2095 1666
rect 2129 1632 2167 1666
rect 2201 1632 2303 1666
rect 1993 1598 2303 1632
rect 1993 1564 2095 1598
rect 2129 1564 2167 1598
rect 2201 1564 2303 1598
rect 1993 1552 2303 1564
rect 2423 2540 2574 2552
rect 2714 2540 2865 2552
rect 2423 2506 2525 2540
rect 2559 2506 2574 2540
rect 2714 2506 2729 2540
rect 2763 2506 2865 2540
rect 2423 2472 2574 2506
rect 2714 2472 2865 2506
rect 2423 2438 2525 2472
rect 2559 2438 2574 2472
rect 2714 2438 2729 2472
rect 2763 2438 2865 2472
rect 2423 2404 2574 2438
rect 2714 2404 2865 2438
rect 2423 2370 2525 2404
rect 2559 2370 2574 2404
rect 2714 2370 2729 2404
rect 2763 2370 2865 2404
rect 2423 2336 2574 2370
rect 2714 2336 2865 2370
rect 2423 2302 2525 2336
rect 2559 2302 2574 2336
rect 2714 2302 2729 2336
rect 2763 2302 2865 2336
rect 2423 2268 2574 2302
rect 2714 2268 2865 2302
rect 2423 2234 2525 2268
rect 2559 2234 2574 2268
rect 2714 2234 2729 2268
rect 2763 2234 2865 2268
rect 2423 2200 2574 2234
rect 2714 2200 2865 2234
rect 2423 2166 2525 2200
rect 2559 2166 2574 2200
rect 2714 2166 2729 2200
rect 2763 2166 2865 2200
rect 2423 2132 2574 2166
rect 2714 2132 2865 2166
rect 2423 2098 2525 2132
rect 2559 2098 2574 2132
rect 2714 2098 2729 2132
rect 2763 2098 2865 2132
rect 2423 2064 2574 2098
rect 2714 2064 2865 2098
rect 2423 2030 2525 2064
rect 2559 2030 2574 2064
rect 2714 2030 2729 2064
rect 2763 2030 2865 2064
rect 2423 1996 2574 2030
rect 2714 1996 2865 2030
rect 2423 1962 2525 1996
rect 2559 1962 2574 1996
rect 2714 1962 2729 1996
rect 2763 1962 2865 1996
rect 2423 1928 2574 1962
rect 2714 1928 2865 1962
rect 2423 1894 2525 1928
rect 2559 1894 2574 1928
rect 2714 1894 2729 1928
rect 2763 1894 2865 1928
rect 2423 1860 2574 1894
rect 2714 1860 2865 1894
rect 2423 1826 2525 1860
rect 2559 1826 2574 1860
rect 2714 1826 2729 1860
rect 2763 1826 2865 1860
rect 2423 1792 2574 1826
rect 2714 1792 2865 1826
rect 2423 1758 2525 1792
rect 2559 1758 2574 1792
rect 2714 1758 2729 1792
rect 2763 1758 2865 1792
rect 2423 1724 2574 1758
rect 2714 1724 2865 1758
rect 2423 1690 2525 1724
rect 2559 1690 2574 1724
rect 2714 1690 2729 1724
rect 2763 1690 2865 1724
rect 2423 1656 2574 1690
rect 2714 1656 2865 1690
rect 2423 1622 2525 1656
rect 2559 1622 2574 1656
rect 2714 1622 2729 1656
rect 2763 1622 2865 1656
rect 2423 1552 2574 1622
rect 2714 1552 2865 1622
rect 2985 2482 3295 2552
rect 2985 2448 3087 2482
rect 3121 2448 3159 2482
rect 3193 2448 3295 2482
rect 2985 2414 3295 2448
rect 2985 2380 3087 2414
rect 3121 2380 3159 2414
rect 3193 2380 3295 2414
rect 2985 2346 3295 2380
rect 2985 2312 3087 2346
rect 3121 2312 3159 2346
rect 3193 2312 3295 2346
rect 2985 2278 3295 2312
rect 2985 2244 3087 2278
rect 3121 2244 3159 2278
rect 3193 2244 3295 2278
rect 2985 2210 3295 2244
rect 2985 2176 3087 2210
rect 3121 2176 3159 2210
rect 3193 2176 3295 2210
rect 2985 2142 3295 2176
rect 2985 2108 3087 2142
rect 3121 2108 3159 2142
rect 3193 2108 3295 2142
rect 2985 2074 3295 2108
rect 2985 2040 3087 2074
rect 3121 2040 3159 2074
rect 3193 2040 3295 2074
rect 2985 2006 3295 2040
rect 2985 1972 3087 2006
rect 3121 1972 3159 2006
rect 3193 1972 3295 2006
rect 2985 1938 3295 1972
rect 2985 1904 3087 1938
rect 3121 1904 3159 1938
rect 3193 1904 3295 1938
rect 2985 1870 3295 1904
rect 2985 1836 3087 1870
rect 3121 1836 3159 1870
rect 3193 1836 3295 1870
rect 2985 1802 3295 1836
rect 2985 1768 3087 1802
rect 3121 1768 3159 1802
rect 3193 1768 3295 1802
rect 2985 1734 3295 1768
rect 2985 1700 3087 1734
rect 3121 1700 3159 1734
rect 3193 1700 3295 1734
rect 2985 1666 3295 1700
rect 2985 1632 3087 1666
rect 3121 1632 3159 1666
rect 3193 1632 3295 1666
rect 2985 1598 3295 1632
rect 2985 1564 3087 1598
rect 3121 1564 3159 1598
rect 3193 1564 3295 1598
rect 2985 1552 3295 1564
rect 3415 2540 3566 2552
rect 3706 2540 3857 2552
rect 3415 2506 3517 2540
rect 3551 2506 3566 2540
rect 3706 2506 3721 2540
rect 3755 2506 3857 2540
rect 3415 2472 3566 2506
rect 3706 2472 3857 2506
rect 3415 2438 3517 2472
rect 3551 2438 3566 2472
rect 3706 2438 3721 2472
rect 3755 2438 3857 2472
rect 3415 2404 3566 2438
rect 3706 2404 3857 2438
rect 3415 2370 3517 2404
rect 3551 2370 3566 2404
rect 3706 2370 3721 2404
rect 3755 2370 3857 2404
rect 3415 2336 3566 2370
rect 3706 2336 3857 2370
rect 3415 2302 3517 2336
rect 3551 2302 3566 2336
rect 3706 2302 3721 2336
rect 3755 2302 3857 2336
rect 3415 2268 3566 2302
rect 3706 2268 3857 2302
rect 3415 2234 3517 2268
rect 3551 2234 3566 2268
rect 3706 2234 3721 2268
rect 3755 2234 3857 2268
rect 3415 2200 3566 2234
rect 3706 2200 3857 2234
rect 3415 2166 3517 2200
rect 3551 2166 3566 2200
rect 3706 2166 3721 2200
rect 3755 2166 3857 2200
rect 3415 2132 3566 2166
rect 3706 2132 3857 2166
rect 3415 2098 3517 2132
rect 3551 2098 3566 2132
rect 3706 2098 3721 2132
rect 3755 2098 3857 2132
rect 3415 2064 3566 2098
rect 3706 2064 3857 2098
rect 3415 2030 3517 2064
rect 3551 2030 3566 2064
rect 3706 2030 3721 2064
rect 3755 2030 3857 2064
rect 3415 1996 3566 2030
rect 3706 1996 3857 2030
rect 3415 1962 3517 1996
rect 3551 1962 3566 1996
rect 3706 1962 3721 1996
rect 3755 1962 3857 1996
rect 3415 1928 3566 1962
rect 3706 1928 3857 1962
rect 3415 1894 3517 1928
rect 3551 1894 3566 1928
rect 3706 1894 3721 1928
rect 3755 1894 3857 1928
rect 3415 1860 3566 1894
rect 3706 1860 3857 1894
rect 3415 1826 3517 1860
rect 3551 1826 3566 1860
rect 3706 1826 3721 1860
rect 3755 1826 3857 1860
rect 3415 1792 3566 1826
rect 3706 1792 3857 1826
rect 3415 1758 3517 1792
rect 3551 1758 3566 1792
rect 3706 1758 3721 1792
rect 3755 1758 3857 1792
rect 3415 1724 3566 1758
rect 3706 1724 3857 1758
rect 3415 1690 3517 1724
rect 3551 1690 3566 1724
rect 3706 1690 3721 1724
rect 3755 1690 3857 1724
rect 3415 1656 3566 1690
rect 3706 1656 3857 1690
rect 3415 1622 3517 1656
rect 3551 1622 3566 1656
rect 3706 1622 3721 1656
rect 3755 1622 3857 1656
rect 3415 1552 3566 1622
rect 3706 1552 3857 1622
rect 3977 2482 4287 2552
rect 3977 2448 4079 2482
rect 4113 2448 4151 2482
rect 4185 2448 4287 2482
rect 3977 2414 4287 2448
rect 3977 2380 4079 2414
rect 4113 2380 4151 2414
rect 4185 2380 4287 2414
rect 3977 2346 4287 2380
rect 3977 2312 4079 2346
rect 4113 2312 4151 2346
rect 4185 2312 4287 2346
rect 3977 2278 4287 2312
rect 3977 2244 4079 2278
rect 4113 2244 4151 2278
rect 4185 2244 4287 2278
rect 3977 2210 4287 2244
rect 3977 2176 4079 2210
rect 4113 2176 4151 2210
rect 4185 2176 4287 2210
rect 3977 2142 4287 2176
rect 3977 2108 4079 2142
rect 4113 2108 4151 2142
rect 4185 2108 4287 2142
rect 3977 2074 4287 2108
rect 3977 2040 4079 2074
rect 4113 2040 4151 2074
rect 4185 2040 4287 2074
rect 3977 2006 4287 2040
rect 3977 1972 4079 2006
rect 4113 1972 4151 2006
rect 4185 1972 4287 2006
rect 3977 1938 4287 1972
rect 3977 1904 4079 1938
rect 4113 1904 4151 1938
rect 4185 1904 4287 1938
rect 3977 1870 4287 1904
rect 3977 1836 4079 1870
rect 4113 1836 4151 1870
rect 4185 1836 4287 1870
rect 3977 1802 4287 1836
rect 3977 1768 4079 1802
rect 4113 1768 4151 1802
rect 4185 1768 4287 1802
rect 3977 1734 4287 1768
rect 3977 1700 4079 1734
rect 4113 1700 4151 1734
rect 4185 1700 4287 1734
rect 3977 1666 4287 1700
rect 3977 1632 4079 1666
rect 4113 1632 4151 1666
rect 4185 1632 4287 1666
rect 3977 1598 4287 1632
rect 3977 1564 4079 1598
rect 4113 1564 4151 1598
rect 4185 1564 4287 1598
rect 3977 1552 4287 1564
rect 4407 2540 4558 2552
rect 4698 2540 4849 2552
rect 4407 2506 4509 2540
rect 4543 2506 4558 2540
rect 4698 2506 4713 2540
rect 4747 2506 4849 2540
rect 4407 2472 4558 2506
rect 4698 2472 4849 2506
rect 4407 2438 4509 2472
rect 4543 2438 4558 2472
rect 4698 2438 4713 2472
rect 4747 2438 4849 2472
rect 4407 2404 4558 2438
rect 4698 2404 4849 2438
rect 4407 2370 4509 2404
rect 4543 2370 4558 2404
rect 4698 2370 4713 2404
rect 4747 2370 4849 2404
rect 4407 2336 4558 2370
rect 4698 2336 4849 2370
rect 4407 2302 4509 2336
rect 4543 2302 4558 2336
rect 4698 2302 4713 2336
rect 4747 2302 4849 2336
rect 4407 2268 4558 2302
rect 4698 2268 4849 2302
rect 4407 2234 4509 2268
rect 4543 2234 4558 2268
rect 4698 2234 4713 2268
rect 4747 2234 4849 2268
rect 4407 2200 4558 2234
rect 4698 2200 4849 2234
rect 4407 2166 4509 2200
rect 4543 2166 4558 2200
rect 4698 2166 4713 2200
rect 4747 2166 4849 2200
rect 4407 2132 4558 2166
rect 4698 2132 4849 2166
rect 4407 2098 4509 2132
rect 4543 2098 4558 2132
rect 4698 2098 4713 2132
rect 4747 2098 4849 2132
rect 4407 2064 4558 2098
rect 4698 2064 4849 2098
rect 4407 2030 4509 2064
rect 4543 2030 4558 2064
rect 4698 2030 4713 2064
rect 4747 2030 4849 2064
rect 4407 1996 4558 2030
rect 4698 1996 4849 2030
rect 4407 1962 4509 1996
rect 4543 1962 4558 1996
rect 4698 1962 4713 1996
rect 4747 1962 4849 1996
rect 4407 1928 4558 1962
rect 4698 1928 4849 1962
rect 4407 1894 4509 1928
rect 4543 1894 4558 1928
rect 4698 1894 4713 1928
rect 4747 1894 4849 1928
rect 4407 1860 4558 1894
rect 4698 1860 4849 1894
rect 4407 1826 4509 1860
rect 4543 1826 4558 1860
rect 4698 1826 4713 1860
rect 4747 1826 4849 1860
rect 4407 1792 4558 1826
rect 4698 1792 4849 1826
rect 4407 1758 4509 1792
rect 4543 1758 4558 1792
rect 4698 1758 4713 1792
rect 4747 1758 4849 1792
rect 4407 1724 4558 1758
rect 4698 1724 4849 1758
rect 4407 1690 4509 1724
rect 4543 1690 4558 1724
rect 4698 1690 4713 1724
rect 4747 1690 4849 1724
rect 4407 1656 4558 1690
rect 4698 1656 4849 1690
rect 4407 1622 4509 1656
rect 4543 1622 4558 1656
rect 4698 1622 4713 1656
rect 4747 1622 4849 1656
rect 4407 1552 4558 1622
rect 4698 1552 4849 1622
rect 4969 2482 5279 2552
rect 4969 2448 5071 2482
rect 5105 2448 5143 2482
rect 5177 2448 5279 2482
rect 4969 2414 5279 2448
rect 4969 2380 5071 2414
rect 5105 2380 5143 2414
rect 5177 2380 5279 2414
rect 4969 2346 5279 2380
rect 4969 2312 5071 2346
rect 5105 2312 5143 2346
rect 5177 2312 5279 2346
rect 4969 2278 5279 2312
rect 4969 2244 5071 2278
rect 5105 2244 5143 2278
rect 5177 2244 5279 2278
rect 4969 2210 5279 2244
rect 4969 2176 5071 2210
rect 5105 2176 5143 2210
rect 5177 2176 5279 2210
rect 4969 2142 5279 2176
rect 4969 2108 5071 2142
rect 5105 2108 5143 2142
rect 5177 2108 5279 2142
rect 4969 2074 5279 2108
rect 4969 2040 5071 2074
rect 5105 2040 5143 2074
rect 5177 2040 5279 2074
rect 4969 2006 5279 2040
rect 4969 1972 5071 2006
rect 5105 1972 5143 2006
rect 5177 1972 5279 2006
rect 4969 1938 5279 1972
rect 4969 1904 5071 1938
rect 5105 1904 5143 1938
rect 5177 1904 5279 1938
rect 4969 1870 5279 1904
rect 4969 1836 5071 1870
rect 5105 1836 5143 1870
rect 5177 1836 5279 1870
rect 4969 1802 5279 1836
rect 4969 1768 5071 1802
rect 5105 1768 5143 1802
rect 5177 1768 5279 1802
rect 4969 1734 5279 1768
rect 4969 1700 5071 1734
rect 5105 1700 5143 1734
rect 5177 1700 5279 1734
rect 4969 1666 5279 1700
rect 4969 1632 5071 1666
rect 5105 1632 5143 1666
rect 5177 1632 5279 1666
rect 4969 1598 5279 1632
rect 4969 1564 5071 1598
rect 5105 1564 5143 1598
rect 5177 1564 5279 1598
rect 4969 1552 5279 1564
rect 5399 2540 5550 2552
rect 5690 2540 5841 2552
rect 5399 2506 5501 2540
rect 5535 2506 5550 2540
rect 5690 2506 5705 2540
rect 5739 2506 5841 2540
rect 5399 2472 5550 2506
rect 5690 2472 5841 2506
rect 5399 2438 5501 2472
rect 5535 2438 5550 2472
rect 5690 2438 5705 2472
rect 5739 2438 5841 2472
rect 5399 2404 5550 2438
rect 5690 2404 5841 2438
rect 5399 2370 5501 2404
rect 5535 2370 5550 2404
rect 5690 2370 5705 2404
rect 5739 2370 5841 2404
rect 5399 2336 5550 2370
rect 5690 2336 5841 2370
rect 5399 2302 5501 2336
rect 5535 2302 5550 2336
rect 5690 2302 5705 2336
rect 5739 2302 5841 2336
rect 5399 2268 5550 2302
rect 5690 2268 5841 2302
rect 5399 2234 5501 2268
rect 5535 2234 5550 2268
rect 5690 2234 5705 2268
rect 5739 2234 5841 2268
rect 5399 2200 5550 2234
rect 5690 2200 5841 2234
rect 5399 2166 5501 2200
rect 5535 2166 5550 2200
rect 5690 2166 5705 2200
rect 5739 2166 5841 2200
rect 5399 2132 5550 2166
rect 5690 2132 5841 2166
rect 5399 2098 5501 2132
rect 5535 2098 5550 2132
rect 5690 2098 5705 2132
rect 5739 2098 5841 2132
rect 5399 2064 5550 2098
rect 5690 2064 5841 2098
rect 5399 2030 5501 2064
rect 5535 2030 5550 2064
rect 5690 2030 5705 2064
rect 5739 2030 5841 2064
rect 5399 1996 5550 2030
rect 5690 1996 5841 2030
rect 5399 1962 5501 1996
rect 5535 1962 5550 1996
rect 5690 1962 5705 1996
rect 5739 1962 5841 1996
rect 5399 1928 5550 1962
rect 5690 1928 5841 1962
rect 5399 1894 5501 1928
rect 5535 1894 5550 1928
rect 5690 1894 5705 1928
rect 5739 1894 5841 1928
rect 5399 1860 5550 1894
rect 5690 1860 5841 1894
rect 5399 1826 5501 1860
rect 5535 1826 5550 1860
rect 5690 1826 5705 1860
rect 5739 1826 5841 1860
rect 5399 1792 5550 1826
rect 5690 1792 5841 1826
rect 5399 1758 5501 1792
rect 5535 1758 5550 1792
rect 5690 1758 5705 1792
rect 5739 1758 5841 1792
rect 5399 1724 5550 1758
rect 5690 1724 5841 1758
rect 5399 1690 5501 1724
rect 5535 1690 5550 1724
rect 5690 1690 5705 1724
rect 5739 1690 5841 1724
rect 5399 1656 5550 1690
rect 5690 1656 5841 1690
rect 5399 1622 5501 1656
rect 5535 1622 5550 1656
rect 5690 1622 5705 1656
rect 5739 1622 5841 1656
rect 5399 1552 5550 1622
rect 5690 1552 5841 1622
rect 5961 2482 6271 2552
rect 5961 2448 6063 2482
rect 6097 2448 6135 2482
rect 6169 2448 6271 2482
rect 5961 2414 6271 2448
rect 5961 2380 6063 2414
rect 6097 2380 6135 2414
rect 6169 2380 6271 2414
rect 5961 2346 6271 2380
rect 5961 2312 6063 2346
rect 6097 2312 6135 2346
rect 6169 2312 6271 2346
rect 5961 2278 6271 2312
rect 5961 2244 6063 2278
rect 6097 2244 6135 2278
rect 6169 2244 6271 2278
rect 5961 2210 6271 2244
rect 5961 2176 6063 2210
rect 6097 2176 6135 2210
rect 6169 2176 6271 2210
rect 5961 2142 6271 2176
rect 5961 2108 6063 2142
rect 6097 2108 6135 2142
rect 6169 2108 6271 2142
rect 5961 2074 6271 2108
rect 5961 2040 6063 2074
rect 6097 2040 6135 2074
rect 6169 2040 6271 2074
rect 5961 2006 6271 2040
rect 5961 1972 6063 2006
rect 6097 1972 6135 2006
rect 6169 1972 6271 2006
rect 5961 1938 6271 1972
rect 5961 1904 6063 1938
rect 6097 1904 6135 1938
rect 6169 1904 6271 1938
rect 5961 1870 6271 1904
rect 5961 1836 6063 1870
rect 6097 1836 6135 1870
rect 6169 1836 6271 1870
rect 5961 1802 6271 1836
rect 5961 1768 6063 1802
rect 6097 1768 6135 1802
rect 6169 1768 6271 1802
rect 5961 1734 6271 1768
rect 5961 1700 6063 1734
rect 6097 1700 6135 1734
rect 6169 1700 6271 1734
rect 5961 1666 6271 1700
rect 5961 1632 6063 1666
rect 6097 1632 6135 1666
rect 6169 1632 6271 1666
rect 5961 1598 6271 1632
rect 5961 1564 6063 1598
rect 6097 1564 6135 1598
rect 6169 1564 6271 1598
rect 5961 1552 6271 1564
rect 6391 2540 6542 2552
rect 6682 2540 6833 2552
rect 6391 2506 6493 2540
rect 6527 2506 6542 2540
rect 6682 2506 6697 2540
rect 6731 2506 6833 2540
rect 6391 2472 6542 2506
rect 6682 2472 6833 2506
rect 6391 2438 6493 2472
rect 6527 2438 6542 2472
rect 6682 2438 6697 2472
rect 6731 2438 6833 2472
rect 6391 2404 6542 2438
rect 6682 2404 6833 2438
rect 6391 2370 6493 2404
rect 6527 2370 6542 2404
rect 6682 2370 6697 2404
rect 6731 2370 6833 2404
rect 6391 2336 6542 2370
rect 6682 2336 6833 2370
rect 6391 2302 6493 2336
rect 6527 2302 6542 2336
rect 6682 2302 6697 2336
rect 6731 2302 6833 2336
rect 6391 2268 6542 2302
rect 6682 2268 6833 2302
rect 6391 2234 6493 2268
rect 6527 2234 6542 2268
rect 6682 2234 6697 2268
rect 6731 2234 6833 2268
rect 6391 2200 6542 2234
rect 6682 2200 6833 2234
rect 6391 2166 6493 2200
rect 6527 2166 6542 2200
rect 6682 2166 6697 2200
rect 6731 2166 6833 2200
rect 6391 2132 6542 2166
rect 6682 2132 6833 2166
rect 6391 2098 6493 2132
rect 6527 2098 6542 2132
rect 6682 2098 6697 2132
rect 6731 2098 6833 2132
rect 6391 2064 6542 2098
rect 6682 2064 6833 2098
rect 6391 2030 6493 2064
rect 6527 2030 6542 2064
rect 6682 2030 6697 2064
rect 6731 2030 6833 2064
rect 6391 1996 6542 2030
rect 6682 1996 6833 2030
rect 6391 1962 6493 1996
rect 6527 1962 6542 1996
rect 6682 1962 6697 1996
rect 6731 1962 6833 1996
rect 6391 1928 6542 1962
rect 6682 1928 6833 1962
rect 6391 1894 6493 1928
rect 6527 1894 6542 1928
rect 6682 1894 6697 1928
rect 6731 1894 6833 1928
rect 6391 1860 6542 1894
rect 6682 1860 6833 1894
rect 6391 1826 6493 1860
rect 6527 1826 6542 1860
rect 6682 1826 6697 1860
rect 6731 1826 6833 1860
rect 6391 1792 6542 1826
rect 6682 1792 6833 1826
rect 6391 1758 6493 1792
rect 6527 1758 6542 1792
rect 6682 1758 6697 1792
rect 6731 1758 6833 1792
rect 6391 1724 6542 1758
rect 6682 1724 6833 1758
rect 6391 1690 6493 1724
rect 6527 1690 6542 1724
rect 6682 1690 6697 1724
rect 6731 1690 6833 1724
rect 6391 1656 6542 1690
rect 6682 1656 6833 1690
rect 6391 1622 6493 1656
rect 6527 1622 6542 1656
rect 6682 1622 6697 1656
rect 6731 1622 6833 1656
rect 6391 1552 6542 1622
rect 6682 1552 6833 1622
rect 6953 2482 7263 2552
rect 6953 2448 7055 2482
rect 7089 2448 7127 2482
rect 7161 2448 7263 2482
rect 6953 2414 7263 2448
rect 6953 2380 7055 2414
rect 7089 2380 7127 2414
rect 7161 2380 7263 2414
rect 6953 2346 7263 2380
rect 6953 2312 7055 2346
rect 7089 2312 7127 2346
rect 7161 2312 7263 2346
rect 6953 2278 7263 2312
rect 6953 2244 7055 2278
rect 7089 2244 7127 2278
rect 7161 2244 7263 2278
rect 6953 2210 7263 2244
rect 6953 2176 7055 2210
rect 7089 2176 7127 2210
rect 7161 2176 7263 2210
rect 6953 2142 7263 2176
rect 6953 2108 7055 2142
rect 7089 2108 7127 2142
rect 7161 2108 7263 2142
rect 6953 2074 7263 2108
rect 6953 2040 7055 2074
rect 7089 2040 7127 2074
rect 7161 2040 7263 2074
rect 6953 2006 7263 2040
rect 6953 1972 7055 2006
rect 7089 1972 7127 2006
rect 7161 1972 7263 2006
rect 6953 1938 7263 1972
rect 6953 1904 7055 1938
rect 7089 1904 7127 1938
rect 7161 1904 7263 1938
rect 6953 1870 7263 1904
rect 6953 1836 7055 1870
rect 7089 1836 7127 1870
rect 7161 1836 7263 1870
rect 6953 1802 7263 1836
rect 6953 1768 7055 1802
rect 7089 1768 7127 1802
rect 7161 1768 7263 1802
rect 6953 1734 7263 1768
rect 6953 1700 7055 1734
rect 7089 1700 7127 1734
rect 7161 1700 7263 1734
rect 6953 1666 7263 1700
rect 6953 1632 7055 1666
rect 7089 1632 7127 1666
rect 7161 1632 7263 1666
rect 6953 1598 7263 1632
rect 6953 1564 7055 1598
rect 7089 1564 7127 1598
rect 7161 1564 7263 1598
rect 6953 1552 7263 1564
rect 7383 2540 7534 2552
rect 7674 2540 7825 2552
rect 7383 2506 7485 2540
rect 7519 2506 7534 2540
rect 7674 2506 7689 2540
rect 7723 2506 7825 2540
rect 7383 2472 7534 2506
rect 7674 2472 7825 2506
rect 7383 2438 7485 2472
rect 7519 2438 7534 2472
rect 7674 2438 7689 2472
rect 7723 2438 7825 2472
rect 7383 2404 7534 2438
rect 7674 2404 7825 2438
rect 7383 2370 7485 2404
rect 7519 2370 7534 2404
rect 7674 2370 7689 2404
rect 7723 2370 7825 2404
rect 7383 2336 7534 2370
rect 7674 2336 7825 2370
rect 7383 2302 7485 2336
rect 7519 2302 7534 2336
rect 7674 2302 7689 2336
rect 7723 2302 7825 2336
rect 7383 2268 7534 2302
rect 7674 2268 7825 2302
rect 7383 2234 7485 2268
rect 7519 2234 7534 2268
rect 7674 2234 7689 2268
rect 7723 2234 7825 2268
rect 7383 2200 7534 2234
rect 7674 2200 7825 2234
rect 7383 2166 7485 2200
rect 7519 2166 7534 2200
rect 7674 2166 7689 2200
rect 7723 2166 7825 2200
rect 7383 2132 7534 2166
rect 7674 2132 7825 2166
rect 7383 2098 7485 2132
rect 7519 2098 7534 2132
rect 7674 2098 7689 2132
rect 7723 2098 7825 2132
rect 7383 2064 7534 2098
rect 7674 2064 7825 2098
rect 7383 2030 7485 2064
rect 7519 2030 7534 2064
rect 7674 2030 7689 2064
rect 7723 2030 7825 2064
rect 7383 1996 7534 2030
rect 7674 1996 7825 2030
rect 7383 1962 7485 1996
rect 7519 1962 7534 1996
rect 7674 1962 7689 1996
rect 7723 1962 7825 1996
rect 7383 1928 7534 1962
rect 7674 1928 7825 1962
rect 7383 1894 7485 1928
rect 7519 1894 7534 1928
rect 7674 1894 7689 1928
rect 7723 1894 7825 1928
rect 7383 1860 7534 1894
rect 7674 1860 7825 1894
rect 7383 1826 7485 1860
rect 7519 1826 7534 1860
rect 7674 1826 7689 1860
rect 7723 1826 7825 1860
rect 7383 1792 7534 1826
rect 7674 1792 7825 1826
rect 7383 1758 7485 1792
rect 7519 1758 7534 1792
rect 7674 1758 7689 1792
rect 7723 1758 7825 1792
rect 7383 1724 7534 1758
rect 7674 1724 7825 1758
rect 7383 1690 7485 1724
rect 7519 1690 7534 1724
rect 7674 1690 7689 1724
rect 7723 1690 7825 1724
rect 7383 1656 7534 1690
rect 7674 1656 7825 1690
rect 7383 1622 7485 1656
rect 7519 1622 7534 1656
rect 7674 1622 7689 1656
rect 7723 1622 7825 1656
rect 7383 1552 7534 1622
rect 7674 1552 7825 1622
rect 7945 2482 8255 2552
rect 7945 2448 8047 2482
rect 8081 2448 8119 2482
rect 8153 2448 8255 2482
rect 7945 2414 8255 2448
rect 7945 2380 8047 2414
rect 8081 2380 8119 2414
rect 8153 2380 8255 2414
rect 7945 2346 8255 2380
rect 7945 2312 8047 2346
rect 8081 2312 8119 2346
rect 8153 2312 8255 2346
rect 7945 2278 8255 2312
rect 7945 2244 8047 2278
rect 8081 2244 8119 2278
rect 8153 2244 8255 2278
rect 7945 2210 8255 2244
rect 7945 2176 8047 2210
rect 8081 2176 8119 2210
rect 8153 2176 8255 2210
rect 7945 2142 8255 2176
rect 7945 2108 8047 2142
rect 8081 2108 8119 2142
rect 8153 2108 8255 2142
rect 7945 2074 8255 2108
rect 7945 2040 8047 2074
rect 8081 2040 8119 2074
rect 8153 2040 8255 2074
rect 7945 2006 8255 2040
rect 7945 1972 8047 2006
rect 8081 1972 8119 2006
rect 8153 1972 8255 2006
rect 7945 1938 8255 1972
rect 7945 1904 8047 1938
rect 8081 1904 8119 1938
rect 8153 1904 8255 1938
rect 7945 1870 8255 1904
rect 7945 1836 8047 1870
rect 8081 1836 8119 1870
rect 8153 1836 8255 1870
rect 7945 1802 8255 1836
rect 7945 1768 8047 1802
rect 8081 1768 8119 1802
rect 8153 1768 8255 1802
rect 7945 1734 8255 1768
rect 7945 1700 8047 1734
rect 8081 1700 8119 1734
rect 8153 1700 8255 1734
rect 7945 1666 8255 1700
rect 7945 1632 8047 1666
rect 8081 1632 8119 1666
rect 8153 1632 8255 1666
rect 7945 1598 8255 1632
rect 7945 1564 8047 1598
rect 8081 1564 8119 1598
rect 8153 1564 8255 1598
rect 7945 1552 8255 1564
rect 8375 2540 8526 2552
rect 8666 2540 8817 2552
rect 8375 2506 8477 2540
rect 8511 2506 8526 2540
rect 8666 2506 8681 2540
rect 8715 2506 8817 2540
rect 8375 2472 8526 2506
rect 8666 2472 8817 2506
rect 8375 2438 8477 2472
rect 8511 2438 8526 2472
rect 8666 2438 8681 2472
rect 8715 2438 8817 2472
rect 8375 2404 8526 2438
rect 8666 2404 8817 2438
rect 8375 2370 8477 2404
rect 8511 2370 8526 2404
rect 8666 2370 8681 2404
rect 8715 2370 8817 2404
rect 8375 2336 8526 2370
rect 8666 2336 8817 2370
rect 8375 2302 8477 2336
rect 8511 2302 8526 2336
rect 8666 2302 8681 2336
rect 8715 2302 8817 2336
rect 8375 2268 8526 2302
rect 8666 2268 8817 2302
rect 8375 2234 8477 2268
rect 8511 2234 8526 2268
rect 8666 2234 8681 2268
rect 8715 2234 8817 2268
rect 8375 2200 8526 2234
rect 8666 2200 8817 2234
rect 8375 2166 8477 2200
rect 8511 2166 8526 2200
rect 8666 2166 8681 2200
rect 8715 2166 8817 2200
rect 8375 2132 8526 2166
rect 8666 2132 8817 2166
rect 8375 2098 8477 2132
rect 8511 2098 8526 2132
rect 8666 2098 8681 2132
rect 8715 2098 8817 2132
rect 8375 2064 8526 2098
rect 8666 2064 8817 2098
rect 8375 2030 8477 2064
rect 8511 2030 8526 2064
rect 8666 2030 8681 2064
rect 8715 2030 8817 2064
rect 8375 1996 8526 2030
rect 8666 1996 8817 2030
rect 8375 1962 8477 1996
rect 8511 1962 8526 1996
rect 8666 1962 8681 1996
rect 8715 1962 8817 1996
rect 8375 1928 8526 1962
rect 8666 1928 8817 1962
rect 8375 1894 8477 1928
rect 8511 1894 8526 1928
rect 8666 1894 8681 1928
rect 8715 1894 8817 1928
rect 8375 1860 8526 1894
rect 8666 1860 8817 1894
rect 8375 1826 8477 1860
rect 8511 1826 8526 1860
rect 8666 1826 8681 1860
rect 8715 1826 8817 1860
rect 8375 1792 8526 1826
rect 8666 1792 8817 1826
rect 8375 1758 8477 1792
rect 8511 1758 8526 1792
rect 8666 1758 8681 1792
rect 8715 1758 8817 1792
rect 8375 1724 8526 1758
rect 8666 1724 8817 1758
rect 8375 1690 8477 1724
rect 8511 1690 8526 1724
rect 8666 1690 8681 1724
rect 8715 1690 8817 1724
rect 8375 1656 8526 1690
rect 8666 1656 8817 1690
rect 8375 1622 8477 1656
rect 8511 1622 8526 1656
rect 8666 1622 8681 1656
rect 8715 1622 8817 1656
rect 8375 1552 8526 1622
rect 8666 1552 8817 1622
rect 8937 2482 9247 2552
rect 8937 2448 9039 2482
rect 9073 2448 9111 2482
rect 9145 2448 9247 2482
rect 8937 2414 9247 2448
rect 8937 2380 9039 2414
rect 9073 2380 9111 2414
rect 9145 2380 9247 2414
rect 8937 2346 9247 2380
rect 8937 2312 9039 2346
rect 9073 2312 9111 2346
rect 9145 2312 9247 2346
rect 8937 2278 9247 2312
rect 8937 2244 9039 2278
rect 9073 2244 9111 2278
rect 9145 2244 9247 2278
rect 8937 2210 9247 2244
rect 8937 2176 9039 2210
rect 9073 2176 9111 2210
rect 9145 2176 9247 2210
rect 8937 2142 9247 2176
rect 8937 2108 9039 2142
rect 9073 2108 9111 2142
rect 9145 2108 9247 2142
rect 8937 2074 9247 2108
rect 8937 2040 9039 2074
rect 9073 2040 9111 2074
rect 9145 2040 9247 2074
rect 8937 2006 9247 2040
rect 8937 1972 9039 2006
rect 9073 1972 9111 2006
rect 9145 1972 9247 2006
rect 8937 1938 9247 1972
rect 8937 1904 9039 1938
rect 9073 1904 9111 1938
rect 9145 1904 9247 1938
rect 8937 1870 9247 1904
rect 8937 1836 9039 1870
rect 9073 1836 9111 1870
rect 9145 1836 9247 1870
rect 8937 1802 9247 1836
rect 8937 1768 9039 1802
rect 9073 1768 9111 1802
rect 9145 1768 9247 1802
rect 8937 1734 9247 1768
rect 8937 1700 9039 1734
rect 9073 1700 9111 1734
rect 9145 1700 9247 1734
rect 8937 1666 9247 1700
rect 8937 1632 9039 1666
rect 9073 1632 9111 1666
rect 9145 1632 9247 1666
rect 8937 1598 9247 1632
rect 8937 1564 9039 1598
rect 9073 1564 9111 1598
rect 9145 1564 9247 1598
rect 8937 1552 9247 1564
rect 9367 2540 9518 2552
rect 9658 2540 9809 2552
rect 9367 2506 9469 2540
rect 9503 2506 9518 2540
rect 9658 2506 9673 2540
rect 9707 2506 9809 2540
rect 9367 2472 9518 2506
rect 9658 2472 9809 2506
rect 9367 2438 9469 2472
rect 9503 2438 9518 2472
rect 9658 2438 9673 2472
rect 9707 2438 9809 2472
rect 9367 2404 9518 2438
rect 9658 2404 9809 2438
rect 9367 2370 9469 2404
rect 9503 2370 9518 2404
rect 9658 2370 9673 2404
rect 9707 2370 9809 2404
rect 9367 2336 9518 2370
rect 9658 2336 9809 2370
rect 9367 2302 9469 2336
rect 9503 2302 9518 2336
rect 9658 2302 9673 2336
rect 9707 2302 9809 2336
rect 9367 2268 9518 2302
rect 9658 2268 9809 2302
rect 9367 2234 9469 2268
rect 9503 2234 9518 2268
rect 9658 2234 9673 2268
rect 9707 2234 9809 2268
rect 9367 2200 9518 2234
rect 9658 2200 9809 2234
rect 9367 2166 9469 2200
rect 9503 2166 9518 2200
rect 9658 2166 9673 2200
rect 9707 2166 9809 2200
rect 9367 2132 9518 2166
rect 9658 2132 9809 2166
rect 9367 2098 9469 2132
rect 9503 2098 9518 2132
rect 9658 2098 9673 2132
rect 9707 2098 9809 2132
rect 9367 2064 9518 2098
rect 9658 2064 9809 2098
rect 9367 2030 9469 2064
rect 9503 2030 9518 2064
rect 9658 2030 9673 2064
rect 9707 2030 9809 2064
rect 9367 1996 9518 2030
rect 9658 1996 9809 2030
rect 9367 1962 9469 1996
rect 9503 1962 9518 1996
rect 9658 1962 9673 1996
rect 9707 1962 9809 1996
rect 9367 1928 9518 1962
rect 9658 1928 9809 1962
rect 9367 1894 9469 1928
rect 9503 1894 9518 1928
rect 9658 1894 9673 1928
rect 9707 1894 9809 1928
rect 9367 1860 9518 1894
rect 9658 1860 9809 1894
rect 9367 1826 9469 1860
rect 9503 1826 9518 1860
rect 9658 1826 9673 1860
rect 9707 1826 9809 1860
rect 9367 1792 9518 1826
rect 9658 1792 9809 1826
rect 9367 1758 9469 1792
rect 9503 1758 9518 1792
rect 9658 1758 9673 1792
rect 9707 1758 9809 1792
rect 9367 1724 9518 1758
rect 9658 1724 9809 1758
rect 9367 1690 9469 1724
rect 9503 1690 9518 1724
rect 9658 1690 9673 1724
rect 9707 1690 9809 1724
rect 9367 1656 9518 1690
rect 9658 1656 9809 1690
rect 9367 1622 9469 1656
rect 9503 1622 9518 1656
rect 9658 1622 9673 1656
rect 9707 1622 9809 1656
rect 9367 1552 9518 1622
rect 9658 1552 9809 1622
rect 9929 2482 10239 2552
rect 9929 2448 10031 2482
rect 10065 2448 10103 2482
rect 10137 2448 10239 2482
rect 9929 2414 10239 2448
rect 9929 2380 10031 2414
rect 10065 2380 10103 2414
rect 10137 2380 10239 2414
rect 9929 2346 10239 2380
rect 9929 2312 10031 2346
rect 10065 2312 10103 2346
rect 10137 2312 10239 2346
rect 9929 2278 10239 2312
rect 9929 2244 10031 2278
rect 10065 2244 10103 2278
rect 10137 2244 10239 2278
rect 9929 2210 10239 2244
rect 9929 2176 10031 2210
rect 10065 2176 10103 2210
rect 10137 2176 10239 2210
rect 9929 2142 10239 2176
rect 9929 2108 10031 2142
rect 10065 2108 10103 2142
rect 10137 2108 10239 2142
rect 9929 2074 10239 2108
rect 9929 2040 10031 2074
rect 10065 2040 10103 2074
rect 10137 2040 10239 2074
rect 9929 2006 10239 2040
rect 9929 1972 10031 2006
rect 10065 1972 10103 2006
rect 10137 1972 10239 2006
rect 9929 1938 10239 1972
rect 9929 1904 10031 1938
rect 10065 1904 10103 1938
rect 10137 1904 10239 1938
rect 9929 1870 10239 1904
rect 9929 1836 10031 1870
rect 10065 1836 10103 1870
rect 10137 1836 10239 1870
rect 9929 1802 10239 1836
rect 9929 1768 10031 1802
rect 10065 1768 10103 1802
rect 10137 1768 10239 1802
rect 9929 1734 10239 1768
rect 9929 1700 10031 1734
rect 10065 1700 10103 1734
rect 10137 1700 10239 1734
rect 9929 1666 10239 1700
rect 9929 1632 10031 1666
rect 10065 1632 10103 1666
rect 10137 1632 10239 1666
rect 9929 1598 10239 1632
rect 9929 1564 10031 1598
rect 10065 1564 10103 1598
rect 10137 1564 10239 1598
rect 9929 1552 10239 1564
rect 10359 2540 10510 2552
rect 10650 2540 10801 2552
rect 10359 2506 10461 2540
rect 10495 2506 10510 2540
rect 10650 2506 10665 2540
rect 10699 2506 10801 2540
rect 10359 2472 10510 2506
rect 10650 2472 10801 2506
rect 10359 2438 10461 2472
rect 10495 2438 10510 2472
rect 10650 2438 10665 2472
rect 10699 2438 10801 2472
rect 10359 2404 10510 2438
rect 10650 2404 10801 2438
rect 10359 2370 10461 2404
rect 10495 2370 10510 2404
rect 10650 2370 10665 2404
rect 10699 2370 10801 2404
rect 10359 2336 10510 2370
rect 10650 2336 10801 2370
rect 10359 2302 10461 2336
rect 10495 2302 10510 2336
rect 10650 2302 10665 2336
rect 10699 2302 10801 2336
rect 10359 2268 10510 2302
rect 10650 2268 10801 2302
rect 10359 2234 10461 2268
rect 10495 2234 10510 2268
rect 10650 2234 10665 2268
rect 10699 2234 10801 2268
rect 10359 2200 10510 2234
rect 10650 2200 10801 2234
rect 10359 2166 10461 2200
rect 10495 2166 10510 2200
rect 10650 2166 10665 2200
rect 10699 2166 10801 2200
rect 10359 2132 10510 2166
rect 10650 2132 10801 2166
rect 10359 2098 10461 2132
rect 10495 2098 10510 2132
rect 10650 2098 10665 2132
rect 10699 2098 10801 2132
rect 10359 2064 10510 2098
rect 10650 2064 10801 2098
rect 10359 2030 10461 2064
rect 10495 2030 10510 2064
rect 10650 2030 10665 2064
rect 10699 2030 10801 2064
rect 10359 1996 10510 2030
rect 10650 1996 10801 2030
rect 10359 1962 10461 1996
rect 10495 1962 10510 1996
rect 10650 1962 10665 1996
rect 10699 1962 10801 1996
rect 10359 1928 10510 1962
rect 10650 1928 10801 1962
rect 10359 1894 10461 1928
rect 10495 1894 10510 1928
rect 10650 1894 10665 1928
rect 10699 1894 10801 1928
rect 10359 1860 10510 1894
rect 10650 1860 10801 1894
rect 10359 1826 10461 1860
rect 10495 1826 10510 1860
rect 10650 1826 10665 1860
rect 10699 1826 10801 1860
rect 10359 1792 10510 1826
rect 10650 1792 10801 1826
rect 10359 1758 10461 1792
rect 10495 1758 10510 1792
rect 10650 1758 10665 1792
rect 10699 1758 10801 1792
rect 10359 1724 10510 1758
rect 10650 1724 10801 1758
rect 10359 1690 10461 1724
rect 10495 1690 10510 1724
rect 10650 1690 10665 1724
rect 10699 1690 10801 1724
rect 10359 1656 10510 1690
rect 10650 1656 10801 1690
rect 10359 1622 10461 1656
rect 10495 1622 10510 1656
rect 10650 1622 10665 1656
rect 10699 1622 10801 1656
rect 10359 1552 10510 1622
rect 10650 1552 10801 1622
rect 10921 2482 11231 2552
rect 10921 2448 11023 2482
rect 11057 2448 11095 2482
rect 11129 2448 11231 2482
rect 10921 2414 11231 2448
rect 10921 2380 11023 2414
rect 11057 2380 11095 2414
rect 11129 2380 11231 2414
rect 10921 2346 11231 2380
rect 10921 2312 11023 2346
rect 11057 2312 11095 2346
rect 11129 2312 11231 2346
rect 10921 2278 11231 2312
rect 10921 2244 11023 2278
rect 11057 2244 11095 2278
rect 11129 2244 11231 2278
rect 10921 2210 11231 2244
rect 10921 2176 11023 2210
rect 11057 2176 11095 2210
rect 11129 2176 11231 2210
rect 10921 2142 11231 2176
rect 10921 2108 11023 2142
rect 11057 2108 11095 2142
rect 11129 2108 11231 2142
rect 10921 2074 11231 2108
rect 10921 2040 11023 2074
rect 11057 2040 11095 2074
rect 11129 2040 11231 2074
rect 10921 2006 11231 2040
rect 10921 1972 11023 2006
rect 11057 1972 11095 2006
rect 11129 1972 11231 2006
rect 10921 1938 11231 1972
rect 10921 1904 11023 1938
rect 11057 1904 11095 1938
rect 11129 1904 11231 1938
rect 10921 1870 11231 1904
rect 10921 1836 11023 1870
rect 11057 1836 11095 1870
rect 11129 1836 11231 1870
rect 10921 1802 11231 1836
rect 10921 1768 11023 1802
rect 11057 1768 11095 1802
rect 11129 1768 11231 1802
rect 10921 1734 11231 1768
rect 10921 1700 11023 1734
rect 11057 1700 11095 1734
rect 11129 1700 11231 1734
rect 10921 1666 11231 1700
rect 10921 1632 11023 1666
rect 11057 1632 11095 1666
rect 11129 1632 11231 1666
rect 10921 1598 11231 1632
rect 10921 1564 11023 1598
rect 11057 1564 11095 1598
rect 11129 1564 11231 1598
rect 10921 1552 11231 1564
rect 11351 2540 11502 2552
rect 11642 2540 11793 2552
rect 11351 2506 11453 2540
rect 11487 2506 11502 2540
rect 11642 2506 11657 2540
rect 11691 2506 11793 2540
rect 11351 2472 11502 2506
rect 11642 2472 11793 2506
rect 11351 2438 11453 2472
rect 11487 2438 11502 2472
rect 11642 2438 11657 2472
rect 11691 2438 11793 2472
rect 11351 2404 11502 2438
rect 11642 2404 11793 2438
rect 11351 2370 11453 2404
rect 11487 2370 11502 2404
rect 11642 2370 11657 2404
rect 11691 2370 11793 2404
rect 11351 2336 11502 2370
rect 11642 2336 11793 2370
rect 11351 2302 11453 2336
rect 11487 2302 11502 2336
rect 11642 2302 11657 2336
rect 11691 2302 11793 2336
rect 11351 2268 11502 2302
rect 11642 2268 11793 2302
rect 11351 2234 11453 2268
rect 11487 2234 11502 2268
rect 11642 2234 11657 2268
rect 11691 2234 11793 2268
rect 11351 2200 11502 2234
rect 11642 2200 11793 2234
rect 11351 2166 11453 2200
rect 11487 2166 11502 2200
rect 11642 2166 11657 2200
rect 11691 2166 11793 2200
rect 11351 2132 11502 2166
rect 11642 2132 11793 2166
rect 11351 2098 11453 2132
rect 11487 2098 11502 2132
rect 11642 2098 11657 2132
rect 11691 2098 11793 2132
rect 11351 2064 11502 2098
rect 11642 2064 11793 2098
rect 11351 2030 11453 2064
rect 11487 2030 11502 2064
rect 11642 2030 11657 2064
rect 11691 2030 11793 2064
rect 11351 1996 11502 2030
rect 11642 1996 11793 2030
rect 11351 1962 11453 1996
rect 11487 1962 11502 1996
rect 11642 1962 11657 1996
rect 11691 1962 11793 1996
rect 11351 1928 11502 1962
rect 11642 1928 11793 1962
rect 11351 1894 11453 1928
rect 11487 1894 11502 1928
rect 11642 1894 11657 1928
rect 11691 1894 11793 1928
rect 11351 1860 11502 1894
rect 11642 1860 11793 1894
rect 11351 1826 11453 1860
rect 11487 1826 11502 1860
rect 11642 1826 11657 1860
rect 11691 1826 11793 1860
rect 11351 1792 11502 1826
rect 11642 1792 11793 1826
rect 11351 1758 11453 1792
rect 11487 1758 11502 1792
rect 11642 1758 11657 1792
rect 11691 1758 11793 1792
rect 11351 1724 11502 1758
rect 11642 1724 11793 1758
rect 11351 1690 11453 1724
rect 11487 1690 11502 1724
rect 11642 1690 11657 1724
rect 11691 1690 11793 1724
rect 11351 1656 11502 1690
rect 11642 1656 11793 1690
rect 11351 1622 11453 1656
rect 11487 1622 11502 1656
rect 11642 1622 11657 1656
rect 11691 1622 11793 1656
rect 11351 1552 11502 1622
rect 11642 1552 11793 1622
rect 11913 2482 12223 2552
rect 11913 2448 12015 2482
rect 12049 2448 12087 2482
rect 12121 2448 12223 2482
rect 11913 2414 12223 2448
rect 11913 2380 12015 2414
rect 12049 2380 12087 2414
rect 12121 2380 12223 2414
rect 11913 2346 12223 2380
rect 11913 2312 12015 2346
rect 12049 2312 12087 2346
rect 12121 2312 12223 2346
rect 11913 2278 12223 2312
rect 11913 2244 12015 2278
rect 12049 2244 12087 2278
rect 12121 2244 12223 2278
rect 11913 2210 12223 2244
rect 11913 2176 12015 2210
rect 12049 2176 12087 2210
rect 12121 2176 12223 2210
rect 11913 2142 12223 2176
rect 11913 2108 12015 2142
rect 12049 2108 12087 2142
rect 12121 2108 12223 2142
rect 11913 2074 12223 2108
rect 11913 2040 12015 2074
rect 12049 2040 12087 2074
rect 12121 2040 12223 2074
rect 11913 2006 12223 2040
rect 11913 1972 12015 2006
rect 12049 1972 12087 2006
rect 12121 1972 12223 2006
rect 11913 1938 12223 1972
rect 11913 1904 12015 1938
rect 12049 1904 12087 1938
rect 12121 1904 12223 1938
rect 11913 1870 12223 1904
rect 11913 1836 12015 1870
rect 12049 1836 12087 1870
rect 12121 1836 12223 1870
rect 11913 1802 12223 1836
rect 11913 1768 12015 1802
rect 12049 1768 12087 1802
rect 12121 1768 12223 1802
rect 11913 1734 12223 1768
rect 11913 1700 12015 1734
rect 12049 1700 12087 1734
rect 12121 1700 12223 1734
rect 11913 1666 12223 1700
rect 11913 1632 12015 1666
rect 12049 1632 12087 1666
rect 12121 1632 12223 1666
rect 11913 1598 12223 1632
rect 11913 1564 12015 1598
rect 12049 1564 12087 1598
rect 12121 1564 12223 1598
rect 11913 1552 12223 1564
rect 12343 2540 12494 2552
rect 12634 2540 12785 2552
rect 12343 2506 12445 2540
rect 12479 2506 12494 2540
rect 12634 2506 12649 2540
rect 12683 2506 12785 2540
rect 12343 2472 12494 2506
rect 12634 2472 12785 2506
rect 12343 2438 12445 2472
rect 12479 2438 12494 2472
rect 12634 2438 12649 2472
rect 12683 2438 12785 2472
rect 12343 2404 12494 2438
rect 12634 2404 12785 2438
rect 12343 2370 12445 2404
rect 12479 2370 12494 2404
rect 12634 2370 12649 2404
rect 12683 2370 12785 2404
rect 12343 2336 12494 2370
rect 12634 2336 12785 2370
rect 12343 2302 12445 2336
rect 12479 2302 12494 2336
rect 12634 2302 12649 2336
rect 12683 2302 12785 2336
rect 12343 2268 12494 2302
rect 12634 2268 12785 2302
rect 12343 2234 12445 2268
rect 12479 2234 12494 2268
rect 12634 2234 12649 2268
rect 12683 2234 12785 2268
rect 12343 2200 12494 2234
rect 12634 2200 12785 2234
rect 12343 2166 12445 2200
rect 12479 2166 12494 2200
rect 12634 2166 12649 2200
rect 12683 2166 12785 2200
rect 12343 2132 12494 2166
rect 12634 2132 12785 2166
rect 12343 2098 12445 2132
rect 12479 2098 12494 2132
rect 12634 2098 12649 2132
rect 12683 2098 12785 2132
rect 12343 2064 12494 2098
rect 12634 2064 12785 2098
rect 12343 2030 12445 2064
rect 12479 2030 12494 2064
rect 12634 2030 12649 2064
rect 12683 2030 12785 2064
rect 12343 1996 12494 2030
rect 12634 1996 12785 2030
rect 12343 1962 12445 1996
rect 12479 1962 12494 1996
rect 12634 1962 12649 1996
rect 12683 1962 12785 1996
rect 12343 1928 12494 1962
rect 12634 1928 12785 1962
rect 12343 1894 12445 1928
rect 12479 1894 12494 1928
rect 12634 1894 12649 1928
rect 12683 1894 12785 1928
rect 12343 1860 12494 1894
rect 12634 1860 12785 1894
rect 12343 1826 12445 1860
rect 12479 1826 12494 1860
rect 12634 1826 12649 1860
rect 12683 1826 12785 1860
rect 12343 1792 12494 1826
rect 12634 1792 12785 1826
rect 12343 1758 12445 1792
rect 12479 1758 12494 1792
rect 12634 1758 12649 1792
rect 12683 1758 12785 1792
rect 12343 1724 12494 1758
rect 12634 1724 12785 1758
rect 12343 1690 12445 1724
rect 12479 1690 12494 1724
rect 12634 1690 12649 1724
rect 12683 1690 12785 1724
rect 12343 1656 12494 1690
rect 12634 1656 12785 1690
rect 12343 1622 12445 1656
rect 12479 1622 12494 1656
rect 12634 1622 12649 1656
rect 12683 1622 12785 1656
rect 12343 1552 12494 1622
rect 12634 1552 12785 1622
rect 12905 2482 13215 2552
rect 12905 2448 13007 2482
rect 13041 2448 13079 2482
rect 13113 2448 13215 2482
rect 12905 2414 13215 2448
rect 12905 2380 13007 2414
rect 13041 2380 13079 2414
rect 13113 2380 13215 2414
rect 12905 2346 13215 2380
rect 12905 2312 13007 2346
rect 13041 2312 13079 2346
rect 13113 2312 13215 2346
rect 12905 2278 13215 2312
rect 12905 2244 13007 2278
rect 13041 2244 13079 2278
rect 13113 2244 13215 2278
rect 12905 2210 13215 2244
rect 12905 2176 13007 2210
rect 13041 2176 13079 2210
rect 13113 2176 13215 2210
rect 12905 2142 13215 2176
rect 12905 2108 13007 2142
rect 13041 2108 13079 2142
rect 13113 2108 13215 2142
rect 12905 2074 13215 2108
rect 12905 2040 13007 2074
rect 13041 2040 13079 2074
rect 13113 2040 13215 2074
rect 12905 2006 13215 2040
rect 12905 1972 13007 2006
rect 13041 1972 13079 2006
rect 13113 1972 13215 2006
rect 12905 1938 13215 1972
rect 12905 1904 13007 1938
rect 13041 1904 13079 1938
rect 13113 1904 13215 1938
rect 12905 1870 13215 1904
rect 12905 1836 13007 1870
rect 13041 1836 13079 1870
rect 13113 1836 13215 1870
rect 12905 1802 13215 1836
rect 12905 1768 13007 1802
rect 13041 1768 13079 1802
rect 13113 1768 13215 1802
rect 12905 1734 13215 1768
rect 12905 1700 13007 1734
rect 13041 1700 13079 1734
rect 13113 1700 13215 1734
rect 12905 1666 13215 1700
rect 12905 1632 13007 1666
rect 13041 1632 13079 1666
rect 13113 1632 13215 1666
rect 12905 1598 13215 1632
rect 12905 1564 13007 1598
rect 13041 1564 13079 1598
rect 13113 1564 13215 1598
rect 12905 1552 13215 1564
rect 13335 2540 13486 2552
rect 13626 2540 13777 2552
rect 13335 2506 13437 2540
rect 13471 2506 13486 2540
rect 13626 2506 13641 2540
rect 13675 2506 13777 2540
rect 13335 2472 13486 2506
rect 13626 2472 13777 2506
rect 13335 2438 13437 2472
rect 13471 2438 13486 2472
rect 13626 2438 13641 2472
rect 13675 2438 13777 2472
rect 13335 2404 13486 2438
rect 13626 2404 13777 2438
rect 13335 2370 13437 2404
rect 13471 2370 13486 2404
rect 13626 2370 13641 2404
rect 13675 2370 13777 2404
rect 13335 2336 13486 2370
rect 13626 2336 13777 2370
rect 13335 2302 13437 2336
rect 13471 2302 13486 2336
rect 13626 2302 13641 2336
rect 13675 2302 13777 2336
rect 13335 2268 13486 2302
rect 13626 2268 13777 2302
rect 13335 2234 13437 2268
rect 13471 2234 13486 2268
rect 13626 2234 13641 2268
rect 13675 2234 13777 2268
rect 13335 2200 13486 2234
rect 13626 2200 13777 2234
rect 13335 2166 13437 2200
rect 13471 2166 13486 2200
rect 13626 2166 13641 2200
rect 13675 2166 13777 2200
rect 13335 2132 13486 2166
rect 13626 2132 13777 2166
rect 13335 2098 13437 2132
rect 13471 2098 13486 2132
rect 13626 2098 13641 2132
rect 13675 2098 13777 2132
rect 13335 2064 13486 2098
rect 13626 2064 13777 2098
rect 13335 2030 13437 2064
rect 13471 2030 13486 2064
rect 13626 2030 13641 2064
rect 13675 2030 13777 2064
rect 13335 1996 13486 2030
rect 13626 1996 13777 2030
rect 13335 1962 13437 1996
rect 13471 1962 13486 1996
rect 13626 1962 13641 1996
rect 13675 1962 13777 1996
rect 13335 1928 13486 1962
rect 13626 1928 13777 1962
rect 13335 1894 13437 1928
rect 13471 1894 13486 1928
rect 13626 1894 13641 1928
rect 13675 1894 13777 1928
rect 13335 1860 13486 1894
rect 13626 1860 13777 1894
rect 13335 1826 13437 1860
rect 13471 1826 13486 1860
rect 13626 1826 13641 1860
rect 13675 1826 13777 1860
rect 13335 1792 13486 1826
rect 13626 1792 13777 1826
rect 13335 1758 13437 1792
rect 13471 1758 13486 1792
rect 13626 1758 13641 1792
rect 13675 1758 13777 1792
rect 13335 1724 13486 1758
rect 13626 1724 13777 1758
rect 13335 1690 13437 1724
rect 13471 1690 13486 1724
rect 13626 1690 13641 1724
rect 13675 1690 13777 1724
rect 13335 1656 13486 1690
rect 13626 1656 13777 1690
rect 13335 1622 13437 1656
rect 13471 1622 13486 1656
rect 13626 1622 13641 1656
rect 13675 1622 13777 1656
rect 13335 1552 13486 1622
rect 13626 1552 13777 1622
rect 13897 2482 14135 2552
rect 13897 2448 13999 2482
rect 14033 2448 14135 2482
rect 13897 2414 14135 2448
rect 13897 2380 13999 2414
rect 14033 2380 14135 2414
rect 13897 2346 14135 2380
rect 13897 2312 13999 2346
rect 14033 2312 14135 2346
rect 13897 2278 14135 2312
rect 13897 2244 13999 2278
rect 14033 2244 14135 2278
rect 13897 2210 14135 2244
rect 13897 2176 13999 2210
rect 14033 2176 14135 2210
rect 13897 2142 14135 2176
rect 13897 2108 13999 2142
rect 14033 2108 14135 2142
rect 13897 2074 14135 2108
rect 13897 2040 13999 2074
rect 14033 2040 14135 2074
rect 13897 2006 14135 2040
rect 13897 1972 13999 2006
rect 14033 1972 14135 2006
rect 13897 1938 14135 1972
rect 13897 1904 13999 1938
rect 14033 1904 14135 1938
rect 13897 1870 14135 1904
rect 13897 1836 13999 1870
rect 14033 1836 14135 1870
rect 13897 1802 14135 1836
rect 13897 1768 13999 1802
rect 14033 1768 14135 1802
rect 13897 1734 14135 1768
rect 13897 1700 13999 1734
rect 14033 1700 14135 1734
rect 13897 1666 14135 1700
rect 13897 1632 13999 1666
rect 14033 1632 14135 1666
rect 13897 1598 14135 1632
rect 13897 1564 13999 1598
rect 14033 1564 14135 1598
rect 13897 1552 14135 1564
rect 14255 2482 14427 2552
rect 14255 2448 14356 2482
rect 14390 2448 14427 2482
rect 14255 2414 14427 2448
rect 14255 2380 14356 2414
rect 14390 2380 14427 2414
rect 14255 2346 14427 2380
rect 14255 2312 14356 2346
rect 14390 2312 14427 2346
rect 14255 2278 14427 2312
rect 14255 2244 14356 2278
rect 14390 2244 14427 2278
rect 14255 2210 14427 2244
rect 14255 2176 14356 2210
rect 14390 2176 14427 2210
rect 14255 2142 14427 2176
rect 14255 2108 14356 2142
rect 14390 2108 14427 2142
rect 14255 2074 14427 2108
rect 14255 2040 14356 2074
rect 14390 2040 14427 2074
rect 14255 2006 14427 2040
rect 14255 1972 14356 2006
rect 14390 1972 14427 2006
rect 14255 1938 14427 1972
rect 14255 1904 14356 1938
rect 14390 1904 14427 1938
rect 14255 1870 14427 1904
rect 14255 1836 14356 1870
rect 14390 1836 14427 1870
rect 14255 1802 14427 1836
rect 14255 1768 14356 1802
rect 14390 1768 14427 1802
rect 14255 1734 14427 1768
rect 14255 1700 14356 1734
rect 14390 1700 14427 1734
rect 14255 1666 14427 1700
rect 14255 1632 14356 1666
rect 14390 1632 14427 1666
rect 14255 1598 14427 1632
rect 14255 1564 14356 1598
rect 14390 1564 14427 1598
rect 14255 1552 14427 1564
<< mvpdiffc >>
rect 745 4048 779 4082
rect 745 3980 779 4014
rect 745 3912 779 3946
rect 745 3844 779 3878
rect 745 3776 779 3810
rect 745 3708 779 3742
rect 745 3640 779 3674
rect 745 3572 779 3606
rect 745 3504 779 3538
rect 745 3436 779 3470
rect 745 3368 779 3402
rect 745 3300 779 3334
rect 745 3232 779 3266
rect 745 3164 779 3198
rect 1103 4048 1137 4082
rect 1175 4048 1209 4082
rect 1103 3980 1137 4014
rect 1175 3980 1209 4014
rect 1103 3912 1137 3946
rect 1175 3912 1209 3946
rect 1103 3844 1137 3878
rect 1175 3844 1209 3878
rect 1103 3776 1137 3810
rect 1175 3776 1209 3810
rect 1103 3708 1137 3742
rect 1175 3708 1209 3742
rect 1103 3640 1137 3674
rect 1175 3640 1209 3674
rect 1103 3572 1137 3606
rect 1175 3572 1209 3606
rect 1103 3504 1137 3538
rect 1175 3504 1209 3538
rect 1103 3436 1137 3470
rect 1175 3436 1209 3470
rect 1103 3368 1137 3402
rect 1175 3368 1209 3402
rect 1103 3300 1137 3334
rect 1175 3300 1209 3334
rect 1103 3232 1137 3266
rect 1175 3232 1209 3266
rect 1103 3164 1137 3198
rect 1175 3164 1209 3198
rect 1533 4048 1567 4082
rect 1737 4048 1771 4082
rect 1533 3980 1567 4014
rect 1737 3980 1771 4014
rect 1533 3912 1567 3946
rect 1737 3912 1771 3946
rect 1533 3844 1567 3878
rect 1737 3844 1771 3878
rect 1533 3776 1567 3810
rect 1737 3776 1771 3810
rect 1533 3708 1567 3742
rect 1737 3708 1771 3742
rect 1533 3640 1567 3674
rect 1737 3640 1771 3674
rect 1533 3572 1567 3606
rect 1737 3572 1771 3606
rect 1533 3504 1567 3538
rect 1737 3504 1771 3538
rect 1533 3436 1567 3470
rect 1737 3436 1771 3470
rect 1533 3368 1567 3402
rect 1737 3368 1771 3402
rect 1533 3300 1567 3334
rect 1737 3300 1771 3334
rect 1533 3232 1567 3266
rect 1737 3232 1771 3266
rect 1533 3164 1567 3198
rect 1737 3164 1771 3198
rect 2095 4048 2129 4082
rect 2167 4048 2201 4082
rect 2095 3980 2129 4014
rect 2167 3980 2201 4014
rect 2095 3912 2129 3946
rect 2167 3912 2201 3946
rect 2095 3844 2129 3878
rect 2167 3844 2201 3878
rect 2095 3776 2129 3810
rect 2167 3776 2201 3810
rect 2095 3708 2129 3742
rect 2167 3708 2201 3742
rect 2095 3640 2129 3674
rect 2167 3640 2201 3674
rect 2095 3572 2129 3606
rect 2167 3572 2201 3606
rect 2095 3504 2129 3538
rect 2167 3504 2201 3538
rect 2095 3436 2129 3470
rect 2167 3436 2201 3470
rect 2095 3368 2129 3402
rect 2167 3368 2201 3402
rect 2095 3300 2129 3334
rect 2167 3300 2201 3334
rect 2095 3232 2129 3266
rect 2167 3232 2201 3266
rect 2095 3164 2129 3198
rect 2167 3164 2201 3198
rect 2525 4048 2559 4082
rect 2729 4048 2763 4082
rect 2525 3980 2559 4014
rect 2729 3980 2763 4014
rect 2525 3912 2559 3946
rect 2729 3912 2763 3946
rect 2525 3844 2559 3878
rect 2729 3844 2763 3878
rect 2525 3776 2559 3810
rect 2729 3776 2763 3810
rect 2525 3708 2559 3742
rect 2729 3708 2763 3742
rect 2525 3640 2559 3674
rect 2729 3640 2763 3674
rect 2525 3572 2559 3606
rect 2729 3572 2763 3606
rect 2525 3504 2559 3538
rect 2729 3504 2763 3538
rect 2525 3436 2559 3470
rect 2729 3436 2763 3470
rect 2525 3368 2559 3402
rect 2729 3368 2763 3402
rect 2525 3300 2559 3334
rect 2729 3300 2763 3334
rect 2525 3232 2559 3266
rect 2729 3232 2763 3266
rect 2525 3164 2559 3198
rect 2729 3164 2763 3198
rect 3087 4048 3121 4082
rect 3159 4048 3193 4082
rect 3087 3980 3121 4014
rect 3159 3980 3193 4014
rect 3087 3912 3121 3946
rect 3159 3912 3193 3946
rect 3087 3844 3121 3878
rect 3159 3844 3193 3878
rect 3087 3776 3121 3810
rect 3159 3776 3193 3810
rect 3087 3708 3121 3742
rect 3159 3708 3193 3742
rect 3087 3640 3121 3674
rect 3159 3640 3193 3674
rect 3087 3572 3121 3606
rect 3159 3572 3193 3606
rect 3087 3504 3121 3538
rect 3159 3504 3193 3538
rect 3087 3436 3121 3470
rect 3159 3436 3193 3470
rect 3087 3368 3121 3402
rect 3159 3368 3193 3402
rect 3087 3300 3121 3334
rect 3159 3300 3193 3334
rect 3087 3232 3121 3266
rect 3159 3232 3193 3266
rect 3087 3164 3121 3198
rect 3159 3164 3193 3198
rect 3517 4048 3551 4082
rect 3721 4048 3755 4082
rect 3517 3980 3551 4014
rect 3721 3980 3755 4014
rect 3517 3912 3551 3946
rect 3721 3912 3755 3946
rect 3517 3844 3551 3878
rect 3721 3844 3755 3878
rect 3517 3776 3551 3810
rect 3721 3776 3755 3810
rect 3517 3708 3551 3742
rect 3721 3708 3755 3742
rect 3517 3640 3551 3674
rect 3721 3640 3755 3674
rect 3517 3572 3551 3606
rect 3721 3572 3755 3606
rect 3517 3504 3551 3538
rect 3721 3504 3755 3538
rect 3517 3436 3551 3470
rect 3721 3436 3755 3470
rect 3517 3368 3551 3402
rect 3721 3368 3755 3402
rect 3517 3300 3551 3334
rect 3721 3300 3755 3334
rect 3517 3232 3551 3266
rect 3721 3232 3755 3266
rect 3517 3164 3551 3198
rect 3721 3164 3755 3198
rect 4079 4048 4113 4082
rect 4151 4048 4185 4082
rect 4079 3980 4113 4014
rect 4151 3980 4185 4014
rect 4079 3912 4113 3946
rect 4151 3912 4185 3946
rect 4079 3844 4113 3878
rect 4151 3844 4185 3878
rect 4079 3776 4113 3810
rect 4151 3776 4185 3810
rect 4079 3708 4113 3742
rect 4151 3708 4185 3742
rect 4079 3640 4113 3674
rect 4151 3640 4185 3674
rect 4079 3572 4113 3606
rect 4151 3572 4185 3606
rect 4079 3504 4113 3538
rect 4151 3504 4185 3538
rect 4079 3436 4113 3470
rect 4151 3436 4185 3470
rect 4079 3368 4113 3402
rect 4151 3368 4185 3402
rect 4079 3300 4113 3334
rect 4151 3300 4185 3334
rect 4079 3232 4113 3266
rect 4151 3232 4185 3266
rect 4079 3164 4113 3198
rect 4151 3164 4185 3198
rect 4509 4048 4543 4082
rect 4713 4048 4747 4082
rect 4509 3980 4543 4014
rect 4713 3980 4747 4014
rect 4509 3912 4543 3946
rect 4713 3912 4747 3946
rect 4509 3844 4543 3878
rect 4713 3844 4747 3878
rect 4509 3776 4543 3810
rect 4713 3776 4747 3810
rect 4509 3708 4543 3742
rect 4713 3708 4747 3742
rect 4509 3640 4543 3674
rect 4713 3640 4747 3674
rect 4509 3572 4543 3606
rect 4713 3572 4747 3606
rect 4509 3504 4543 3538
rect 4713 3504 4747 3538
rect 4509 3436 4543 3470
rect 4713 3436 4747 3470
rect 4509 3368 4543 3402
rect 4713 3368 4747 3402
rect 4509 3300 4543 3334
rect 4713 3300 4747 3334
rect 4509 3232 4543 3266
rect 4713 3232 4747 3266
rect 4509 3164 4543 3198
rect 4713 3164 4747 3198
rect 5071 4048 5105 4082
rect 5143 4048 5177 4082
rect 5071 3980 5105 4014
rect 5143 3980 5177 4014
rect 5071 3912 5105 3946
rect 5143 3912 5177 3946
rect 5071 3844 5105 3878
rect 5143 3844 5177 3878
rect 5071 3776 5105 3810
rect 5143 3776 5177 3810
rect 5071 3708 5105 3742
rect 5143 3708 5177 3742
rect 5071 3640 5105 3674
rect 5143 3640 5177 3674
rect 5071 3572 5105 3606
rect 5143 3572 5177 3606
rect 5071 3504 5105 3538
rect 5143 3504 5177 3538
rect 5071 3436 5105 3470
rect 5143 3436 5177 3470
rect 5071 3368 5105 3402
rect 5143 3368 5177 3402
rect 5071 3300 5105 3334
rect 5143 3300 5177 3334
rect 5071 3232 5105 3266
rect 5143 3232 5177 3266
rect 5071 3164 5105 3198
rect 5143 3164 5177 3198
rect 5501 4048 5535 4082
rect 5705 4048 5739 4082
rect 5501 3980 5535 4014
rect 5705 3980 5739 4014
rect 5501 3912 5535 3946
rect 5705 3912 5739 3946
rect 5501 3844 5535 3878
rect 5705 3844 5739 3878
rect 5501 3776 5535 3810
rect 5705 3776 5739 3810
rect 5501 3708 5535 3742
rect 5705 3708 5739 3742
rect 5501 3640 5535 3674
rect 5705 3640 5739 3674
rect 5501 3572 5535 3606
rect 5705 3572 5739 3606
rect 5501 3504 5535 3538
rect 5705 3504 5739 3538
rect 5501 3436 5535 3470
rect 5705 3436 5739 3470
rect 5501 3368 5535 3402
rect 5705 3368 5739 3402
rect 5501 3300 5535 3334
rect 5705 3300 5739 3334
rect 5501 3232 5535 3266
rect 5705 3232 5739 3266
rect 5501 3164 5535 3198
rect 5705 3164 5739 3198
rect 6063 4048 6097 4082
rect 6135 4048 6169 4082
rect 6063 3980 6097 4014
rect 6135 3980 6169 4014
rect 6063 3912 6097 3946
rect 6135 3912 6169 3946
rect 6063 3844 6097 3878
rect 6135 3844 6169 3878
rect 6063 3776 6097 3810
rect 6135 3776 6169 3810
rect 6063 3708 6097 3742
rect 6135 3708 6169 3742
rect 6063 3640 6097 3674
rect 6135 3640 6169 3674
rect 6063 3572 6097 3606
rect 6135 3572 6169 3606
rect 6063 3504 6097 3538
rect 6135 3504 6169 3538
rect 6063 3436 6097 3470
rect 6135 3436 6169 3470
rect 6063 3368 6097 3402
rect 6135 3368 6169 3402
rect 6063 3300 6097 3334
rect 6135 3300 6169 3334
rect 6063 3232 6097 3266
rect 6135 3232 6169 3266
rect 6063 3164 6097 3198
rect 6135 3164 6169 3198
rect 6493 4048 6527 4082
rect 6697 4048 6731 4082
rect 6493 3980 6527 4014
rect 6697 3980 6731 4014
rect 6493 3912 6527 3946
rect 6697 3912 6731 3946
rect 6493 3844 6527 3878
rect 6697 3844 6731 3878
rect 6493 3776 6527 3810
rect 6697 3776 6731 3810
rect 6493 3708 6527 3742
rect 6697 3708 6731 3742
rect 6493 3640 6527 3674
rect 6697 3640 6731 3674
rect 6493 3572 6527 3606
rect 6697 3572 6731 3606
rect 6493 3504 6527 3538
rect 6697 3504 6731 3538
rect 6493 3436 6527 3470
rect 6697 3436 6731 3470
rect 6493 3368 6527 3402
rect 6697 3368 6731 3402
rect 6493 3300 6527 3334
rect 6697 3300 6731 3334
rect 6493 3232 6527 3266
rect 6697 3232 6731 3266
rect 6493 3164 6527 3198
rect 6697 3164 6731 3198
rect 7055 4048 7089 4082
rect 7127 4048 7161 4082
rect 7055 3980 7089 4014
rect 7127 3980 7161 4014
rect 7055 3912 7089 3946
rect 7127 3912 7161 3946
rect 7055 3844 7089 3878
rect 7127 3844 7161 3878
rect 7055 3776 7089 3810
rect 7127 3776 7161 3810
rect 7055 3708 7089 3742
rect 7127 3708 7161 3742
rect 7055 3640 7089 3674
rect 7127 3640 7161 3674
rect 7055 3572 7089 3606
rect 7127 3572 7161 3606
rect 7055 3504 7089 3538
rect 7127 3504 7161 3538
rect 7055 3436 7089 3470
rect 7127 3436 7161 3470
rect 7055 3368 7089 3402
rect 7127 3368 7161 3402
rect 7055 3300 7089 3334
rect 7127 3300 7161 3334
rect 7055 3232 7089 3266
rect 7127 3232 7161 3266
rect 7055 3164 7089 3198
rect 7127 3164 7161 3198
rect 7485 4048 7519 4082
rect 7689 4048 7723 4082
rect 7485 3980 7519 4014
rect 7689 3980 7723 4014
rect 7485 3912 7519 3946
rect 7689 3912 7723 3946
rect 7485 3844 7519 3878
rect 7689 3844 7723 3878
rect 7485 3776 7519 3810
rect 7689 3776 7723 3810
rect 7485 3708 7519 3742
rect 7689 3708 7723 3742
rect 7485 3640 7519 3674
rect 7689 3640 7723 3674
rect 7485 3572 7519 3606
rect 7689 3572 7723 3606
rect 7485 3504 7519 3538
rect 7689 3504 7723 3538
rect 7485 3436 7519 3470
rect 7689 3436 7723 3470
rect 7485 3368 7519 3402
rect 7689 3368 7723 3402
rect 7485 3300 7519 3334
rect 7689 3300 7723 3334
rect 7485 3232 7519 3266
rect 7689 3232 7723 3266
rect 7485 3164 7519 3198
rect 7689 3164 7723 3198
rect 8047 4048 8081 4082
rect 8119 4048 8153 4082
rect 8047 3980 8081 4014
rect 8119 3980 8153 4014
rect 8047 3912 8081 3946
rect 8119 3912 8153 3946
rect 8047 3844 8081 3878
rect 8119 3844 8153 3878
rect 8047 3776 8081 3810
rect 8119 3776 8153 3810
rect 8047 3708 8081 3742
rect 8119 3708 8153 3742
rect 8047 3640 8081 3674
rect 8119 3640 8153 3674
rect 8047 3572 8081 3606
rect 8119 3572 8153 3606
rect 8047 3504 8081 3538
rect 8119 3504 8153 3538
rect 8047 3436 8081 3470
rect 8119 3436 8153 3470
rect 8047 3368 8081 3402
rect 8119 3368 8153 3402
rect 8047 3300 8081 3334
rect 8119 3300 8153 3334
rect 8047 3232 8081 3266
rect 8119 3232 8153 3266
rect 8047 3164 8081 3198
rect 8119 3164 8153 3198
rect 8477 4048 8511 4082
rect 8681 4048 8715 4082
rect 8477 3980 8511 4014
rect 8681 3980 8715 4014
rect 8477 3912 8511 3946
rect 8681 3912 8715 3946
rect 8477 3844 8511 3878
rect 8681 3844 8715 3878
rect 8477 3776 8511 3810
rect 8681 3776 8715 3810
rect 8477 3708 8511 3742
rect 8681 3708 8715 3742
rect 8477 3640 8511 3674
rect 8681 3640 8715 3674
rect 8477 3572 8511 3606
rect 8681 3572 8715 3606
rect 8477 3504 8511 3538
rect 8681 3504 8715 3538
rect 8477 3436 8511 3470
rect 8681 3436 8715 3470
rect 8477 3368 8511 3402
rect 8681 3368 8715 3402
rect 8477 3300 8511 3334
rect 8681 3300 8715 3334
rect 8477 3232 8511 3266
rect 8681 3232 8715 3266
rect 8477 3164 8511 3198
rect 8681 3164 8715 3198
rect 9039 4048 9073 4082
rect 9111 4048 9145 4082
rect 9039 3980 9073 4014
rect 9111 3980 9145 4014
rect 9039 3912 9073 3946
rect 9111 3912 9145 3946
rect 9039 3844 9073 3878
rect 9111 3844 9145 3878
rect 9039 3776 9073 3810
rect 9111 3776 9145 3810
rect 9039 3708 9073 3742
rect 9111 3708 9145 3742
rect 9039 3640 9073 3674
rect 9111 3640 9145 3674
rect 9039 3572 9073 3606
rect 9111 3572 9145 3606
rect 9039 3504 9073 3538
rect 9111 3504 9145 3538
rect 9039 3436 9073 3470
rect 9111 3436 9145 3470
rect 9039 3368 9073 3402
rect 9111 3368 9145 3402
rect 9039 3300 9073 3334
rect 9111 3300 9145 3334
rect 9039 3232 9073 3266
rect 9111 3232 9145 3266
rect 9039 3164 9073 3198
rect 9111 3164 9145 3198
rect 9469 4048 9503 4082
rect 9673 4048 9707 4082
rect 9469 3980 9503 4014
rect 9673 3980 9707 4014
rect 9469 3912 9503 3946
rect 9673 3912 9707 3946
rect 9469 3844 9503 3878
rect 9673 3844 9707 3878
rect 9469 3776 9503 3810
rect 9673 3776 9707 3810
rect 9469 3708 9503 3742
rect 9673 3708 9707 3742
rect 9469 3640 9503 3674
rect 9673 3640 9707 3674
rect 9469 3572 9503 3606
rect 9673 3572 9707 3606
rect 9469 3504 9503 3538
rect 9673 3504 9707 3538
rect 9469 3436 9503 3470
rect 9673 3436 9707 3470
rect 9469 3368 9503 3402
rect 9673 3368 9707 3402
rect 9469 3300 9503 3334
rect 9673 3300 9707 3334
rect 9469 3232 9503 3266
rect 9673 3232 9707 3266
rect 9469 3164 9503 3198
rect 9673 3164 9707 3198
rect 10031 4048 10065 4082
rect 10103 4048 10137 4082
rect 10031 3980 10065 4014
rect 10103 3980 10137 4014
rect 10031 3912 10065 3946
rect 10103 3912 10137 3946
rect 10031 3844 10065 3878
rect 10103 3844 10137 3878
rect 10031 3776 10065 3810
rect 10103 3776 10137 3810
rect 10031 3708 10065 3742
rect 10103 3708 10137 3742
rect 10031 3640 10065 3674
rect 10103 3640 10137 3674
rect 10031 3572 10065 3606
rect 10103 3572 10137 3606
rect 10031 3504 10065 3538
rect 10103 3504 10137 3538
rect 10031 3436 10065 3470
rect 10103 3436 10137 3470
rect 10031 3368 10065 3402
rect 10103 3368 10137 3402
rect 10031 3300 10065 3334
rect 10103 3300 10137 3334
rect 10031 3232 10065 3266
rect 10103 3232 10137 3266
rect 10031 3164 10065 3198
rect 10103 3164 10137 3198
rect 10461 4048 10495 4082
rect 10665 4048 10699 4082
rect 10461 3980 10495 4014
rect 10665 3980 10699 4014
rect 10461 3912 10495 3946
rect 10665 3912 10699 3946
rect 10461 3844 10495 3878
rect 10665 3844 10699 3878
rect 10461 3776 10495 3810
rect 10665 3776 10699 3810
rect 10461 3708 10495 3742
rect 10665 3708 10699 3742
rect 10461 3640 10495 3674
rect 10665 3640 10699 3674
rect 10461 3572 10495 3606
rect 10665 3572 10699 3606
rect 10461 3504 10495 3538
rect 10665 3504 10699 3538
rect 10461 3436 10495 3470
rect 10665 3436 10699 3470
rect 10461 3368 10495 3402
rect 10665 3368 10699 3402
rect 10461 3300 10495 3334
rect 10665 3300 10699 3334
rect 10461 3232 10495 3266
rect 10665 3232 10699 3266
rect 10461 3164 10495 3198
rect 10665 3164 10699 3198
rect 11023 4048 11057 4082
rect 11095 4048 11129 4082
rect 11023 3980 11057 4014
rect 11095 3980 11129 4014
rect 11023 3912 11057 3946
rect 11095 3912 11129 3946
rect 11023 3844 11057 3878
rect 11095 3844 11129 3878
rect 11023 3776 11057 3810
rect 11095 3776 11129 3810
rect 11023 3708 11057 3742
rect 11095 3708 11129 3742
rect 11023 3640 11057 3674
rect 11095 3640 11129 3674
rect 11023 3572 11057 3606
rect 11095 3572 11129 3606
rect 11023 3504 11057 3538
rect 11095 3504 11129 3538
rect 11023 3436 11057 3470
rect 11095 3436 11129 3470
rect 11023 3368 11057 3402
rect 11095 3368 11129 3402
rect 11023 3300 11057 3334
rect 11095 3300 11129 3334
rect 11023 3232 11057 3266
rect 11095 3232 11129 3266
rect 11023 3164 11057 3198
rect 11095 3164 11129 3198
rect 11453 4048 11487 4082
rect 11657 4048 11691 4082
rect 11453 3980 11487 4014
rect 11657 3980 11691 4014
rect 11453 3912 11487 3946
rect 11657 3912 11691 3946
rect 11453 3844 11487 3878
rect 11657 3844 11691 3878
rect 11453 3776 11487 3810
rect 11657 3776 11691 3810
rect 11453 3708 11487 3742
rect 11657 3708 11691 3742
rect 11453 3640 11487 3674
rect 11657 3640 11691 3674
rect 11453 3572 11487 3606
rect 11657 3572 11691 3606
rect 11453 3504 11487 3538
rect 11657 3504 11691 3538
rect 11453 3436 11487 3470
rect 11657 3436 11691 3470
rect 11453 3368 11487 3402
rect 11657 3368 11691 3402
rect 11453 3300 11487 3334
rect 11657 3300 11691 3334
rect 11453 3232 11487 3266
rect 11657 3232 11691 3266
rect 11453 3164 11487 3198
rect 11657 3164 11691 3198
rect 12015 4048 12049 4082
rect 12087 4048 12121 4082
rect 12015 3980 12049 4014
rect 12087 3980 12121 4014
rect 12015 3912 12049 3946
rect 12087 3912 12121 3946
rect 12015 3844 12049 3878
rect 12087 3844 12121 3878
rect 12015 3776 12049 3810
rect 12087 3776 12121 3810
rect 12015 3708 12049 3742
rect 12087 3708 12121 3742
rect 12015 3640 12049 3674
rect 12087 3640 12121 3674
rect 12015 3572 12049 3606
rect 12087 3572 12121 3606
rect 12015 3504 12049 3538
rect 12087 3504 12121 3538
rect 12015 3436 12049 3470
rect 12087 3436 12121 3470
rect 12015 3368 12049 3402
rect 12087 3368 12121 3402
rect 12015 3300 12049 3334
rect 12087 3300 12121 3334
rect 12015 3232 12049 3266
rect 12087 3232 12121 3266
rect 12015 3164 12049 3198
rect 12087 3164 12121 3198
rect 12445 4048 12479 4082
rect 12649 4048 12683 4082
rect 12445 3980 12479 4014
rect 12649 3980 12683 4014
rect 12445 3912 12479 3946
rect 12649 3912 12683 3946
rect 12445 3844 12479 3878
rect 12649 3844 12683 3878
rect 12445 3776 12479 3810
rect 12649 3776 12683 3810
rect 12445 3708 12479 3742
rect 12649 3708 12683 3742
rect 12445 3640 12479 3674
rect 12649 3640 12683 3674
rect 12445 3572 12479 3606
rect 12649 3572 12683 3606
rect 12445 3504 12479 3538
rect 12649 3504 12683 3538
rect 12445 3436 12479 3470
rect 12649 3436 12683 3470
rect 12445 3368 12479 3402
rect 12649 3368 12683 3402
rect 12445 3300 12479 3334
rect 12649 3300 12683 3334
rect 12445 3232 12479 3266
rect 12649 3232 12683 3266
rect 12445 3164 12479 3198
rect 12649 3164 12683 3198
rect 13007 4048 13041 4082
rect 13079 4048 13113 4082
rect 13007 3980 13041 4014
rect 13079 3980 13113 4014
rect 13007 3912 13041 3946
rect 13079 3912 13113 3946
rect 13007 3844 13041 3878
rect 13079 3844 13113 3878
rect 13007 3776 13041 3810
rect 13079 3776 13113 3810
rect 13007 3708 13041 3742
rect 13079 3708 13113 3742
rect 13007 3640 13041 3674
rect 13079 3640 13113 3674
rect 13007 3572 13041 3606
rect 13079 3572 13113 3606
rect 13007 3504 13041 3538
rect 13079 3504 13113 3538
rect 13007 3436 13041 3470
rect 13079 3436 13113 3470
rect 13007 3368 13041 3402
rect 13079 3368 13113 3402
rect 13007 3300 13041 3334
rect 13079 3300 13113 3334
rect 13007 3232 13041 3266
rect 13079 3232 13113 3266
rect 13007 3164 13041 3198
rect 13079 3164 13113 3198
rect 13437 4048 13471 4082
rect 13641 4048 13675 4082
rect 13437 3980 13471 4014
rect 13641 3980 13675 4014
rect 13437 3912 13471 3946
rect 13641 3912 13675 3946
rect 13437 3844 13471 3878
rect 13641 3844 13675 3878
rect 13437 3776 13471 3810
rect 13641 3776 13675 3810
rect 13437 3708 13471 3742
rect 13641 3708 13675 3742
rect 13437 3640 13471 3674
rect 13641 3640 13675 3674
rect 13437 3572 13471 3606
rect 13641 3572 13675 3606
rect 13437 3504 13471 3538
rect 13641 3504 13675 3538
rect 13437 3436 13471 3470
rect 13641 3436 13675 3470
rect 13437 3368 13471 3402
rect 13641 3368 13675 3402
rect 13437 3300 13471 3334
rect 13641 3300 13675 3334
rect 13437 3232 13471 3266
rect 13641 3232 13675 3266
rect 13437 3164 13471 3198
rect 13641 3164 13675 3198
rect 13999 4048 14033 4082
rect 13999 3980 14033 4014
rect 13999 3912 14033 3946
rect 13999 3844 14033 3878
rect 13999 3776 14033 3810
rect 13999 3708 14033 3742
rect 13999 3640 14033 3674
rect 13999 3572 14033 3606
rect 13999 3504 14033 3538
rect 13999 3436 14033 3470
rect 13999 3368 14033 3402
rect 13999 3300 14033 3334
rect 13999 3232 14033 3266
rect 13999 3164 14033 3198
rect 14356 4048 14390 4082
rect 14356 3980 14390 4014
rect 14356 3912 14390 3946
rect 14356 3844 14390 3878
rect 14356 3776 14390 3810
rect 14356 3708 14390 3742
rect 14356 3640 14390 3674
rect 14356 3572 14390 3606
rect 14356 3504 14390 3538
rect 14356 3436 14390 3470
rect 14356 3368 14390 3402
rect 14356 3300 14390 3334
rect 14356 3232 14390 3266
rect 14356 3164 14390 3198
rect 745 2448 779 2482
rect 745 2380 779 2414
rect 745 2312 779 2346
rect 745 2244 779 2278
rect 745 2176 779 2210
rect 745 2108 779 2142
rect 745 2040 779 2074
rect 745 1972 779 2006
rect 745 1904 779 1938
rect 745 1836 779 1870
rect 745 1768 779 1802
rect 745 1700 779 1734
rect 745 1632 779 1666
rect 745 1564 779 1598
rect 1103 2448 1137 2482
rect 1175 2448 1209 2482
rect 1103 2380 1137 2414
rect 1175 2380 1209 2414
rect 1103 2312 1137 2346
rect 1175 2312 1209 2346
rect 1103 2244 1137 2278
rect 1175 2244 1209 2278
rect 1103 2176 1137 2210
rect 1175 2176 1209 2210
rect 1103 2108 1137 2142
rect 1175 2108 1209 2142
rect 1103 2040 1137 2074
rect 1175 2040 1209 2074
rect 1103 1972 1137 2006
rect 1175 1972 1209 2006
rect 1103 1904 1137 1938
rect 1175 1904 1209 1938
rect 1103 1836 1137 1870
rect 1175 1836 1209 1870
rect 1103 1768 1137 1802
rect 1175 1768 1209 1802
rect 1103 1700 1137 1734
rect 1175 1700 1209 1734
rect 1103 1632 1137 1666
rect 1175 1632 1209 1666
rect 1103 1564 1137 1598
rect 1175 1564 1209 1598
rect 1533 2506 1567 2540
rect 1737 2506 1771 2540
rect 1533 2438 1567 2472
rect 1737 2438 1771 2472
rect 1533 2370 1567 2404
rect 1737 2370 1771 2404
rect 1533 2302 1567 2336
rect 1737 2302 1771 2336
rect 1533 2234 1567 2268
rect 1737 2234 1771 2268
rect 1533 2166 1567 2200
rect 1737 2166 1771 2200
rect 1533 2098 1567 2132
rect 1737 2098 1771 2132
rect 1533 2030 1567 2064
rect 1737 2030 1771 2064
rect 1533 1962 1567 1996
rect 1737 1962 1771 1996
rect 1533 1894 1567 1928
rect 1737 1894 1771 1928
rect 1533 1826 1567 1860
rect 1737 1826 1771 1860
rect 1533 1758 1567 1792
rect 1737 1758 1771 1792
rect 1533 1690 1567 1724
rect 1737 1690 1771 1724
rect 1533 1622 1567 1656
rect 1737 1622 1771 1656
rect 2095 2448 2129 2482
rect 2167 2448 2201 2482
rect 2095 2380 2129 2414
rect 2167 2380 2201 2414
rect 2095 2312 2129 2346
rect 2167 2312 2201 2346
rect 2095 2244 2129 2278
rect 2167 2244 2201 2278
rect 2095 2176 2129 2210
rect 2167 2176 2201 2210
rect 2095 2108 2129 2142
rect 2167 2108 2201 2142
rect 2095 2040 2129 2074
rect 2167 2040 2201 2074
rect 2095 1972 2129 2006
rect 2167 1972 2201 2006
rect 2095 1904 2129 1938
rect 2167 1904 2201 1938
rect 2095 1836 2129 1870
rect 2167 1836 2201 1870
rect 2095 1768 2129 1802
rect 2167 1768 2201 1802
rect 2095 1700 2129 1734
rect 2167 1700 2201 1734
rect 2095 1632 2129 1666
rect 2167 1632 2201 1666
rect 2095 1564 2129 1598
rect 2167 1564 2201 1598
rect 2525 2506 2559 2540
rect 2729 2506 2763 2540
rect 2525 2438 2559 2472
rect 2729 2438 2763 2472
rect 2525 2370 2559 2404
rect 2729 2370 2763 2404
rect 2525 2302 2559 2336
rect 2729 2302 2763 2336
rect 2525 2234 2559 2268
rect 2729 2234 2763 2268
rect 2525 2166 2559 2200
rect 2729 2166 2763 2200
rect 2525 2098 2559 2132
rect 2729 2098 2763 2132
rect 2525 2030 2559 2064
rect 2729 2030 2763 2064
rect 2525 1962 2559 1996
rect 2729 1962 2763 1996
rect 2525 1894 2559 1928
rect 2729 1894 2763 1928
rect 2525 1826 2559 1860
rect 2729 1826 2763 1860
rect 2525 1758 2559 1792
rect 2729 1758 2763 1792
rect 2525 1690 2559 1724
rect 2729 1690 2763 1724
rect 2525 1622 2559 1656
rect 2729 1622 2763 1656
rect 3087 2448 3121 2482
rect 3159 2448 3193 2482
rect 3087 2380 3121 2414
rect 3159 2380 3193 2414
rect 3087 2312 3121 2346
rect 3159 2312 3193 2346
rect 3087 2244 3121 2278
rect 3159 2244 3193 2278
rect 3087 2176 3121 2210
rect 3159 2176 3193 2210
rect 3087 2108 3121 2142
rect 3159 2108 3193 2142
rect 3087 2040 3121 2074
rect 3159 2040 3193 2074
rect 3087 1972 3121 2006
rect 3159 1972 3193 2006
rect 3087 1904 3121 1938
rect 3159 1904 3193 1938
rect 3087 1836 3121 1870
rect 3159 1836 3193 1870
rect 3087 1768 3121 1802
rect 3159 1768 3193 1802
rect 3087 1700 3121 1734
rect 3159 1700 3193 1734
rect 3087 1632 3121 1666
rect 3159 1632 3193 1666
rect 3087 1564 3121 1598
rect 3159 1564 3193 1598
rect 3517 2506 3551 2540
rect 3721 2506 3755 2540
rect 3517 2438 3551 2472
rect 3721 2438 3755 2472
rect 3517 2370 3551 2404
rect 3721 2370 3755 2404
rect 3517 2302 3551 2336
rect 3721 2302 3755 2336
rect 3517 2234 3551 2268
rect 3721 2234 3755 2268
rect 3517 2166 3551 2200
rect 3721 2166 3755 2200
rect 3517 2098 3551 2132
rect 3721 2098 3755 2132
rect 3517 2030 3551 2064
rect 3721 2030 3755 2064
rect 3517 1962 3551 1996
rect 3721 1962 3755 1996
rect 3517 1894 3551 1928
rect 3721 1894 3755 1928
rect 3517 1826 3551 1860
rect 3721 1826 3755 1860
rect 3517 1758 3551 1792
rect 3721 1758 3755 1792
rect 3517 1690 3551 1724
rect 3721 1690 3755 1724
rect 3517 1622 3551 1656
rect 3721 1622 3755 1656
rect 4079 2448 4113 2482
rect 4151 2448 4185 2482
rect 4079 2380 4113 2414
rect 4151 2380 4185 2414
rect 4079 2312 4113 2346
rect 4151 2312 4185 2346
rect 4079 2244 4113 2278
rect 4151 2244 4185 2278
rect 4079 2176 4113 2210
rect 4151 2176 4185 2210
rect 4079 2108 4113 2142
rect 4151 2108 4185 2142
rect 4079 2040 4113 2074
rect 4151 2040 4185 2074
rect 4079 1972 4113 2006
rect 4151 1972 4185 2006
rect 4079 1904 4113 1938
rect 4151 1904 4185 1938
rect 4079 1836 4113 1870
rect 4151 1836 4185 1870
rect 4079 1768 4113 1802
rect 4151 1768 4185 1802
rect 4079 1700 4113 1734
rect 4151 1700 4185 1734
rect 4079 1632 4113 1666
rect 4151 1632 4185 1666
rect 4079 1564 4113 1598
rect 4151 1564 4185 1598
rect 4509 2506 4543 2540
rect 4713 2506 4747 2540
rect 4509 2438 4543 2472
rect 4713 2438 4747 2472
rect 4509 2370 4543 2404
rect 4713 2370 4747 2404
rect 4509 2302 4543 2336
rect 4713 2302 4747 2336
rect 4509 2234 4543 2268
rect 4713 2234 4747 2268
rect 4509 2166 4543 2200
rect 4713 2166 4747 2200
rect 4509 2098 4543 2132
rect 4713 2098 4747 2132
rect 4509 2030 4543 2064
rect 4713 2030 4747 2064
rect 4509 1962 4543 1996
rect 4713 1962 4747 1996
rect 4509 1894 4543 1928
rect 4713 1894 4747 1928
rect 4509 1826 4543 1860
rect 4713 1826 4747 1860
rect 4509 1758 4543 1792
rect 4713 1758 4747 1792
rect 4509 1690 4543 1724
rect 4713 1690 4747 1724
rect 4509 1622 4543 1656
rect 4713 1622 4747 1656
rect 5071 2448 5105 2482
rect 5143 2448 5177 2482
rect 5071 2380 5105 2414
rect 5143 2380 5177 2414
rect 5071 2312 5105 2346
rect 5143 2312 5177 2346
rect 5071 2244 5105 2278
rect 5143 2244 5177 2278
rect 5071 2176 5105 2210
rect 5143 2176 5177 2210
rect 5071 2108 5105 2142
rect 5143 2108 5177 2142
rect 5071 2040 5105 2074
rect 5143 2040 5177 2074
rect 5071 1972 5105 2006
rect 5143 1972 5177 2006
rect 5071 1904 5105 1938
rect 5143 1904 5177 1938
rect 5071 1836 5105 1870
rect 5143 1836 5177 1870
rect 5071 1768 5105 1802
rect 5143 1768 5177 1802
rect 5071 1700 5105 1734
rect 5143 1700 5177 1734
rect 5071 1632 5105 1666
rect 5143 1632 5177 1666
rect 5071 1564 5105 1598
rect 5143 1564 5177 1598
rect 5501 2506 5535 2540
rect 5705 2506 5739 2540
rect 5501 2438 5535 2472
rect 5705 2438 5739 2472
rect 5501 2370 5535 2404
rect 5705 2370 5739 2404
rect 5501 2302 5535 2336
rect 5705 2302 5739 2336
rect 5501 2234 5535 2268
rect 5705 2234 5739 2268
rect 5501 2166 5535 2200
rect 5705 2166 5739 2200
rect 5501 2098 5535 2132
rect 5705 2098 5739 2132
rect 5501 2030 5535 2064
rect 5705 2030 5739 2064
rect 5501 1962 5535 1996
rect 5705 1962 5739 1996
rect 5501 1894 5535 1928
rect 5705 1894 5739 1928
rect 5501 1826 5535 1860
rect 5705 1826 5739 1860
rect 5501 1758 5535 1792
rect 5705 1758 5739 1792
rect 5501 1690 5535 1724
rect 5705 1690 5739 1724
rect 5501 1622 5535 1656
rect 5705 1622 5739 1656
rect 6063 2448 6097 2482
rect 6135 2448 6169 2482
rect 6063 2380 6097 2414
rect 6135 2380 6169 2414
rect 6063 2312 6097 2346
rect 6135 2312 6169 2346
rect 6063 2244 6097 2278
rect 6135 2244 6169 2278
rect 6063 2176 6097 2210
rect 6135 2176 6169 2210
rect 6063 2108 6097 2142
rect 6135 2108 6169 2142
rect 6063 2040 6097 2074
rect 6135 2040 6169 2074
rect 6063 1972 6097 2006
rect 6135 1972 6169 2006
rect 6063 1904 6097 1938
rect 6135 1904 6169 1938
rect 6063 1836 6097 1870
rect 6135 1836 6169 1870
rect 6063 1768 6097 1802
rect 6135 1768 6169 1802
rect 6063 1700 6097 1734
rect 6135 1700 6169 1734
rect 6063 1632 6097 1666
rect 6135 1632 6169 1666
rect 6063 1564 6097 1598
rect 6135 1564 6169 1598
rect 6493 2506 6527 2540
rect 6697 2506 6731 2540
rect 6493 2438 6527 2472
rect 6697 2438 6731 2472
rect 6493 2370 6527 2404
rect 6697 2370 6731 2404
rect 6493 2302 6527 2336
rect 6697 2302 6731 2336
rect 6493 2234 6527 2268
rect 6697 2234 6731 2268
rect 6493 2166 6527 2200
rect 6697 2166 6731 2200
rect 6493 2098 6527 2132
rect 6697 2098 6731 2132
rect 6493 2030 6527 2064
rect 6697 2030 6731 2064
rect 6493 1962 6527 1996
rect 6697 1962 6731 1996
rect 6493 1894 6527 1928
rect 6697 1894 6731 1928
rect 6493 1826 6527 1860
rect 6697 1826 6731 1860
rect 6493 1758 6527 1792
rect 6697 1758 6731 1792
rect 6493 1690 6527 1724
rect 6697 1690 6731 1724
rect 6493 1622 6527 1656
rect 6697 1622 6731 1656
rect 7055 2448 7089 2482
rect 7127 2448 7161 2482
rect 7055 2380 7089 2414
rect 7127 2380 7161 2414
rect 7055 2312 7089 2346
rect 7127 2312 7161 2346
rect 7055 2244 7089 2278
rect 7127 2244 7161 2278
rect 7055 2176 7089 2210
rect 7127 2176 7161 2210
rect 7055 2108 7089 2142
rect 7127 2108 7161 2142
rect 7055 2040 7089 2074
rect 7127 2040 7161 2074
rect 7055 1972 7089 2006
rect 7127 1972 7161 2006
rect 7055 1904 7089 1938
rect 7127 1904 7161 1938
rect 7055 1836 7089 1870
rect 7127 1836 7161 1870
rect 7055 1768 7089 1802
rect 7127 1768 7161 1802
rect 7055 1700 7089 1734
rect 7127 1700 7161 1734
rect 7055 1632 7089 1666
rect 7127 1632 7161 1666
rect 7055 1564 7089 1598
rect 7127 1564 7161 1598
rect 7485 2506 7519 2540
rect 7689 2506 7723 2540
rect 7485 2438 7519 2472
rect 7689 2438 7723 2472
rect 7485 2370 7519 2404
rect 7689 2370 7723 2404
rect 7485 2302 7519 2336
rect 7689 2302 7723 2336
rect 7485 2234 7519 2268
rect 7689 2234 7723 2268
rect 7485 2166 7519 2200
rect 7689 2166 7723 2200
rect 7485 2098 7519 2132
rect 7689 2098 7723 2132
rect 7485 2030 7519 2064
rect 7689 2030 7723 2064
rect 7485 1962 7519 1996
rect 7689 1962 7723 1996
rect 7485 1894 7519 1928
rect 7689 1894 7723 1928
rect 7485 1826 7519 1860
rect 7689 1826 7723 1860
rect 7485 1758 7519 1792
rect 7689 1758 7723 1792
rect 7485 1690 7519 1724
rect 7689 1690 7723 1724
rect 7485 1622 7519 1656
rect 7689 1622 7723 1656
rect 8047 2448 8081 2482
rect 8119 2448 8153 2482
rect 8047 2380 8081 2414
rect 8119 2380 8153 2414
rect 8047 2312 8081 2346
rect 8119 2312 8153 2346
rect 8047 2244 8081 2278
rect 8119 2244 8153 2278
rect 8047 2176 8081 2210
rect 8119 2176 8153 2210
rect 8047 2108 8081 2142
rect 8119 2108 8153 2142
rect 8047 2040 8081 2074
rect 8119 2040 8153 2074
rect 8047 1972 8081 2006
rect 8119 1972 8153 2006
rect 8047 1904 8081 1938
rect 8119 1904 8153 1938
rect 8047 1836 8081 1870
rect 8119 1836 8153 1870
rect 8047 1768 8081 1802
rect 8119 1768 8153 1802
rect 8047 1700 8081 1734
rect 8119 1700 8153 1734
rect 8047 1632 8081 1666
rect 8119 1632 8153 1666
rect 8047 1564 8081 1598
rect 8119 1564 8153 1598
rect 8477 2506 8511 2540
rect 8681 2506 8715 2540
rect 8477 2438 8511 2472
rect 8681 2438 8715 2472
rect 8477 2370 8511 2404
rect 8681 2370 8715 2404
rect 8477 2302 8511 2336
rect 8681 2302 8715 2336
rect 8477 2234 8511 2268
rect 8681 2234 8715 2268
rect 8477 2166 8511 2200
rect 8681 2166 8715 2200
rect 8477 2098 8511 2132
rect 8681 2098 8715 2132
rect 8477 2030 8511 2064
rect 8681 2030 8715 2064
rect 8477 1962 8511 1996
rect 8681 1962 8715 1996
rect 8477 1894 8511 1928
rect 8681 1894 8715 1928
rect 8477 1826 8511 1860
rect 8681 1826 8715 1860
rect 8477 1758 8511 1792
rect 8681 1758 8715 1792
rect 8477 1690 8511 1724
rect 8681 1690 8715 1724
rect 8477 1622 8511 1656
rect 8681 1622 8715 1656
rect 9039 2448 9073 2482
rect 9111 2448 9145 2482
rect 9039 2380 9073 2414
rect 9111 2380 9145 2414
rect 9039 2312 9073 2346
rect 9111 2312 9145 2346
rect 9039 2244 9073 2278
rect 9111 2244 9145 2278
rect 9039 2176 9073 2210
rect 9111 2176 9145 2210
rect 9039 2108 9073 2142
rect 9111 2108 9145 2142
rect 9039 2040 9073 2074
rect 9111 2040 9145 2074
rect 9039 1972 9073 2006
rect 9111 1972 9145 2006
rect 9039 1904 9073 1938
rect 9111 1904 9145 1938
rect 9039 1836 9073 1870
rect 9111 1836 9145 1870
rect 9039 1768 9073 1802
rect 9111 1768 9145 1802
rect 9039 1700 9073 1734
rect 9111 1700 9145 1734
rect 9039 1632 9073 1666
rect 9111 1632 9145 1666
rect 9039 1564 9073 1598
rect 9111 1564 9145 1598
rect 9469 2506 9503 2540
rect 9673 2506 9707 2540
rect 9469 2438 9503 2472
rect 9673 2438 9707 2472
rect 9469 2370 9503 2404
rect 9673 2370 9707 2404
rect 9469 2302 9503 2336
rect 9673 2302 9707 2336
rect 9469 2234 9503 2268
rect 9673 2234 9707 2268
rect 9469 2166 9503 2200
rect 9673 2166 9707 2200
rect 9469 2098 9503 2132
rect 9673 2098 9707 2132
rect 9469 2030 9503 2064
rect 9673 2030 9707 2064
rect 9469 1962 9503 1996
rect 9673 1962 9707 1996
rect 9469 1894 9503 1928
rect 9673 1894 9707 1928
rect 9469 1826 9503 1860
rect 9673 1826 9707 1860
rect 9469 1758 9503 1792
rect 9673 1758 9707 1792
rect 9469 1690 9503 1724
rect 9673 1690 9707 1724
rect 9469 1622 9503 1656
rect 9673 1622 9707 1656
rect 10031 2448 10065 2482
rect 10103 2448 10137 2482
rect 10031 2380 10065 2414
rect 10103 2380 10137 2414
rect 10031 2312 10065 2346
rect 10103 2312 10137 2346
rect 10031 2244 10065 2278
rect 10103 2244 10137 2278
rect 10031 2176 10065 2210
rect 10103 2176 10137 2210
rect 10031 2108 10065 2142
rect 10103 2108 10137 2142
rect 10031 2040 10065 2074
rect 10103 2040 10137 2074
rect 10031 1972 10065 2006
rect 10103 1972 10137 2006
rect 10031 1904 10065 1938
rect 10103 1904 10137 1938
rect 10031 1836 10065 1870
rect 10103 1836 10137 1870
rect 10031 1768 10065 1802
rect 10103 1768 10137 1802
rect 10031 1700 10065 1734
rect 10103 1700 10137 1734
rect 10031 1632 10065 1666
rect 10103 1632 10137 1666
rect 10031 1564 10065 1598
rect 10103 1564 10137 1598
rect 10461 2506 10495 2540
rect 10665 2506 10699 2540
rect 10461 2438 10495 2472
rect 10665 2438 10699 2472
rect 10461 2370 10495 2404
rect 10665 2370 10699 2404
rect 10461 2302 10495 2336
rect 10665 2302 10699 2336
rect 10461 2234 10495 2268
rect 10665 2234 10699 2268
rect 10461 2166 10495 2200
rect 10665 2166 10699 2200
rect 10461 2098 10495 2132
rect 10665 2098 10699 2132
rect 10461 2030 10495 2064
rect 10665 2030 10699 2064
rect 10461 1962 10495 1996
rect 10665 1962 10699 1996
rect 10461 1894 10495 1928
rect 10665 1894 10699 1928
rect 10461 1826 10495 1860
rect 10665 1826 10699 1860
rect 10461 1758 10495 1792
rect 10665 1758 10699 1792
rect 10461 1690 10495 1724
rect 10665 1690 10699 1724
rect 10461 1622 10495 1656
rect 10665 1622 10699 1656
rect 11023 2448 11057 2482
rect 11095 2448 11129 2482
rect 11023 2380 11057 2414
rect 11095 2380 11129 2414
rect 11023 2312 11057 2346
rect 11095 2312 11129 2346
rect 11023 2244 11057 2278
rect 11095 2244 11129 2278
rect 11023 2176 11057 2210
rect 11095 2176 11129 2210
rect 11023 2108 11057 2142
rect 11095 2108 11129 2142
rect 11023 2040 11057 2074
rect 11095 2040 11129 2074
rect 11023 1972 11057 2006
rect 11095 1972 11129 2006
rect 11023 1904 11057 1938
rect 11095 1904 11129 1938
rect 11023 1836 11057 1870
rect 11095 1836 11129 1870
rect 11023 1768 11057 1802
rect 11095 1768 11129 1802
rect 11023 1700 11057 1734
rect 11095 1700 11129 1734
rect 11023 1632 11057 1666
rect 11095 1632 11129 1666
rect 11023 1564 11057 1598
rect 11095 1564 11129 1598
rect 11453 2506 11487 2540
rect 11657 2506 11691 2540
rect 11453 2438 11487 2472
rect 11657 2438 11691 2472
rect 11453 2370 11487 2404
rect 11657 2370 11691 2404
rect 11453 2302 11487 2336
rect 11657 2302 11691 2336
rect 11453 2234 11487 2268
rect 11657 2234 11691 2268
rect 11453 2166 11487 2200
rect 11657 2166 11691 2200
rect 11453 2098 11487 2132
rect 11657 2098 11691 2132
rect 11453 2030 11487 2064
rect 11657 2030 11691 2064
rect 11453 1962 11487 1996
rect 11657 1962 11691 1996
rect 11453 1894 11487 1928
rect 11657 1894 11691 1928
rect 11453 1826 11487 1860
rect 11657 1826 11691 1860
rect 11453 1758 11487 1792
rect 11657 1758 11691 1792
rect 11453 1690 11487 1724
rect 11657 1690 11691 1724
rect 11453 1622 11487 1656
rect 11657 1622 11691 1656
rect 12015 2448 12049 2482
rect 12087 2448 12121 2482
rect 12015 2380 12049 2414
rect 12087 2380 12121 2414
rect 12015 2312 12049 2346
rect 12087 2312 12121 2346
rect 12015 2244 12049 2278
rect 12087 2244 12121 2278
rect 12015 2176 12049 2210
rect 12087 2176 12121 2210
rect 12015 2108 12049 2142
rect 12087 2108 12121 2142
rect 12015 2040 12049 2074
rect 12087 2040 12121 2074
rect 12015 1972 12049 2006
rect 12087 1972 12121 2006
rect 12015 1904 12049 1938
rect 12087 1904 12121 1938
rect 12015 1836 12049 1870
rect 12087 1836 12121 1870
rect 12015 1768 12049 1802
rect 12087 1768 12121 1802
rect 12015 1700 12049 1734
rect 12087 1700 12121 1734
rect 12015 1632 12049 1666
rect 12087 1632 12121 1666
rect 12015 1564 12049 1598
rect 12087 1564 12121 1598
rect 12445 2506 12479 2540
rect 12649 2506 12683 2540
rect 12445 2438 12479 2472
rect 12649 2438 12683 2472
rect 12445 2370 12479 2404
rect 12649 2370 12683 2404
rect 12445 2302 12479 2336
rect 12649 2302 12683 2336
rect 12445 2234 12479 2268
rect 12649 2234 12683 2268
rect 12445 2166 12479 2200
rect 12649 2166 12683 2200
rect 12445 2098 12479 2132
rect 12649 2098 12683 2132
rect 12445 2030 12479 2064
rect 12649 2030 12683 2064
rect 12445 1962 12479 1996
rect 12649 1962 12683 1996
rect 12445 1894 12479 1928
rect 12649 1894 12683 1928
rect 12445 1826 12479 1860
rect 12649 1826 12683 1860
rect 12445 1758 12479 1792
rect 12649 1758 12683 1792
rect 12445 1690 12479 1724
rect 12649 1690 12683 1724
rect 12445 1622 12479 1656
rect 12649 1622 12683 1656
rect 13007 2448 13041 2482
rect 13079 2448 13113 2482
rect 13007 2380 13041 2414
rect 13079 2380 13113 2414
rect 13007 2312 13041 2346
rect 13079 2312 13113 2346
rect 13007 2244 13041 2278
rect 13079 2244 13113 2278
rect 13007 2176 13041 2210
rect 13079 2176 13113 2210
rect 13007 2108 13041 2142
rect 13079 2108 13113 2142
rect 13007 2040 13041 2074
rect 13079 2040 13113 2074
rect 13007 1972 13041 2006
rect 13079 1972 13113 2006
rect 13007 1904 13041 1938
rect 13079 1904 13113 1938
rect 13007 1836 13041 1870
rect 13079 1836 13113 1870
rect 13007 1768 13041 1802
rect 13079 1768 13113 1802
rect 13007 1700 13041 1734
rect 13079 1700 13113 1734
rect 13007 1632 13041 1666
rect 13079 1632 13113 1666
rect 13007 1564 13041 1598
rect 13079 1564 13113 1598
rect 13437 2506 13471 2540
rect 13641 2506 13675 2540
rect 13437 2438 13471 2472
rect 13641 2438 13675 2472
rect 13437 2370 13471 2404
rect 13641 2370 13675 2404
rect 13437 2302 13471 2336
rect 13641 2302 13675 2336
rect 13437 2234 13471 2268
rect 13641 2234 13675 2268
rect 13437 2166 13471 2200
rect 13641 2166 13675 2200
rect 13437 2098 13471 2132
rect 13641 2098 13675 2132
rect 13437 2030 13471 2064
rect 13641 2030 13675 2064
rect 13437 1962 13471 1996
rect 13641 1962 13675 1996
rect 13437 1894 13471 1928
rect 13641 1894 13675 1928
rect 13437 1826 13471 1860
rect 13641 1826 13675 1860
rect 13437 1758 13471 1792
rect 13641 1758 13675 1792
rect 13437 1690 13471 1724
rect 13641 1690 13675 1724
rect 13437 1622 13471 1656
rect 13641 1622 13675 1656
rect 13999 2448 14033 2482
rect 13999 2380 14033 2414
rect 13999 2312 14033 2346
rect 13999 2244 14033 2278
rect 13999 2176 14033 2210
rect 13999 2108 14033 2142
rect 13999 2040 14033 2074
rect 13999 1972 14033 2006
rect 13999 1904 14033 1938
rect 13999 1836 14033 1870
rect 13999 1768 14033 1802
rect 13999 1700 14033 1734
rect 13999 1632 14033 1666
rect 13999 1564 14033 1598
rect 14356 2448 14390 2482
rect 14356 2380 14390 2414
rect 14356 2312 14390 2346
rect 14356 2244 14390 2278
rect 14356 2176 14390 2210
rect 14356 2108 14390 2142
rect 14356 2040 14390 2074
rect 14356 1972 14390 2006
rect 14356 1904 14390 1938
rect 14356 1836 14390 1870
rect 14356 1768 14390 1802
rect 14356 1700 14390 1734
rect 14356 1632 14390 1666
rect 14356 1564 14390 1598
<< mvpsubdiff >>
rect 159 5082 14940 5083
rect 159 5048 252 5082
rect 286 5048 320 5082
rect 354 5048 388 5082
rect 422 5048 456 5082
rect 490 5048 524 5082
rect 558 5048 592 5082
rect 626 5048 660 5082
rect 694 5048 728 5082
rect 762 5048 796 5082
rect 830 5048 864 5082
rect 898 5048 932 5082
rect 966 5048 1000 5082
rect 1034 5048 1068 5082
rect 1102 5048 1136 5082
rect 1170 5048 1204 5082
rect 1238 5048 1272 5082
rect 1306 5048 1340 5082
rect 1374 5048 1408 5082
rect 1442 5048 1476 5082
rect 1510 5048 1544 5082
rect 1578 5048 1612 5082
rect 1646 5048 1680 5082
rect 1714 5048 1748 5082
rect 1782 5048 1816 5082
rect 1850 5048 1884 5082
rect 1918 5048 1952 5082
rect 1986 5048 2020 5082
rect 2054 5048 2088 5082
rect 2122 5048 2156 5082
rect 2190 5048 2224 5082
rect 2258 5048 2292 5082
rect 2326 5048 2360 5082
rect 2394 5048 2428 5082
rect 2462 5048 2496 5082
rect 2530 5048 2564 5082
rect 2598 5048 2632 5082
rect 2666 5048 2700 5082
rect 2734 5048 2768 5082
rect 2802 5048 2836 5082
rect 2870 5048 2904 5082
rect 2938 5048 2972 5082
rect 3006 5048 3040 5082
rect 3074 5048 3108 5082
rect 3142 5048 3176 5082
rect 3210 5048 3244 5082
rect 3278 5048 3312 5082
rect 3346 5048 3380 5082
rect 3414 5048 3448 5082
rect 3482 5048 3516 5082
rect 3550 5048 3584 5082
rect 3618 5048 3652 5082
rect 3686 5048 3720 5082
rect 3754 5048 3788 5082
rect 3822 5048 3856 5082
rect 3890 5048 3924 5082
rect 3958 5048 3992 5082
rect 4026 5048 4060 5082
rect 4094 5048 4128 5082
rect 4162 5048 4196 5082
rect 4230 5048 4264 5082
rect 4298 5048 4332 5082
rect 4366 5048 4400 5082
rect 4434 5048 4468 5082
rect 4502 5048 4536 5082
rect 4570 5048 4604 5082
rect 4638 5048 4672 5082
rect 4706 5048 4740 5082
rect 4774 5048 4808 5082
rect 4842 5048 4876 5082
rect 4910 5048 4944 5082
rect 4978 5048 5012 5082
rect 5046 5048 5080 5082
rect 5114 5048 5148 5082
rect 5182 5048 5216 5082
rect 5250 5048 5284 5082
rect 5318 5048 5352 5082
rect 5386 5048 5420 5082
rect 5454 5048 5488 5082
rect 5522 5048 5556 5082
rect 5590 5048 5624 5082
rect 5658 5048 5692 5082
rect 5726 5048 5760 5082
rect 5794 5048 5828 5082
rect 5862 5048 5896 5082
rect 5930 5048 5964 5082
rect 5998 5048 6032 5082
rect 6066 5048 6100 5082
rect 6134 5048 6168 5082
rect 6202 5048 6236 5082
rect 6270 5048 6304 5082
rect 6338 5048 6372 5082
rect 6406 5048 6440 5082
rect 6474 5048 6508 5082
rect 6542 5048 6576 5082
rect 6610 5048 6644 5082
rect 6678 5048 6712 5082
rect 6746 5048 6780 5082
rect 6814 5048 6848 5082
rect 6882 5048 6916 5082
rect 6950 5048 6984 5082
rect 7018 5048 7052 5082
rect 7086 5048 7120 5082
rect 7154 5048 7188 5082
rect 7222 5048 7256 5082
rect 7290 5048 7324 5082
rect 7358 5048 7392 5082
rect 7426 5048 7460 5082
rect 7494 5048 7528 5082
rect 7562 5048 7596 5082
rect 7630 5048 7664 5082
rect 7698 5048 7732 5082
rect 7766 5048 7800 5082
rect 7834 5048 7868 5082
rect 7902 5048 7936 5082
rect 7970 5048 8004 5082
rect 8038 5048 8072 5082
rect 8106 5048 8140 5082
rect 8174 5048 8208 5082
rect 8242 5048 8276 5082
rect 8310 5048 8344 5082
rect 8378 5048 8412 5082
rect 8446 5048 8480 5082
rect 8514 5048 8548 5082
rect 8582 5048 8616 5082
rect 8650 5048 8684 5082
rect 8718 5048 8752 5082
rect 8786 5048 8820 5082
rect 8854 5048 8888 5082
rect 8922 5048 8956 5082
rect 8990 5048 9024 5082
rect 9058 5048 9092 5082
rect 9126 5048 9160 5082
rect 9194 5048 9228 5082
rect 9262 5048 9296 5082
rect 9330 5048 9364 5082
rect 9398 5048 9432 5082
rect 9466 5048 9500 5082
rect 9534 5048 9568 5082
rect 9602 5048 9636 5082
rect 9670 5048 9704 5082
rect 9738 5048 9772 5082
rect 9806 5048 9840 5082
rect 9874 5048 9908 5082
rect 9942 5048 9976 5082
rect 10010 5048 10044 5082
rect 10078 5048 10112 5082
rect 10146 5048 10180 5082
rect 10214 5048 10248 5082
rect 10282 5048 10316 5082
rect 10350 5048 10384 5082
rect 10418 5048 10452 5082
rect 10486 5048 10520 5082
rect 10554 5048 10588 5082
rect 10622 5048 10656 5082
rect 10690 5048 10724 5082
rect 10758 5048 10792 5082
rect 10826 5048 10860 5082
rect 10894 5048 10928 5082
rect 10962 5048 10996 5082
rect 11030 5048 11064 5082
rect 11098 5048 11132 5082
rect 11166 5048 11200 5082
rect 11234 5048 11268 5082
rect 11302 5048 11336 5082
rect 11370 5048 11404 5082
rect 11438 5048 11472 5082
rect 11506 5048 11540 5082
rect 11574 5048 11608 5082
rect 11642 5048 11676 5082
rect 11710 5048 11744 5082
rect 11778 5048 11812 5082
rect 11846 5048 11880 5082
rect 11914 5048 11948 5082
rect 11982 5048 12016 5082
rect 12050 5048 12084 5082
rect 12118 5048 12152 5082
rect 12186 5048 12220 5082
rect 12254 5048 12288 5082
rect 12322 5048 12356 5082
rect 12390 5048 12424 5082
rect 12458 5048 12492 5082
rect 12526 5048 12560 5082
rect 12594 5048 12628 5082
rect 12662 5048 12696 5082
rect 12730 5048 12764 5082
rect 12798 5048 12832 5082
rect 12866 5048 12900 5082
rect 12934 5048 12968 5082
rect 13002 5048 13036 5082
rect 13070 5048 13104 5082
rect 13138 5048 13172 5082
rect 13206 5048 13240 5082
rect 13274 5048 13308 5082
rect 13342 5048 13376 5082
rect 13410 5048 13444 5082
rect 13478 5048 13512 5082
rect 13546 5048 13580 5082
rect 13614 5048 13648 5082
rect 13682 5048 13716 5082
rect 13750 5048 13784 5082
rect 13818 5048 13852 5082
rect 13886 5048 13920 5082
rect 13954 5048 13988 5082
rect 14022 5048 14056 5082
rect 14090 5048 14124 5082
rect 14158 5048 14192 5082
rect 14226 5048 14260 5082
rect 14294 5048 14328 5082
rect 14362 5048 14396 5082
rect 14430 5048 14464 5082
rect 14498 5048 14532 5082
rect 14566 5048 14600 5082
rect 14634 5048 14668 5082
rect 14702 5048 14736 5082
rect 14770 5048 14804 5082
rect 14838 5048 14872 5082
rect 14906 5048 14940 5082
rect 159 5000 14940 5048
rect 159 4966 252 5000
rect 286 4966 320 5000
rect 354 4966 388 5000
rect 422 4966 456 5000
rect 490 4966 524 5000
rect 558 4966 592 5000
rect 626 4966 660 5000
rect 694 4966 728 5000
rect 762 4966 796 5000
rect 830 4966 864 5000
rect 898 4966 932 5000
rect 966 4966 1000 5000
rect 1034 4966 1068 5000
rect 1102 4966 1136 5000
rect 1170 4966 1204 5000
rect 1238 4966 1272 5000
rect 1306 4966 1340 5000
rect 1374 4966 1408 5000
rect 1442 4966 1476 5000
rect 1510 4966 1544 5000
rect 1578 4966 1612 5000
rect 1646 4966 1680 5000
rect 1714 4966 1748 5000
rect 1782 4966 1816 5000
rect 1850 4966 1884 5000
rect 1918 4966 1952 5000
rect 1986 4966 2020 5000
rect 2054 4966 2088 5000
rect 2122 4966 2156 5000
rect 2190 4966 2224 5000
rect 2258 4966 2292 5000
rect 2326 4966 2360 5000
rect 2394 4966 2428 5000
rect 2462 4966 2496 5000
rect 2530 4966 2564 5000
rect 2598 4966 2632 5000
rect 2666 4966 2700 5000
rect 2734 4966 2768 5000
rect 2802 4966 2836 5000
rect 2870 4966 2904 5000
rect 2938 4966 2972 5000
rect 3006 4966 3040 5000
rect 3074 4966 3108 5000
rect 3142 4966 3176 5000
rect 3210 4966 3244 5000
rect 3278 4966 3312 5000
rect 3346 4966 3380 5000
rect 3414 4966 3448 5000
rect 3482 4966 3516 5000
rect 3550 4966 3584 5000
rect 3618 4966 3652 5000
rect 3686 4966 3720 5000
rect 3754 4966 3788 5000
rect 3822 4966 3856 5000
rect 3890 4966 3924 5000
rect 3958 4966 3992 5000
rect 4026 4966 4060 5000
rect 4094 4966 4128 5000
rect 4162 4966 4196 5000
rect 4230 4966 4264 5000
rect 4298 4966 4332 5000
rect 4366 4966 4400 5000
rect 4434 4966 4468 5000
rect 4502 4966 4536 5000
rect 4570 4966 4604 5000
rect 4638 4966 4672 5000
rect 4706 4966 4740 5000
rect 4774 4966 4808 5000
rect 4842 4966 4876 5000
rect 4910 4966 4944 5000
rect 4978 4966 5012 5000
rect 5046 4966 5080 5000
rect 5114 4966 5148 5000
rect 5182 4966 5216 5000
rect 5250 4966 5284 5000
rect 5318 4966 5352 5000
rect 5386 4966 5420 5000
rect 5454 4966 5488 5000
rect 5522 4966 5556 5000
rect 5590 4966 5624 5000
rect 5658 4966 5692 5000
rect 5726 4966 5760 5000
rect 5794 4966 5828 5000
rect 5862 4966 5896 5000
rect 5930 4966 5964 5000
rect 5998 4966 6032 5000
rect 6066 4966 6100 5000
rect 6134 4966 6168 5000
rect 6202 4966 6236 5000
rect 6270 4966 6304 5000
rect 6338 4966 6372 5000
rect 6406 4966 6440 5000
rect 6474 4966 6508 5000
rect 6542 4966 6576 5000
rect 6610 4966 6644 5000
rect 6678 4966 6712 5000
rect 6746 4966 6780 5000
rect 6814 4966 6848 5000
rect 6882 4966 6916 5000
rect 6950 4966 6984 5000
rect 7018 4966 7052 5000
rect 7086 4966 7120 5000
rect 7154 4966 7188 5000
rect 7222 4966 7256 5000
rect 7290 4966 7324 5000
rect 7358 4966 7392 5000
rect 7426 4966 7460 5000
rect 7494 4966 7528 5000
rect 7562 4966 7596 5000
rect 7630 4966 7664 5000
rect 7698 4966 7732 5000
rect 7766 4966 7800 5000
rect 7834 4966 7868 5000
rect 7902 4966 7936 5000
rect 7970 4966 8004 5000
rect 8038 4966 8072 5000
rect 8106 4966 8140 5000
rect 8174 4966 8208 5000
rect 8242 4966 8276 5000
rect 8310 4966 8344 5000
rect 8378 4966 8412 5000
rect 8446 4966 8480 5000
rect 8514 4966 8548 5000
rect 8582 4966 8616 5000
rect 8650 4966 8684 5000
rect 8718 4966 8752 5000
rect 8786 4966 8820 5000
rect 8854 4966 8888 5000
rect 8922 4966 8956 5000
rect 8990 4966 9024 5000
rect 9058 4966 9092 5000
rect 9126 4966 9160 5000
rect 9194 4966 9228 5000
rect 9262 4966 9296 5000
rect 9330 4966 9364 5000
rect 9398 4966 9432 5000
rect 9466 4966 9500 5000
rect 9534 4966 9568 5000
rect 9602 4966 9636 5000
rect 9670 4966 9704 5000
rect 9738 4966 9772 5000
rect 9806 4966 9840 5000
rect 9874 4966 9908 5000
rect 9942 4966 9976 5000
rect 10010 4966 10044 5000
rect 10078 4966 10112 5000
rect 10146 4966 10180 5000
rect 10214 4966 10248 5000
rect 10282 4966 10316 5000
rect 10350 4966 10384 5000
rect 10418 4966 10452 5000
rect 10486 4966 10520 5000
rect 10554 4966 10588 5000
rect 10622 4966 10656 5000
rect 10690 4966 10724 5000
rect 10758 4966 10792 5000
rect 10826 4966 10860 5000
rect 10894 4966 10928 5000
rect 10962 4966 10996 5000
rect 11030 4966 11064 5000
rect 11098 4966 11132 5000
rect 11166 4966 11200 5000
rect 11234 4966 11268 5000
rect 11302 4966 11336 5000
rect 11370 4966 11404 5000
rect 11438 4966 11472 5000
rect 11506 4966 11540 5000
rect 11574 4966 11608 5000
rect 11642 4966 11676 5000
rect 11710 4966 11744 5000
rect 11778 4966 11812 5000
rect 11846 4966 11880 5000
rect 11914 4966 11948 5000
rect 11982 4966 12016 5000
rect 12050 4966 12084 5000
rect 12118 4966 12152 5000
rect 12186 4966 12220 5000
rect 12254 4966 12288 5000
rect 12322 4966 12356 5000
rect 12390 4966 12424 5000
rect 12458 4966 12492 5000
rect 12526 4966 12560 5000
rect 12594 4966 12628 5000
rect 12662 4966 12696 5000
rect 12730 4966 12764 5000
rect 12798 4966 12832 5000
rect 12866 4966 12900 5000
rect 12934 4966 12968 5000
rect 13002 4966 13036 5000
rect 13070 4966 13104 5000
rect 13138 4966 13172 5000
rect 13206 4966 13240 5000
rect 13274 4966 13308 5000
rect 13342 4966 13376 5000
rect 13410 4966 13444 5000
rect 13478 4966 13512 5000
rect 13546 4966 13580 5000
rect 13614 4966 13648 5000
rect 13682 4966 13716 5000
rect 13750 4966 13784 5000
rect 13818 4966 13852 5000
rect 13886 4966 13920 5000
rect 13954 4966 13988 5000
rect 14022 4966 14056 5000
rect 14090 4966 14124 5000
rect 14158 4966 14192 5000
rect 14226 4966 14260 5000
rect 14294 4966 14328 5000
rect 14362 4966 14396 5000
rect 14430 4966 14464 5000
rect 14498 4966 14532 5000
rect 14566 4966 14600 5000
rect 14634 4966 14668 5000
rect 14702 4966 14736 5000
rect 14770 4966 14804 5000
rect 14838 4966 14872 5000
rect 14906 4966 14940 5000
rect 159 4918 14940 4966
rect 159 4884 252 4918
rect 286 4884 320 4918
rect 354 4884 388 4918
rect 422 4884 456 4918
rect 490 4884 524 4918
rect 558 4884 592 4918
rect 626 4884 660 4918
rect 694 4884 728 4918
rect 762 4884 796 4918
rect 830 4884 864 4918
rect 898 4884 932 4918
rect 966 4884 1000 4918
rect 1034 4884 1068 4918
rect 1102 4884 1136 4918
rect 1170 4884 1204 4918
rect 1238 4884 1272 4918
rect 1306 4884 1340 4918
rect 1374 4884 1408 4918
rect 1442 4884 1476 4918
rect 1510 4884 1544 4918
rect 1578 4884 1612 4918
rect 1646 4884 1680 4918
rect 1714 4884 1748 4918
rect 1782 4884 1816 4918
rect 1850 4884 1884 4918
rect 1918 4884 1952 4918
rect 1986 4884 2020 4918
rect 2054 4884 2088 4918
rect 2122 4884 2156 4918
rect 2190 4884 2224 4918
rect 2258 4884 2292 4918
rect 2326 4884 2360 4918
rect 2394 4884 2428 4918
rect 2462 4884 2496 4918
rect 2530 4884 2564 4918
rect 2598 4884 2632 4918
rect 2666 4884 2700 4918
rect 2734 4884 2768 4918
rect 2802 4884 2836 4918
rect 2870 4884 2904 4918
rect 2938 4884 2972 4918
rect 3006 4884 3040 4918
rect 3074 4884 3108 4918
rect 3142 4884 3176 4918
rect 3210 4884 3244 4918
rect 3278 4884 3312 4918
rect 3346 4884 3380 4918
rect 3414 4884 3448 4918
rect 3482 4884 3516 4918
rect 3550 4884 3584 4918
rect 3618 4884 3652 4918
rect 3686 4884 3720 4918
rect 3754 4884 3788 4918
rect 3822 4884 3856 4918
rect 3890 4884 3924 4918
rect 3958 4884 3992 4918
rect 4026 4884 4060 4918
rect 4094 4884 4128 4918
rect 4162 4884 4196 4918
rect 4230 4884 4264 4918
rect 4298 4884 4332 4918
rect 4366 4884 4400 4918
rect 4434 4884 4468 4918
rect 4502 4884 4536 4918
rect 4570 4884 4604 4918
rect 4638 4884 4672 4918
rect 4706 4884 4740 4918
rect 4774 4884 4808 4918
rect 4842 4884 4876 4918
rect 4910 4884 4944 4918
rect 4978 4884 5012 4918
rect 5046 4884 5080 4918
rect 5114 4884 5148 4918
rect 5182 4884 5216 4918
rect 5250 4884 5284 4918
rect 5318 4884 5352 4918
rect 5386 4884 5420 4918
rect 5454 4884 5488 4918
rect 5522 4884 5556 4918
rect 5590 4884 5624 4918
rect 5658 4884 5692 4918
rect 5726 4884 5760 4918
rect 5794 4884 5828 4918
rect 5862 4884 5896 4918
rect 5930 4884 5964 4918
rect 5998 4884 6032 4918
rect 6066 4884 6100 4918
rect 6134 4884 6168 4918
rect 6202 4884 6236 4918
rect 6270 4884 6304 4918
rect 6338 4884 6372 4918
rect 6406 4884 6440 4918
rect 6474 4884 6508 4918
rect 6542 4884 6576 4918
rect 6610 4884 6644 4918
rect 6678 4884 6712 4918
rect 6746 4884 6780 4918
rect 6814 4884 6848 4918
rect 6882 4884 6916 4918
rect 6950 4884 6984 4918
rect 7018 4884 7052 4918
rect 7086 4884 7120 4918
rect 7154 4884 7188 4918
rect 7222 4884 7256 4918
rect 7290 4884 7324 4918
rect 7358 4884 7392 4918
rect 7426 4884 7460 4918
rect 7494 4884 7528 4918
rect 7562 4884 7596 4918
rect 7630 4884 7664 4918
rect 7698 4884 7732 4918
rect 7766 4884 7800 4918
rect 7834 4884 7868 4918
rect 7902 4884 7936 4918
rect 7970 4884 8004 4918
rect 8038 4884 8072 4918
rect 8106 4884 8140 4918
rect 8174 4884 8208 4918
rect 8242 4884 8276 4918
rect 8310 4884 8344 4918
rect 8378 4884 8412 4918
rect 8446 4884 8480 4918
rect 8514 4884 8548 4918
rect 8582 4884 8616 4918
rect 8650 4884 8684 4918
rect 8718 4884 8752 4918
rect 8786 4884 8820 4918
rect 8854 4884 8888 4918
rect 8922 4884 8956 4918
rect 8990 4884 9024 4918
rect 9058 4884 9092 4918
rect 9126 4884 9160 4918
rect 9194 4884 9228 4918
rect 9262 4884 9296 4918
rect 9330 4884 9364 4918
rect 9398 4884 9432 4918
rect 9466 4884 9500 4918
rect 9534 4884 9568 4918
rect 9602 4884 9636 4918
rect 9670 4884 9704 4918
rect 9738 4884 9772 4918
rect 9806 4884 9840 4918
rect 9874 4884 9908 4918
rect 9942 4884 9976 4918
rect 10010 4884 10044 4918
rect 10078 4884 10112 4918
rect 10146 4884 10180 4918
rect 10214 4884 10248 4918
rect 10282 4884 10316 4918
rect 10350 4884 10384 4918
rect 10418 4884 10452 4918
rect 10486 4884 10520 4918
rect 10554 4884 10588 4918
rect 10622 4884 10656 4918
rect 10690 4884 10724 4918
rect 10758 4884 10792 4918
rect 10826 4884 10860 4918
rect 10894 4884 10928 4918
rect 10962 4884 10996 4918
rect 11030 4884 11064 4918
rect 11098 4884 11132 4918
rect 11166 4884 11200 4918
rect 11234 4884 11268 4918
rect 11302 4884 11336 4918
rect 11370 4884 11404 4918
rect 11438 4884 11472 4918
rect 11506 4884 11540 4918
rect 11574 4884 11608 4918
rect 11642 4884 11676 4918
rect 11710 4884 11744 4918
rect 11778 4884 11812 4918
rect 11846 4884 11880 4918
rect 11914 4884 11948 4918
rect 11982 4884 12016 4918
rect 12050 4884 12084 4918
rect 12118 4884 12152 4918
rect 12186 4884 12220 4918
rect 12254 4884 12288 4918
rect 12322 4884 12356 4918
rect 12390 4884 12424 4918
rect 12458 4884 12492 4918
rect 12526 4884 12560 4918
rect 12594 4884 12628 4918
rect 12662 4884 12696 4918
rect 12730 4884 12764 4918
rect 12798 4884 12832 4918
rect 12866 4884 12900 4918
rect 12934 4884 12968 4918
rect 13002 4884 13036 4918
rect 13070 4884 13104 4918
rect 13138 4884 13172 4918
rect 13206 4884 13240 4918
rect 13274 4884 13308 4918
rect 13342 4884 13376 4918
rect 13410 4884 13444 4918
rect 13478 4884 13512 4918
rect 13546 4884 13580 4918
rect 13614 4884 13648 4918
rect 13682 4884 13716 4918
rect 13750 4884 13784 4918
rect 13818 4884 13852 4918
rect 13886 4884 13920 4918
rect 13954 4884 13988 4918
rect 14022 4884 14056 4918
rect 14090 4884 14124 4918
rect 14158 4884 14192 4918
rect 14226 4884 14260 4918
rect 14294 4884 14328 4918
rect 14362 4884 14396 4918
rect 14430 4884 14464 4918
rect 14498 4884 14532 4918
rect 14566 4884 14600 4918
rect 14634 4884 14668 4918
rect 14702 4884 14736 4918
rect 14770 4884 14804 4918
rect 14838 4884 14872 4918
rect 14906 4884 14940 4918
rect 159 4883 14940 4884
rect 159 4849 329 4883
rect 159 599 193 4849
rect 295 599 329 4849
rect 14806 4849 14940 4883
rect 14840 4815 14906 4849
rect 14806 4781 14940 4815
rect 14840 4747 14906 4781
rect 14806 4713 14940 4747
rect 14840 4679 14906 4713
rect 14806 4645 14940 4679
rect 14840 4611 14906 4645
rect 14806 4577 14940 4611
rect 14840 4543 14906 4577
rect 14806 4509 14940 4543
rect 14840 4475 14906 4509
rect 14806 4441 14940 4475
rect 14840 4407 14906 4441
rect 14806 4373 14940 4407
rect 14840 4339 14906 4373
rect 14806 4305 14940 4339
rect 14840 4271 14906 4305
rect 14806 4237 14940 4271
rect 14840 4203 14906 4237
rect 14806 4169 14940 4203
rect 14840 4135 14906 4169
rect 14806 4101 14940 4135
rect 14840 4067 14906 4101
rect 14806 4033 14940 4067
rect 14840 3999 14906 4033
rect 14806 3965 14940 3999
rect 14840 3931 14906 3965
rect 14806 3897 14940 3931
rect 14840 3863 14906 3897
rect 14806 3829 14940 3863
rect 14840 3795 14906 3829
rect 14806 3761 14940 3795
rect 14840 3727 14906 3761
rect 14806 3693 14940 3727
rect 14840 3659 14906 3693
rect 14806 3625 14940 3659
rect 14840 3591 14906 3625
rect 14806 3557 14940 3591
rect 14840 3523 14906 3557
rect 14806 3489 14940 3523
rect 14840 3455 14906 3489
rect 14806 3421 14940 3455
rect 14840 3387 14906 3421
rect 14806 3353 14940 3387
rect 14840 3319 14906 3353
rect 14806 3285 14940 3319
rect 14840 3251 14906 3285
rect 14806 3217 14940 3251
rect 14840 3183 14906 3217
rect 14806 3149 14940 3183
rect 14840 3115 14906 3149
rect 14806 3081 14940 3115
rect 14840 3047 14906 3081
rect 14806 3013 14940 3047
rect 14840 2979 14906 3013
rect 14806 2945 14940 2979
rect 14840 2911 14906 2945
rect 14806 2877 14940 2911
rect 14840 2843 14906 2877
rect 14806 2809 14940 2843
rect 14840 2775 14906 2809
rect 14806 2741 14940 2775
rect 14840 2707 14906 2741
rect 14806 2673 14940 2707
rect 14840 2639 14906 2673
rect 14806 2605 14940 2639
rect 14840 2571 14906 2605
rect 14806 2537 14940 2571
rect 14840 2503 14906 2537
rect 14806 2469 14940 2503
rect 14840 2435 14906 2469
rect 14806 2401 14940 2435
rect 14840 2367 14906 2401
rect 14806 2333 14940 2367
rect 14840 2299 14906 2333
rect 14806 2265 14940 2299
rect 14840 2231 14906 2265
rect 14806 2197 14940 2231
rect 14840 2163 14906 2197
rect 14806 2129 14940 2163
rect 14840 2095 14906 2129
rect 14806 2061 14940 2095
rect 14840 2027 14906 2061
rect 14806 1993 14940 2027
rect 14840 1959 14906 1993
rect 14806 1925 14940 1959
rect 14840 1891 14906 1925
rect 14806 1857 14940 1891
rect 14840 1823 14906 1857
rect 14806 1789 14940 1823
rect 14840 1755 14906 1789
rect 14806 1721 14940 1755
rect 14840 1687 14906 1721
rect 14806 1653 14940 1687
rect 14840 1619 14906 1653
rect 14806 1585 14940 1619
rect 14840 1551 14906 1585
rect 14806 1517 14940 1551
rect 14840 1483 14906 1517
rect 14806 1449 14940 1483
rect 14840 1415 14906 1449
rect 14806 1381 14940 1415
rect 14840 1347 14906 1381
rect 14806 1313 14940 1347
rect 14840 1279 14906 1313
rect 14806 1245 14940 1279
rect 14840 1211 14906 1245
rect 14806 1177 14940 1211
rect 14840 1143 14906 1177
rect 14806 1109 14940 1143
rect 14840 1075 14906 1109
rect 14806 1041 14940 1075
rect 14840 1007 14906 1041
rect 14806 973 14940 1007
rect 14840 939 14906 973
rect 14806 905 14940 939
rect 14840 871 14906 905
rect 14806 837 14940 871
rect 14840 803 14906 837
rect 14806 769 14940 803
rect 14840 735 14906 769
rect 14806 701 14940 735
rect 14840 667 14906 701
rect 159 509 329 599
rect 14806 633 14940 667
rect 14840 599 14906 633
rect 14806 509 14940 599
rect 159 407 193 509
rect 14847 407 14940 509
rect 159 309 14940 407
<< mvnsubdiff >>
rect 482 4638 14653 4653
rect 482 4619 584 4638
rect 482 4585 497 4619
rect 531 4585 584 4619
rect 482 4570 584 4585
rect 10410 4604 10445 4638
rect 10479 4604 10514 4638
rect 10548 4604 10583 4638
rect 10617 4604 10652 4638
rect 10686 4604 10721 4638
rect 10755 4604 10790 4638
rect 10824 4604 10859 4638
rect 10893 4604 10928 4638
rect 10962 4604 10997 4638
rect 11031 4604 11066 4638
rect 11100 4604 11135 4638
rect 11169 4604 11204 4638
rect 11238 4604 11273 4638
rect 11307 4604 11342 4638
rect 11376 4604 11411 4638
rect 11445 4604 11480 4638
rect 11514 4604 11549 4638
rect 11583 4604 11618 4638
rect 11652 4604 11687 4638
rect 11721 4604 11756 4638
rect 11790 4604 11825 4638
rect 11859 4604 11894 4638
rect 11928 4604 11963 4638
rect 11997 4604 12032 4638
rect 12066 4604 12101 4638
rect 12135 4604 12170 4638
rect 12204 4604 12239 4638
rect 12273 4604 12308 4638
rect 12342 4604 12377 4638
rect 12411 4604 12446 4638
rect 12480 4604 12515 4638
rect 12549 4604 12584 4638
rect 12618 4604 12653 4638
rect 12687 4604 12722 4638
rect 12756 4604 12791 4638
rect 12825 4604 12860 4638
rect 12894 4604 12929 4638
rect 12963 4604 12998 4638
rect 13032 4604 13067 4638
rect 13101 4604 13136 4638
rect 13170 4604 13205 4638
rect 13239 4604 13274 4638
rect 13308 4604 13343 4638
rect 13377 4604 13412 4638
rect 13446 4604 13481 4638
rect 13515 4604 13550 4638
rect 13584 4604 13619 4638
rect 13653 4604 13688 4638
rect 13722 4604 13757 4638
rect 13791 4604 13826 4638
rect 13860 4604 13895 4638
rect 13929 4604 13964 4638
rect 13998 4604 14033 4638
rect 14067 4604 14102 4638
rect 14136 4604 14171 4638
rect 14205 4604 14240 4638
rect 14274 4604 14309 4638
rect 14343 4604 14378 4638
rect 14412 4604 14447 4638
rect 14481 4604 14516 4638
rect 14550 4604 14585 4638
rect 14619 4604 14653 4638
rect 10410 4570 14653 4604
rect 482 4549 565 4570
rect 482 4515 497 4549
rect 531 4536 565 4549
rect 12363 4536 12397 4570
rect 12431 4536 12466 4570
rect 12500 4536 12535 4570
rect 12569 4536 12604 4570
rect 12638 4536 12673 4570
rect 12707 4536 12742 4570
rect 12776 4536 12811 4570
rect 12845 4536 12880 4570
rect 12914 4536 12949 4570
rect 12983 4536 13018 4570
rect 13052 4536 13087 4570
rect 13121 4536 13156 4570
rect 13190 4536 13225 4570
rect 13259 4536 13294 4570
rect 13328 4536 13363 4570
rect 13397 4536 13432 4570
rect 13466 4536 13501 4570
rect 13535 4536 13570 4570
rect 13604 4536 13639 4570
rect 13673 4536 13708 4570
rect 13742 4536 13777 4570
rect 13811 4536 13846 4570
rect 13880 4536 13915 4570
rect 13949 4536 13984 4570
rect 14018 4536 14053 4570
rect 14087 4536 14122 4570
rect 14156 4536 14191 4570
rect 14225 4536 14260 4570
rect 14294 4536 14329 4570
rect 14363 4536 14398 4570
rect 14432 4536 14467 4570
rect 14501 4536 14536 4570
rect 14570 4551 14653 4570
rect 531 4515 633 4536
rect 482 4498 633 4515
rect 482 4479 565 4498
rect 482 4445 497 4479
rect 531 4464 565 4479
rect 599 4468 633 4498
rect 12363 4502 14536 4536
rect 12363 4468 12398 4502
rect 12432 4468 12467 4502
rect 12501 4468 12536 4502
rect 12570 4468 12605 4502
rect 12639 4468 12674 4502
rect 12708 4468 12743 4502
rect 12777 4468 12812 4502
rect 12846 4468 12881 4502
rect 12915 4468 12950 4502
rect 12984 4468 13019 4502
rect 13053 4468 13088 4502
rect 13122 4468 13157 4502
rect 13191 4468 13226 4502
rect 13260 4468 13295 4502
rect 13329 4468 13364 4502
rect 13398 4468 13433 4502
rect 13467 4468 13502 4502
rect 13536 4468 13571 4502
rect 13605 4468 13640 4502
rect 13674 4468 13709 4502
rect 13743 4468 13778 4502
rect 13812 4468 13847 4502
rect 13881 4468 13916 4502
rect 13950 4468 13985 4502
rect 14019 4468 14054 4502
rect 14088 4468 14123 4502
rect 14157 4468 14192 4502
rect 14226 4468 14261 4502
rect 14295 4468 14330 4502
rect 14364 4468 14399 4502
rect 14433 4468 14468 4502
rect 599 4464 14468 4468
rect 531 4453 14468 4464
rect 531 4445 682 4453
rect 482 4429 682 4445
rect 482 4426 633 4429
rect 482 4409 565 4426
rect 482 4375 497 4409
rect 531 4392 565 4409
rect 599 4395 633 4426
rect 667 4395 682 4429
rect 599 4392 682 4395
rect 531 4375 682 4392
rect 482 4356 682 4375
rect 482 4354 633 4356
rect 482 4339 565 4354
rect 482 4305 497 4339
rect 531 4320 565 4339
rect 599 4322 633 4354
rect 667 4322 682 4356
rect 599 4320 682 4322
rect 531 4305 682 4320
rect 482 4283 682 4305
rect 482 4282 633 4283
rect 482 4269 565 4282
rect 482 4235 497 4269
rect 531 4248 565 4269
rect 599 4249 633 4282
rect 667 4249 682 4283
rect 599 4248 682 4249
rect 531 4235 682 4248
rect 482 4211 682 4235
rect 482 4210 633 4211
rect 482 4199 565 4210
rect 482 4165 497 4199
rect 531 4176 565 4199
rect 599 4177 633 4210
rect 667 4177 682 4211
rect 599 4176 682 4177
rect 531 4165 682 4176
rect 482 4152 682 4165
rect 14453 4152 14468 4453
rect 482 4139 708 4152
rect 482 4138 633 4139
rect 482 4129 565 4138
rect 482 4095 497 4129
rect 531 4104 565 4129
rect 599 4105 633 4138
rect 667 4105 708 4139
rect 599 4104 708 4105
rect 531 4095 708 4104
rect 482 4067 708 4095
rect 482 4066 633 4067
rect 482 4059 565 4066
rect 482 4025 497 4059
rect 531 4032 565 4059
rect 599 4033 633 4066
rect 667 4033 708 4067
rect 599 4032 708 4033
rect 531 4025 708 4032
rect 482 3995 708 4025
rect 482 3994 633 3995
rect 482 3989 565 3994
rect 482 3955 497 3989
rect 531 3960 565 3989
rect 599 3961 633 3994
rect 667 3961 708 3995
rect 599 3960 708 3961
rect 531 3955 708 3960
rect 482 3923 708 3955
rect 482 3922 633 3923
rect 482 3920 565 3922
rect 482 3886 497 3920
rect 531 3888 565 3920
rect 599 3889 633 3922
rect 667 3889 708 3923
rect 599 3888 708 3889
rect 531 3886 708 3888
rect 482 3851 708 3886
rect 482 3817 497 3851
rect 531 3817 565 3851
rect 599 3817 633 3851
rect 667 3817 708 3851
rect 482 3749 708 3817
rect 482 3715 497 3749
rect 531 3715 565 3749
rect 599 3715 633 3749
rect 667 3715 708 3749
rect 482 3680 708 3715
rect 482 3646 497 3680
rect 531 3646 565 3680
rect 599 3646 633 3680
rect 667 3646 708 3680
rect 482 3611 708 3646
rect 482 3577 497 3611
rect 531 3577 565 3611
rect 599 3577 633 3611
rect 667 3577 708 3611
rect 482 3542 708 3577
rect 482 3508 497 3542
rect 531 3508 565 3542
rect 599 3508 633 3542
rect 667 3508 708 3542
rect 482 3473 708 3508
rect 482 3439 497 3473
rect 531 3439 565 3473
rect 599 3439 633 3473
rect 667 3439 708 3473
rect 482 3404 708 3439
rect 482 3370 497 3404
rect 531 3370 565 3404
rect 599 3370 633 3404
rect 667 3370 708 3404
rect 482 3335 708 3370
rect 482 3301 497 3335
rect 531 3301 565 3335
rect 599 3301 633 3335
rect 667 3301 708 3335
rect 482 3266 708 3301
rect 482 3232 497 3266
rect 531 3232 565 3266
rect 599 3232 633 3266
rect 667 3232 708 3266
rect 482 3197 708 3232
rect 482 3163 497 3197
rect 531 3163 565 3197
rect 599 3163 633 3197
rect 667 3163 708 3197
rect 482 3152 708 3163
rect 1582 4082 1722 4152
rect 1582 4048 1635 4082
rect 1669 4048 1722 4082
rect 1582 4014 1722 4048
rect 1582 3980 1635 4014
rect 1669 3980 1722 4014
rect 1582 3946 1722 3980
rect 1582 3912 1635 3946
rect 1669 3912 1722 3946
rect 1582 3878 1722 3912
rect 1582 3844 1635 3878
rect 1669 3844 1722 3878
rect 1582 3810 1722 3844
rect 1582 3776 1635 3810
rect 1669 3776 1722 3810
rect 1582 3742 1722 3776
rect 1582 3708 1635 3742
rect 1669 3708 1722 3742
rect 1582 3674 1722 3708
rect 1582 3640 1635 3674
rect 1669 3640 1722 3674
rect 1582 3606 1722 3640
rect 1582 3572 1635 3606
rect 1669 3572 1722 3606
rect 1582 3538 1722 3572
rect 1582 3504 1635 3538
rect 1669 3504 1722 3538
rect 1582 3470 1722 3504
rect 1582 3436 1635 3470
rect 1669 3436 1722 3470
rect 1582 3402 1722 3436
rect 1582 3368 1635 3402
rect 1669 3368 1722 3402
rect 1582 3334 1722 3368
rect 1582 3300 1635 3334
rect 1669 3300 1722 3334
rect 1582 3266 1722 3300
rect 1582 3232 1635 3266
rect 1669 3232 1722 3266
rect 1582 3198 1722 3232
rect 1582 3164 1635 3198
rect 1669 3164 1722 3198
rect 1582 3152 1722 3164
rect 2574 4082 2714 4152
rect 2574 4048 2627 4082
rect 2661 4048 2714 4082
rect 2574 4014 2714 4048
rect 2574 3980 2627 4014
rect 2661 3980 2714 4014
rect 2574 3946 2714 3980
rect 2574 3912 2627 3946
rect 2661 3912 2714 3946
rect 2574 3878 2714 3912
rect 2574 3844 2627 3878
rect 2661 3844 2714 3878
rect 2574 3810 2714 3844
rect 2574 3776 2627 3810
rect 2661 3776 2714 3810
rect 2574 3742 2714 3776
rect 2574 3708 2627 3742
rect 2661 3708 2714 3742
rect 2574 3674 2714 3708
rect 2574 3640 2627 3674
rect 2661 3640 2714 3674
rect 2574 3606 2714 3640
rect 2574 3572 2627 3606
rect 2661 3572 2714 3606
rect 2574 3538 2714 3572
rect 2574 3504 2627 3538
rect 2661 3504 2714 3538
rect 2574 3470 2714 3504
rect 2574 3436 2627 3470
rect 2661 3436 2714 3470
rect 2574 3402 2714 3436
rect 2574 3368 2627 3402
rect 2661 3368 2714 3402
rect 2574 3334 2714 3368
rect 2574 3300 2627 3334
rect 2661 3300 2714 3334
rect 2574 3266 2714 3300
rect 2574 3232 2627 3266
rect 2661 3232 2714 3266
rect 2574 3198 2714 3232
rect 2574 3164 2627 3198
rect 2661 3164 2714 3198
rect 2574 3152 2714 3164
rect 3566 4082 3706 4152
rect 3566 4048 3619 4082
rect 3653 4048 3706 4082
rect 3566 4014 3706 4048
rect 3566 3980 3619 4014
rect 3653 3980 3706 4014
rect 3566 3946 3706 3980
rect 3566 3912 3619 3946
rect 3653 3912 3706 3946
rect 3566 3878 3706 3912
rect 3566 3844 3619 3878
rect 3653 3844 3706 3878
rect 3566 3810 3706 3844
rect 3566 3776 3619 3810
rect 3653 3776 3706 3810
rect 3566 3742 3706 3776
rect 3566 3708 3619 3742
rect 3653 3708 3706 3742
rect 3566 3674 3706 3708
rect 3566 3640 3619 3674
rect 3653 3640 3706 3674
rect 3566 3606 3706 3640
rect 3566 3572 3619 3606
rect 3653 3572 3706 3606
rect 3566 3538 3706 3572
rect 3566 3504 3619 3538
rect 3653 3504 3706 3538
rect 3566 3470 3706 3504
rect 3566 3436 3619 3470
rect 3653 3436 3706 3470
rect 3566 3402 3706 3436
rect 3566 3368 3619 3402
rect 3653 3368 3706 3402
rect 3566 3334 3706 3368
rect 3566 3300 3619 3334
rect 3653 3300 3706 3334
rect 3566 3266 3706 3300
rect 3566 3232 3619 3266
rect 3653 3232 3706 3266
rect 3566 3198 3706 3232
rect 3566 3164 3619 3198
rect 3653 3164 3706 3198
rect 3566 3152 3706 3164
rect 4558 4082 4698 4152
rect 4558 4048 4611 4082
rect 4645 4048 4698 4082
rect 4558 4014 4698 4048
rect 4558 3980 4611 4014
rect 4645 3980 4698 4014
rect 4558 3946 4698 3980
rect 4558 3912 4611 3946
rect 4645 3912 4698 3946
rect 4558 3878 4698 3912
rect 4558 3844 4611 3878
rect 4645 3844 4698 3878
rect 4558 3810 4698 3844
rect 4558 3776 4611 3810
rect 4645 3776 4698 3810
rect 4558 3742 4698 3776
rect 4558 3708 4611 3742
rect 4645 3708 4698 3742
rect 4558 3674 4698 3708
rect 4558 3640 4611 3674
rect 4645 3640 4698 3674
rect 4558 3606 4698 3640
rect 4558 3572 4611 3606
rect 4645 3572 4698 3606
rect 4558 3538 4698 3572
rect 4558 3504 4611 3538
rect 4645 3504 4698 3538
rect 4558 3470 4698 3504
rect 4558 3436 4611 3470
rect 4645 3436 4698 3470
rect 4558 3402 4698 3436
rect 4558 3368 4611 3402
rect 4645 3368 4698 3402
rect 4558 3334 4698 3368
rect 4558 3300 4611 3334
rect 4645 3300 4698 3334
rect 4558 3266 4698 3300
rect 4558 3232 4611 3266
rect 4645 3232 4698 3266
rect 4558 3198 4698 3232
rect 4558 3164 4611 3198
rect 4645 3164 4698 3198
rect 4558 3152 4698 3164
rect 5550 4082 5690 4152
rect 5550 4048 5603 4082
rect 5637 4048 5690 4082
rect 5550 4014 5690 4048
rect 5550 3980 5603 4014
rect 5637 3980 5690 4014
rect 5550 3946 5690 3980
rect 5550 3912 5603 3946
rect 5637 3912 5690 3946
rect 5550 3878 5690 3912
rect 5550 3844 5603 3878
rect 5637 3844 5690 3878
rect 5550 3810 5690 3844
rect 5550 3776 5603 3810
rect 5637 3776 5690 3810
rect 5550 3742 5690 3776
rect 5550 3708 5603 3742
rect 5637 3708 5690 3742
rect 5550 3674 5690 3708
rect 5550 3640 5603 3674
rect 5637 3640 5690 3674
rect 5550 3606 5690 3640
rect 5550 3572 5603 3606
rect 5637 3572 5690 3606
rect 5550 3538 5690 3572
rect 5550 3504 5603 3538
rect 5637 3504 5690 3538
rect 5550 3470 5690 3504
rect 5550 3436 5603 3470
rect 5637 3436 5690 3470
rect 5550 3402 5690 3436
rect 5550 3368 5603 3402
rect 5637 3368 5690 3402
rect 5550 3334 5690 3368
rect 5550 3300 5603 3334
rect 5637 3300 5690 3334
rect 5550 3266 5690 3300
rect 5550 3232 5603 3266
rect 5637 3232 5690 3266
rect 5550 3198 5690 3232
rect 5550 3164 5603 3198
rect 5637 3164 5690 3198
rect 5550 3152 5690 3164
rect 6542 4082 6682 4152
rect 6542 4048 6595 4082
rect 6629 4048 6682 4082
rect 6542 4014 6682 4048
rect 6542 3980 6595 4014
rect 6629 3980 6682 4014
rect 6542 3946 6682 3980
rect 6542 3912 6595 3946
rect 6629 3912 6682 3946
rect 6542 3878 6682 3912
rect 6542 3844 6595 3878
rect 6629 3844 6682 3878
rect 6542 3810 6682 3844
rect 6542 3776 6595 3810
rect 6629 3776 6682 3810
rect 6542 3742 6682 3776
rect 6542 3708 6595 3742
rect 6629 3708 6682 3742
rect 6542 3674 6682 3708
rect 6542 3640 6595 3674
rect 6629 3640 6682 3674
rect 6542 3606 6682 3640
rect 6542 3572 6595 3606
rect 6629 3572 6682 3606
rect 6542 3538 6682 3572
rect 6542 3504 6595 3538
rect 6629 3504 6682 3538
rect 6542 3470 6682 3504
rect 6542 3436 6595 3470
rect 6629 3436 6682 3470
rect 6542 3402 6682 3436
rect 6542 3368 6595 3402
rect 6629 3368 6682 3402
rect 6542 3334 6682 3368
rect 6542 3300 6595 3334
rect 6629 3300 6682 3334
rect 6542 3266 6682 3300
rect 6542 3232 6595 3266
rect 6629 3232 6682 3266
rect 6542 3198 6682 3232
rect 6542 3164 6595 3198
rect 6629 3164 6682 3198
rect 6542 3152 6682 3164
rect 7534 4082 7674 4152
rect 7534 4048 7587 4082
rect 7621 4048 7674 4082
rect 7534 4014 7674 4048
rect 7534 3980 7587 4014
rect 7621 3980 7674 4014
rect 7534 3946 7674 3980
rect 7534 3912 7587 3946
rect 7621 3912 7674 3946
rect 7534 3878 7674 3912
rect 7534 3844 7587 3878
rect 7621 3844 7674 3878
rect 7534 3810 7674 3844
rect 7534 3776 7587 3810
rect 7621 3776 7674 3810
rect 7534 3742 7674 3776
rect 7534 3708 7587 3742
rect 7621 3708 7674 3742
rect 7534 3674 7674 3708
rect 7534 3640 7587 3674
rect 7621 3640 7674 3674
rect 7534 3606 7674 3640
rect 7534 3572 7587 3606
rect 7621 3572 7674 3606
rect 7534 3538 7674 3572
rect 7534 3504 7587 3538
rect 7621 3504 7674 3538
rect 7534 3470 7674 3504
rect 7534 3436 7587 3470
rect 7621 3436 7674 3470
rect 7534 3402 7674 3436
rect 7534 3368 7587 3402
rect 7621 3368 7674 3402
rect 7534 3334 7674 3368
rect 7534 3300 7587 3334
rect 7621 3300 7674 3334
rect 7534 3266 7674 3300
rect 7534 3232 7587 3266
rect 7621 3232 7674 3266
rect 7534 3198 7674 3232
rect 7534 3164 7587 3198
rect 7621 3164 7674 3198
rect 7534 3152 7674 3164
rect 8526 4082 8666 4152
rect 8526 4048 8579 4082
rect 8613 4048 8666 4082
rect 8526 4014 8666 4048
rect 8526 3980 8579 4014
rect 8613 3980 8666 4014
rect 8526 3946 8666 3980
rect 8526 3912 8579 3946
rect 8613 3912 8666 3946
rect 8526 3878 8666 3912
rect 8526 3844 8579 3878
rect 8613 3844 8666 3878
rect 8526 3810 8666 3844
rect 8526 3776 8579 3810
rect 8613 3776 8666 3810
rect 8526 3742 8666 3776
rect 8526 3708 8579 3742
rect 8613 3708 8666 3742
rect 8526 3674 8666 3708
rect 8526 3640 8579 3674
rect 8613 3640 8666 3674
rect 8526 3606 8666 3640
rect 8526 3572 8579 3606
rect 8613 3572 8666 3606
rect 8526 3538 8666 3572
rect 8526 3504 8579 3538
rect 8613 3504 8666 3538
rect 8526 3470 8666 3504
rect 8526 3436 8579 3470
rect 8613 3436 8666 3470
rect 8526 3402 8666 3436
rect 8526 3368 8579 3402
rect 8613 3368 8666 3402
rect 8526 3334 8666 3368
rect 8526 3300 8579 3334
rect 8613 3300 8666 3334
rect 8526 3266 8666 3300
rect 8526 3232 8579 3266
rect 8613 3232 8666 3266
rect 8526 3198 8666 3232
rect 8526 3164 8579 3198
rect 8613 3164 8666 3198
rect 8526 3152 8666 3164
rect 9518 4082 9658 4152
rect 9518 4048 9571 4082
rect 9605 4048 9658 4082
rect 9518 4014 9658 4048
rect 9518 3980 9571 4014
rect 9605 3980 9658 4014
rect 9518 3946 9658 3980
rect 9518 3912 9571 3946
rect 9605 3912 9658 3946
rect 9518 3878 9658 3912
rect 9518 3844 9571 3878
rect 9605 3844 9658 3878
rect 9518 3810 9658 3844
rect 9518 3776 9571 3810
rect 9605 3776 9658 3810
rect 9518 3742 9658 3776
rect 9518 3708 9571 3742
rect 9605 3708 9658 3742
rect 9518 3674 9658 3708
rect 9518 3640 9571 3674
rect 9605 3640 9658 3674
rect 9518 3606 9658 3640
rect 9518 3572 9571 3606
rect 9605 3572 9658 3606
rect 9518 3538 9658 3572
rect 9518 3504 9571 3538
rect 9605 3504 9658 3538
rect 9518 3470 9658 3504
rect 9518 3436 9571 3470
rect 9605 3436 9658 3470
rect 9518 3402 9658 3436
rect 9518 3368 9571 3402
rect 9605 3368 9658 3402
rect 9518 3334 9658 3368
rect 9518 3300 9571 3334
rect 9605 3300 9658 3334
rect 9518 3266 9658 3300
rect 9518 3232 9571 3266
rect 9605 3232 9658 3266
rect 9518 3198 9658 3232
rect 9518 3164 9571 3198
rect 9605 3164 9658 3198
rect 9518 3152 9658 3164
rect 10510 4082 10650 4152
rect 10510 4048 10563 4082
rect 10597 4048 10650 4082
rect 10510 4014 10650 4048
rect 10510 3980 10563 4014
rect 10597 3980 10650 4014
rect 10510 3946 10650 3980
rect 10510 3912 10563 3946
rect 10597 3912 10650 3946
rect 10510 3878 10650 3912
rect 10510 3844 10563 3878
rect 10597 3844 10650 3878
rect 10510 3810 10650 3844
rect 10510 3776 10563 3810
rect 10597 3776 10650 3810
rect 10510 3742 10650 3776
rect 10510 3708 10563 3742
rect 10597 3708 10650 3742
rect 10510 3674 10650 3708
rect 10510 3640 10563 3674
rect 10597 3640 10650 3674
rect 10510 3606 10650 3640
rect 10510 3572 10563 3606
rect 10597 3572 10650 3606
rect 10510 3538 10650 3572
rect 10510 3504 10563 3538
rect 10597 3504 10650 3538
rect 10510 3470 10650 3504
rect 10510 3436 10563 3470
rect 10597 3436 10650 3470
rect 10510 3402 10650 3436
rect 10510 3368 10563 3402
rect 10597 3368 10650 3402
rect 10510 3334 10650 3368
rect 10510 3300 10563 3334
rect 10597 3300 10650 3334
rect 10510 3266 10650 3300
rect 10510 3232 10563 3266
rect 10597 3232 10650 3266
rect 10510 3198 10650 3232
rect 10510 3164 10563 3198
rect 10597 3164 10650 3198
rect 10510 3152 10650 3164
rect 11502 4082 11642 4152
rect 11502 4048 11555 4082
rect 11589 4048 11642 4082
rect 11502 4014 11642 4048
rect 11502 3980 11555 4014
rect 11589 3980 11642 4014
rect 11502 3946 11642 3980
rect 11502 3912 11555 3946
rect 11589 3912 11642 3946
rect 11502 3878 11642 3912
rect 11502 3844 11555 3878
rect 11589 3844 11642 3878
rect 11502 3810 11642 3844
rect 11502 3776 11555 3810
rect 11589 3776 11642 3810
rect 11502 3742 11642 3776
rect 11502 3708 11555 3742
rect 11589 3708 11642 3742
rect 11502 3674 11642 3708
rect 11502 3640 11555 3674
rect 11589 3640 11642 3674
rect 11502 3606 11642 3640
rect 11502 3572 11555 3606
rect 11589 3572 11642 3606
rect 11502 3538 11642 3572
rect 11502 3504 11555 3538
rect 11589 3504 11642 3538
rect 11502 3470 11642 3504
rect 11502 3436 11555 3470
rect 11589 3436 11642 3470
rect 11502 3402 11642 3436
rect 11502 3368 11555 3402
rect 11589 3368 11642 3402
rect 11502 3334 11642 3368
rect 11502 3300 11555 3334
rect 11589 3300 11642 3334
rect 11502 3266 11642 3300
rect 11502 3232 11555 3266
rect 11589 3232 11642 3266
rect 11502 3198 11642 3232
rect 11502 3164 11555 3198
rect 11589 3164 11642 3198
rect 11502 3152 11642 3164
rect 12494 4082 12634 4152
rect 12494 4048 12547 4082
rect 12581 4048 12634 4082
rect 12494 4014 12634 4048
rect 12494 3980 12547 4014
rect 12581 3980 12634 4014
rect 12494 3946 12634 3980
rect 12494 3912 12547 3946
rect 12581 3912 12634 3946
rect 12494 3878 12634 3912
rect 12494 3844 12547 3878
rect 12581 3844 12634 3878
rect 12494 3810 12634 3844
rect 12494 3776 12547 3810
rect 12581 3776 12634 3810
rect 12494 3742 12634 3776
rect 12494 3708 12547 3742
rect 12581 3708 12634 3742
rect 12494 3674 12634 3708
rect 12494 3640 12547 3674
rect 12581 3640 12634 3674
rect 12494 3606 12634 3640
rect 12494 3572 12547 3606
rect 12581 3572 12634 3606
rect 12494 3538 12634 3572
rect 12494 3504 12547 3538
rect 12581 3504 12634 3538
rect 12494 3470 12634 3504
rect 12494 3436 12547 3470
rect 12581 3436 12634 3470
rect 12494 3402 12634 3436
rect 12494 3368 12547 3402
rect 12581 3368 12634 3402
rect 12494 3334 12634 3368
rect 12494 3300 12547 3334
rect 12581 3300 12634 3334
rect 12494 3266 12634 3300
rect 12494 3232 12547 3266
rect 12581 3232 12634 3266
rect 12494 3198 12634 3232
rect 12494 3164 12547 3198
rect 12581 3164 12634 3198
rect 12494 3152 12634 3164
rect 13486 4082 13626 4152
rect 13486 4048 13539 4082
rect 13573 4048 13626 4082
rect 13486 4014 13626 4048
rect 13486 3980 13539 4014
rect 13573 3980 13626 4014
rect 13486 3946 13626 3980
rect 13486 3912 13539 3946
rect 13573 3912 13626 3946
rect 13486 3878 13626 3912
rect 13486 3844 13539 3878
rect 13573 3844 13626 3878
rect 13486 3810 13626 3844
rect 13486 3776 13539 3810
rect 13573 3776 13626 3810
rect 13486 3742 13626 3776
rect 13486 3708 13539 3742
rect 13573 3708 13626 3742
rect 13486 3674 13626 3708
rect 13486 3640 13539 3674
rect 13573 3640 13626 3674
rect 13486 3606 13626 3640
rect 13486 3572 13539 3606
rect 13573 3572 13626 3606
rect 13486 3538 13626 3572
rect 13486 3504 13539 3538
rect 13573 3504 13626 3538
rect 13486 3470 13626 3504
rect 13486 3436 13539 3470
rect 13573 3436 13626 3470
rect 13486 3402 13626 3436
rect 13486 3368 13539 3402
rect 13573 3368 13626 3402
rect 13486 3334 13626 3368
rect 13486 3300 13539 3334
rect 13573 3300 13626 3334
rect 13486 3266 13626 3300
rect 13486 3232 13539 3266
rect 13573 3232 13626 3266
rect 13486 3198 13626 3232
rect 13486 3164 13539 3198
rect 13573 3164 13626 3198
rect 13486 3152 13626 3164
rect 14427 3992 14468 4152
rect 14427 3957 14536 3992
rect 14427 3923 14468 3957
rect 14502 3924 14536 3957
rect 14502 3923 14604 3924
rect 14427 3905 14604 3923
rect 14638 3905 14653 4551
rect 14427 3889 14653 3905
rect 14427 3888 14536 3889
rect 14427 3854 14468 3888
rect 14502 3855 14536 3888
rect 14570 3871 14653 3889
rect 14570 3855 14604 3871
rect 14502 3854 14604 3855
rect 14427 3837 14604 3854
rect 14638 3837 14653 3871
rect 14427 3820 14653 3837
rect 14427 3819 14536 3820
rect 14427 3785 14468 3819
rect 14502 3786 14536 3819
rect 14570 3803 14653 3820
rect 14570 3786 14604 3803
rect 14502 3785 14604 3786
rect 14427 3769 14604 3785
rect 14638 3769 14653 3803
rect 14427 3751 14653 3769
rect 14427 3750 14536 3751
rect 14427 3716 14468 3750
rect 14502 3717 14536 3750
rect 14570 3735 14653 3751
rect 14570 3717 14604 3735
rect 14502 3716 14604 3717
rect 14427 3701 14604 3716
rect 14638 3701 14653 3735
rect 14427 3682 14653 3701
rect 14427 3681 14536 3682
rect 14427 3647 14468 3681
rect 14502 3648 14536 3681
rect 14570 3667 14653 3682
rect 14570 3648 14604 3667
rect 14502 3647 14604 3648
rect 14427 3633 14604 3647
rect 14638 3633 14653 3667
rect 14427 3613 14653 3633
rect 14427 3612 14536 3613
rect 14427 3578 14468 3612
rect 14502 3579 14536 3612
rect 14570 3599 14653 3613
rect 14570 3579 14604 3599
rect 14502 3578 14604 3579
rect 14427 3565 14604 3578
rect 14638 3565 14653 3599
rect 14427 3544 14653 3565
rect 14427 3543 14536 3544
rect 14427 3509 14468 3543
rect 14502 3510 14536 3543
rect 14570 3531 14653 3544
rect 14570 3510 14604 3531
rect 14502 3509 14604 3510
rect 14427 3497 14604 3509
rect 14638 3497 14653 3531
rect 14427 3475 14653 3497
rect 14427 3474 14536 3475
rect 14427 3440 14468 3474
rect 14502 3441 14536 3474
rect 14570 3463 14653 3475
rect 14570 3441 14604 3463
rect 14502 3440 14604 3441
rect 14427 3429 14604 3440
rect 14638 3429 14653 3463
rect 14427 3406 14653 3429
rect 14427 3405 14536 3406
rect 14427 3371 14468 3405
rect 14502 3372 14536 3405
rect 14570 3395 14653 3406
rect 14570 3372 14604 3395
rect 14502 3371 14604 3372
rect 14427 3361 14604 3371
rect 14638 3361 14653 3395
rect 14427 3337 14653 3361
rect 14427 3336 14536 3337
rect 14427 3302 14468 3336
rect 14502 3303 14536 3336
rect 14570 3327 14653 3337
rect 14570 3303 14604 3327
rect 14502 3302 14604 3303
rect 14427 3293 14604 3302
rect 14638 3293 14653 3327
rect 14427 3268 14653 3293
rect 14427 3267 14536 3268
rect 14427 3233 14468 3267
rect 14502 3234 14536 3267
rect 14570 3259 14653 3268
rect 14570 3234 14604 3259
rect 14502 3233 14604 3234
rect 14427 3225 14604 3233
rect 14638 3225 14653 3259
rect 14427 3199 14653 3225
rect 14427 3198 14536 3199
rect 14427 3164 14468 3198
rect 14502 3165 14536 3198
rect 14570 3191 14653 3199
rect 14570 3165 14604 3191
rect 14502 3164 14604 3165
rect 14427 3157 14604 3164
rect 14638 3157 14653 3191
rect 14427 3152 14653 3157
rect 482 3128 682 3152
rect 482 3094 497 3128
rect 531 3094 565 3128
rect 599 3094 633 3128
rect 667 3094 682 3128
rect 482 3059 682 3094
rect 482 3025 497 3059
rect 531 3025 565 3059
rect 599 3025 633 3059
rect 667 3025 682 3059
rect 482 2990 682 3025
rect 482 2956 497 2990
rect 531 2956 565 2990
rect 599 2956 633 2990
rect 667 2956 682 2990
rect 482 2921 682 2956
rect 482 2887 497 2921
rect 531 2887 565 2921
rect 599 2887 633 2921
rect 667 2887 682 2921
rect 482 2852 682 2887
rect 482 2818 497 2852
rect 531 2818 565 2852
rect 599 2818 633 2852
rect 667 2818 682 2852
rect 482 2783 682 2818
rect 482 2749 497 2783
rect 531 2749 565 2783
rect 599 2749 633 2783
rect 667 2749 682 2783
rect 482 2714 682 2749
rect 482 2680 497 2714
rect 531 2680 565 2714
rect 599 2680 633 2714
rect 667 2680 682 2714
rect 482 2645 682 2680
rect 482 2611 497 2645
rect 531 2611 565 2645
rect 599 2611 633 2645
rect 667 2611 682 2645
rect 482 2576 682 2611
rect 482 2542 497 2576
rect 531 2542 565 2576
rect 599 2542 633 2576
rect 667 2552 682 2576
rect 1541 3044 1763 3078
rect 1541 3010 1601 3044
rect 1635 3010 1669 3044
rect 1703 3010 1763 3044
rect 1541 2974 1763 3010
rect 1541 2940 1601 2974
rect 1635 2940 1669 2974
rect 1703 2940 1763 2974
rect 1541 2904 1763 2940
rect 1541 2870 1601 2904
rect 1635 2870 1669 2904
rect 1703 2870 1763 2904
rect 1541 2834 1763 2870
rect 1541 2800 1601 2834
rect 1635 2800 1669 2834
rect 1703 2800 1763 2834
rect 1541 2764 1763 2800
rect 1541 2730 1601 2764
rect 1635 2730 1669 2764
rect 1703 2730 1763 2764
rect 1541 2694 1763 2730
rect 1541 2660 1601 2694
rect 1635 2660 1669 2694
rect 1703 2660 1763 2694
rect 1541 2626 1763 2660
rect 2533 3044 2755 3078
rect 2533 3010 2593 3044
rect 2627 3010 2661 3044
rect 2695 3010 2755 3044
rect 2533 2974 2755 3010
rect 2533 2940 2593 2974
rect 2627 2940 2661 2974
rect 2695 2940 2755 2974
rect 2533 2904 2755 2940
rect 2533 2870 2593 2904
rect 2627 2870 2661 2904
rect 2695 2870 2755 2904
rect 2533 2834 2755 2870
rect 2533 2800 2593 2834
rect 2627 2800 2661 2834
rect 2695 2800 2755 2834
rect 2533 2764 2755 2800
rect 2533 2730 2593 2764
rect 2627 2730 2661 2764
rect 2695 2730 2755 2764
rect 2533 2694 2755 2730
rect 2533 2660 2593 2694
rect 2627 2660 2661 2694
rect 2695 2660 2755 2694
rect 2533 2626 2755 2660
rect 3525 3044 3747 3078
rect 3525 3010 3585 3044
rect 3619 3010 3653 3044
rect 3687 3010 3747 3044
rect 3525 2974 3747 3010
rect 3525 2940 3585 2974
rect 3619 2940 3653 2974
rect 3687 2940 3747 2974
rect 3525 2904 3747 2940
rect 3525 2870 3585 2904
rect 3619 2870 3653 2904
rect 3687 2870 3747 2904
rect 3525 2834 3747 2870
rect 3525 2800 3585 2834
rect 3619 2800 3653 2834
rect 3687 2800 3747 2834
rect 3525 2764 3747 2800
rect 3525 2730 3585 2764
rect 3619 2730 3653 2764
rect 3687 2730 3747 2764
rect 3525 2694 3747 2730
rect 3525 2660 3585 2694
rect 3619 2660 3653 2694
rect 3687 2660 3747 2694
rect 3525 2626 3747 2660
rect 4517 3044 4739 3078
rect 4517 3010 4577 3044
rect 4611 3010 4645 3044
rect 4679 3010 4739 3044
rect 4517 2974 4739 3010
rect 4517 2940 4577 2974
rect 4611 2940 4645 2974
rect 4679 2940 4739 2974
rect 4517 2904 4739 2940
rect 4517 2870 4577 2904
rect 4611 2870 4645 2904
rect 4679 2870 4739 2904
rect 4517 2834 4739 2870
rect 4517 2800 4577 2834
rect 4611 2800 4645 2834
rect 4679 2800 4739 2834
rect 4517 2764 4739 2800
rect 4517 2730 4577 2764
rect 4611 2730 4645 2764
rect 4679 2730 4739 2764
rect 4517 2694 4739 2730
rect 4517 2660 4577 2694
rect 4611 2660 4645 2694
rect 4679 2660 4739 2694
rect 4517 2626 4739 2660
rect 5509 3044 5731 3078
rect 5509 3010 5569 3044
rect 5603 3010 5637 3044
rect 5671 3010 5731 3044
rect 5509 2974 5731 3010
rect 5509 2940 5569 2974
rect 5603 2940 5637 2974
rect 5671 2940 5731 2974
rect 5509 2904 5731 2940
rect 5509 2870 5569 2904
rect 5603 2870 5637 2904
rect 5671 2870 5731 2904
rect 5509 2834 5731 2870
rect 5509 2800 5569 2834
rect 5603 2800 5637 2834
rect 5671 2800 5731 2834
rect 5509 2764 5731 2800
rect 5509 2730 5569 2764
rect 5603 2730 5637 2764
rect 5671 2730 5731 2764
rect 5509 2694 5731 2730
rect 5509 2660 5569 2694
rect 5603 2660 5637 2694
rect 5671 2660 5731 2694
rect 5509 2626 5731 2660
rect 6501 3044 6723 3078
rect 6501 3010 6561 3044
rect 6595 3010 6629 3044
rect 6663 3010 6723 3044
rect 6501 2974 6723 3010
rect 6501 2940 6561 2974
rect 6595 2940 6629 2974
rect 6663 2940 6723 2974
rect 6501 2904 6723 2940
rect 6501 2870 6561 2904
rect 6595 2870 6629 2904
rect 6663 2870 6723 2904
rect 6501 2834 6723 2870
rect 6501 2800 6561 2834
rect 6595 2800 6629 2834
rect 6663 2800 6723 2834
rect 6501 2764 6723 2800
rect 6501 2730 6561 2764
rect 6595 2730 6629 2764
rect 6663 2730 6723 2764
rect 6501 2694 6723 2730
rect 6501 2660 6561 2694
rect 6595 2660 6629 2694
rect 6663 2660 6723 2694
rect 6501 2626 6723 2660
rect 7493 3044 7715 3078
rect 7493 3010 7553 3044
rect 7587 3010 7621 3044
rect 7655 3010 7715 3044
rect 7493 2974 7715 3010
rect 7493 2940 7553 2974
rect 7587 2940 7621 2974
rect 7655 2940 7715 2974
rect 7493 2904 7715 2940
rect 7493 2870 7553 2904
rect 7587 2870 7621 2904
rect 7655 2870 7715 2904
rect 7493 2834 7715 2870
rect 7493 2800 7553 2834
rect 7587 2800 7621 2834
rect 7655 2800 7715 2834
rect 7493 2764 7715 2800
rect 7493 2730 7553 2764
rect 7587 2730 7621 2764
rect 7655 2730 7715 2764
rect 7493 2694 7715 2730
rect 7493 2660 7553 2694
rect 7587 2660 7621 2694
rect 7655 2660 7715 2694
rect 7493 2626 7715 2660
rect 8485 3044 8707 3078
rect 8485 3010 8545 3044
rect 8579 3010 8613 3044
rect 8647 3010 8707 3044
rect 8485 2974 8707 3010
rect 8485 2940 8545 2974
rect 8579 2940 8613 2974
rect 8647 2940 8707 2974
rect 8485 2904 8707 2940
rect 8485 2870 8545 2904
rect 8579 2870 8613 2904
rect 8647 2870 8707 2904
rect 8485 2834 8707 2870
rect 8485 2800 8545 2834
rect 8579 2800 8613 2834
rect 8647 2800 8707 2834
rect 8485 2764 8707 2800
rect 8485 2730 8545 2764
rect 8579 2730 8613 2764
rect 8647 2730 8707 2764
rect 8485 2694 8707 2730
rect 8485 2660 8545 2694
rect 8579 2660 8613 2694
rect 8647 2660 8707 2694
rect 8485 2626 8707 2660
rect 9477 3044 9699 3078
rect 9477 3010 9537 3044
rect 9571 3010 9605 3044
rect 9639 3010 9699 3044
rect 9477 2974 9699 3010
rect 9477 2940 9537 2974
rect 9571 2940 9605 2974
rect 9639 2940 9699 2974
rect 9477 2904 9699 2940
rect 9477 2870 9537 2904
rect 9571 2870 9605 2904
rect 9639 2870 9699 2904
rect 9477 2834 9699 2870
rect 9477 2800 9537 2834
rect 9571 2800 9605 2834
rect 9639 2800 9699 2834
rect 9477 2764 9699 2800
rect 9477 2730 9537 2764
rect 9571 2730 9605 2764
rect 9639 2730 9699 2764
rect 9477 2694 9699 2730
rect 9477 2660 9537 2694
rect 9571 2660 9605 2694
rect 9639 2660 9699 2694
rect 9477 2626 9699 2660
rect 10469 3044 10691 3078
rect 10469 3010 10529 3044
rect 10563 3010 10597 3044
rect 10631 3010 10691 3044
rect 10469 2974 10691 3010
rect 10469 2940 10529 2974
rect 10563 2940 10597 2974
rect 10631 2940 10691 2974
rect 10469 2904 10691 2940
rect 10469 2870 10529 2904
rect 10563 2870 10597 2904
rect 10631 2870 10691 2904
rect 10469 2834 10691 2870
rect 10469 2800 10529 2834
rect 10563 2800 10597 2834
rect 10631 2800 10691 2834
rect 10469 2764 10691 2800
rect 10469 2730 10529 2764
rect 10563 2730 10597 2764
rect 10631 2730 10691 2764
rect 10469 2694 10691 2730
rect 10469 2660 10529 2694
rect 10563 2660 10597 2694
rect 10631 2660 10691 2694
rect 10469 2626 10691 2660
rect 11461 3044 11683 3078
rect 11461 3010 11521 3044
rect 11555 3010 11589 3044
rect 11623 3010 11683 3044
rect 11461 2974 11683 3010
rect 11461 2940 11521 2974
rect 11555 2940 11589 2974
rect 11623 2940 11683 2974
rect 11461 2904 11683 2940
rect 11461 2870 11521 2904
rect 11555 2870 11589 2904
rect 11623 2870 11683 2904
rect 11461 2834 11683 2870
rect 11461 2800 11521 2834
rect 11555 2800 11589 2834
rect 11623 2800 11683 2834
rect 11461 2764 11683 2800
rect 11461 2730 11521 2764
rect 11555 2730 11589 2764
rect 11623 2730 11683 2764
rect 11461 2694 11683 2730
rect 11461 2660 11521 2694
rect 11555 2660 11589 2694
rect 11623 2660 11683 2694
rect 11461 2626 11683 2660
rect 12453 3044 12675 3078
rect 12453 3010 12513 3044
rect 12547 3010 12581 3044
rect 12615 3010 12675 3044
rect 12453 2974 12675 3010
rect 12453 2940 12513 2974
rect 12547 2940 12581 2974
rect 12615 2940 12675 2974
rect 12453 2904 12675 2940
rect 12453 2870 12513 2904
rect 12547 2870 12581 2904
rect 12615 2870 12675 2904
rect 12453 2834 12675 2870
rect 12453 2800 12513 2834
rect 12547 2800 12581 2834
rect 12615 2800 12675 2834
rect 12453 2764 12675 2800
rect 12453 2730 12513 2764
rect 12547 2730 12581 2764
rect 12615 2730 12675 2764
rect 12453 2694 12675 2730
rect 12453 2660 12513 2694
rect 12547 2660 12581 2694
rect 12615 2660 12675 2694
rect 12453 2626 12675 2660
rect 13445 3044 13667 3078
rect 13445 3010 13505 3044
rect 13539 3010 13573 3044
rect 13607 3010 13667 3044
rect 13445 2974 13667 3010
rect 13445 2940 13505 2974
rect 13539 2940 13573 2974
rect 13607 2940 13667 2974
rect 13445 2904 13667 2940
rect 13445 2870 13505 2904
rect 13539 2870 13573 2904
rect 13607 2870 13667 2904
rect 13445 2834 13667 2870
rect 13445 2800 13505 2834
rect 13539 2800 13573 2834
rect 13607 2800 13667 2834
rect 13445 2764 13667 2800
rect 13445 2730 13505 2764
rect 13539 2730 13573 2764
rect 13607 2730 13667 2764
rect 13445 2694 13667 2730
rect 13445 2660 13505 2694
rect 13539 2660 13573 2694
rect 13607 2660 13667 2694
rect 13445 2626 13667 2660
rect 14453 3130 14653 3152
rect 14453 3129 14536 3130
rect 14453 3095 14468 3129
rect 14502 3096 14536 3129
rect 14570 3123 14653 3130
rect 14570 3096 14604 3123
rect 14502 3095 14604 3096
rect 14453 3089 14604 3095
rect 14638 3089 14653 3123
rect 14453 3061 14653 3089
rect 14453 3060 14536 3061
rect 14453 3026 14468 3060
rect 14502 3027 14536 3060
rect 14570 3055 14653 3061
rect 14570 3027 14604 3055
rect 14502 3026 14604 3027
rect 14453 3021 14604 3026
rect 14638 3021 14653 3055
rect 14453 2992 14653 3021
rect 14453 2991 14536 2992
rect 14453 2957 14468 2991
rect 14502 2958 14536 2991
rect 14570 2987 14653 2992
rect 14570 2958 14604 2987
rect 14502 2957 14604 2958
rect 14453 2953 14604 2957
rect 14638 2953 14653 2987
rect 14453 2923 14653 2953
rect 14453 2922 14536 2923
rect 14453 2888 14468 2922
rect 14502 2889 14536 2922
rect 14570 2919 14653 2923
rect 14570 2889 14604 2919
rect 14502 2888 14604 2889
rect 14453 2885 14604 2888
rect 14638 2885 14653 2919
rect 14453 2854 14653 2885
rect 14453 2853 14536 2854
rect 14453 2819 14468 2853
rect 14502 2820 14536 2853
rect 14570 2851 14653 2854
rect 14570 2820 14604 2851
rect 14502 2819 14604 2820
rect 14453 2817 14604 2819
rect 14638 2817 14653 2851
rect 14453 2785 14653 2817
rect 14453 2784 14536 2785
rect 14453 2750 14468 2784
rect 14502 2751 14536 2784
rect 14570 2783 14653 2785
rect 14570 2751 14604 2783
rect 14502 2750 14604 2751
rect 14453 2749 14604 2750
rect 14638 2749 14653 2783
rect 14453 2716 14653 2749
rect 14453 2715 14536 2716
rect 14453 2681 14468 2715
rect 14502 2682 14536 2715
rect 14570 2715 14653 2716
rect 14570 2682 14604 2715
rect 14502 2681 14604 2682
rect 14638 2681 14653 2715
rect 14453 2647 14653 2681
rect 14453 2646 14536 2647
rect 14453 2612 14468 2646
rect 14502 2613 14536 2646
rect 14570 2613 14604 2647
rect 14638 2613 14653 2647
rect 14502 2612 14653 2613
rect 14453 2579 14653 2612
rect 14453 2578 14604 2579
rect 14453 2577 14536 2578
rect 14453 2552 14468 2577
rect 667 2542 708 2552
rect 482 2507 708 2542
rect 482 2473 497 2507
rect 531 2473 565 2507
rect 599 2473 633 2507
rect 667 2473 708 2507
rect 482 2438 708 2473
rect 482 2404 497 2438
rect 531 2404 565 2438
rect 599 2404 633 2438
rect 667 2404 708 2438
rect 482 2369 708 2404
rect 482 2335 497 2369
rect 531 2335 565 2369
rect 599 2335 633 2369
rect 667 2335 708 2369
rect 482 2300 708 2335
rect 482 2266 497 2300
rect 531 2266 565 2300
rect 599 2266 633 2300
rect 667 2266 708 2300
rect 482 2231 708 2266
rect 482 2197 497 2231
rect 531 2197 565 2231
rect 599 2197 633 2231
rect 667 2197 708 2231
rect 482 2163 708 2197
rect 482 2129 497 2163
rect 531 2162 708 2163
rect 531 2129 565 2162
rect 482 2128 565 2129
rect 599 2128 633 2162
rect 667 2128 708 2162
rect 482 2095 708 2128
rect 482 2061 497 2095
rect 531 2093 708 2095
rect 531 2061 565 2093
rect 482 2059 565 2061
rect 599 2059 633 2093
rect 667 2059 708 2093
rect 482 2027 708 2059
rect 482 1993 497 2027
rect 531 2024 708 2027
rect 531 1993 565 2024
rect 482 1990 565 1993
rect 599 1990 633 2024
rect 667 1990 708 2024
rect 482 1959 708 1990
rect 482 1925 497 1959
rect 531 1955 708 1959
rect 531 1925 565 1955
rect 482 1921 565 1925
rect 599 1921 633 1955
rect 667 1921 708 1955
rect 482 1891 708 1921
rect 482 1857 497 1891
rect 531 1886 708 1891
rect 531 1857 565 1886
rect 482 1852 565 1857
rect 599 1852 633 1886
rect 667 1852 708 1886
rect 482 1823 708 1852
rect 482 1789 497 1823
rect 531 1817 708 1823
rect 531 1789 565 1817
rect 482 1783 565 1789
rect 599 1783 633 1817
rect 667 1783 708 1817
rect 482 1755 708 1783
rect 482 1721 497 1755
rect 531 1748 708 1755
rect 531 1721 565 1748
rect 482 1714 565 1721
rect 599 1714 633 1748
rect 667 1714 708 1748
rect 482 1687 708 1714
rect 482 1653 497 1687
rect 531 1679 708 1687
rect 531 1653 565 1679
rect 482 1645 565 1653
rect 599 1645 633 1679
rect 667 1645 708 1679
rect 482 1619 708 1645
rect 482 1585 497 1619
rect 531 1610 708 1619
rect 531 1585 565 1610
rect 482 1576 565 1585
rect 599 1576 633 1610
rect 667 1576 708 1610
rect 482 1552 708 1576
rect 1582 2540 1722 2552
rect 1582 2506 1635 2540
rect 1669 2506 1722 2540
rect 1582 2472 1722 2506
rect 1582 2438 1635 2472
rect 1669 2438 1722 2472
rect 1582 2404 1722 2438
rect 1582 2370 1635 2404
rect 1669 2370 1722 2404
rect 1582 2336 1722 2370
rect 1582 2302 1635 2336
rect 1669 2302 1722 2336
rect 1582 2268 1722 2302
rect 1582 2234 1635 2268
rect 1669 2234 1722 2268
rect 1582 2200 1722 2234
rect 1582 2166 1635 2200
rect 1669 2166 1722 2200
rect 1582 2132 1722 2166
rect 1582 2098 1635 2132
rect 1669 2098 1722 2132
rect 1582 2064 1722 2098
rect 1582 2030 1635 2064
rect 1669 2030 1722 2064
rect 1582 1996 1722 2030
rect 1582 1962 1635 1996
rect 1669 1962 1722 1996
rect 1582 1928 1722 1962
rect 1582 1894 1635 1928
rect 1669 1894 1722 1928
rect 1582 1860 1722 1894
rect 1582 1826 1635 1860
rect 1669 1826 1722 1860
rect 1582 1792 1722 1826
rect 1582 1758 1635 1792
rect 1669 1758 1722 1792
rect 1582 1724 1722 1758
rect 1582 1690 1635 1724
rect 1669 1690 1722 1724
rect 1582 1656 1722 1690
rect 1582 1622 1635 1656
rect 1669 1622 1722 1656
rect 1582 1552 1722 1622
rect 2574 2540 2714 2552
rect 2574 2506 2627 2540
rect 2661 2506 2714 2540
rect 2574 2472 2714 2506
rect 2574 2438 2627 2472
rect 2661 2438 2714 2472
rect 2574 2404 2714 2438
rect 2574 2370 2627 2404
rect 2661 2370 2714 2404
rect 2574 2336 2714 2370
rect 2574 2302 2627 2336
rect 2661 2302 2714 2336
rect 2574 2268 2714 2302
rect 2574 2234 2627 2268
rect 2661 2234 2714 2268
rect 2574 2200 2714 2234
rect 2574 2166 2627 2200
rect 2661 2166 2714 2200
rect 2574 2132 2714 2166
rect 2574 2098 2627 2132
rect 2661 2098 2714 2132
rect 2574 2064 2714 2098
rect 2574 2030 2627 2064
rect 2661 2030 2714 2064
rect 2574 1996 2714 2030
rect 2574 1962 2627 1996
rect 2661 1962 2714 1996
rect 2574 1928 2714 1962
rect 2574 1894 2627 1928
rect 2661 1894 2714 1928
rect 2574 1860 2714 1894
rect 2574 1826 2627 1860
rect 2661 1826 2714 1860
rect 2574 1792 2714 1826
rect 2574 1758 2627 1792
rect 2661 1758 2714 1792
rect 2574 1724 2714 1758
rect 2574 1690 2627 1724
rect 2661 1690 2714 1724
rect 2574 1656 2714 1690
rect 2574 1622 2627 1656
rect 2661 1622 2714 1656
rect 2574 1552 2714 1622
rect 3566 2540 3706 2552
rect 3566 2506 3619 2540
rect 3653 2506 3706 2540
rect 3566 2472 3706 2506
rect 3566 2438 3619 2472
rect 3653 2438 3706 2472
rect 3566 2404 3706 2438
rect 3566 2370 3619 2404
rect 3653 2370 3706 2404
rect 3566 2336 3706 2370
rect 3566 2302 3619 2336
rect 3653 2302 3706 2336
rect 3566 2268 3706 2302
rect 3566 2234 3619 2268
rect 3653 2234 3706 2268
rect 3566 2200 3706 2234
rect 3566 2166 3619 2200
rect 3653 2166 3706 2200
rect 3566 2132 3706 2166
rect 3566 2098 3619 2132
rect 3653 2098 3706 2132
rect 3566 2064 3706 2098
rect 3566 2030 3619 2064
rect 3653 2030 3706 2064
rect 3566 1996 3706 2030
rect 3566 1962 3619 1996
rect 3653 1962 3706 1996
rect 3566 1928 3706 1962
rect 3566 1894 3619 1928
rect 3653 1894 3706 1928
rect 3566 1860 3706 1894
rect 3566 1826 3619 1860
rect 3653 1826 3706 1860
rect 3566 1792 3706 1826
rect 3566 1758 3619 1792
rect 3653 1758 3706 1792
rect 3566 1724 3706 1758
rect 3566 1690 3619 1724
rect 3653 1690 3706 1724
rect 3566 1656 3706 1690
rect 3566 1622 3619 1656
rect 3653 1622 3706 1656
rect 3566 1552 3706 1622
rect 4558 2540 4698 2552
rect 4558 2506 4611 2540
rect 4645 2506 4698 2540
rect 4558 2472 4698 2506
rect 4558 2438 4611 2472
rect 4645 2438 4698 2472
rect 4558 2404 4698 2438
rect 4558 2370 4611 2404
rect 4645 2370 4698 2404
rect 4558 2336 4698 2370
rect 4558 2302 4611 2336
rect 4645 2302 4698 2336
rect 4558 2268 4698 2302
rect 4558 2234 4611 2268
rect 4645 2234 4698 2268
rect 4558 2200 4698 2234
rect 4558 2166 4611 2200
rect 4645 2166 4698 2200
rect 4558 2132 4698 2166
rect 4558 2098 4611 2132
rect 4645 2098 4698 2132
rect 4558 2064 4698 2098
rect 4558 2030 4611 2064
rect 4645 2030 4698 2064
rect 4558 1996 4698 2030
rect 4558 1962 4611 1996
rect 4645 1962 4698 1996
rect 4558 1928 4698 1962
rect 4558 1894 4611 1928
rect 4645 1894 4698 1928
rect 4558 1860 4698 1894
rect 4558 1826 4611 1860
rect 4645 1826 4698 1860
rect 4558 1792 4698 1826
rect 4558 1758 4611 1792
rect 4645 1758 4698 1792
rect 4558 1724 4698 1758
rect 4558 1690 4611 1724
rect 4645 1690 4698 1724
rect 4558 1656 4698 1690
rect 4558 1622 4611 1656
rect 4645 1622 4698 1656
rect 4558 1552 4698 1622
rect 5550 2540 5690 2552
rect 5550 2506 5603 2540
rect 5637 2506 5690 2540
rect 5550 2472 5690 2506
rect 5550 2438 5603 2472
rect 5637 2438 5690 2472
rect 5550 2404 5690 2438
rect 5550 2370 5603 2404
rect 5637 2370 5690 2404
rect 5550 2336 5690 2370
rect 5550 2302 5603 2336
rect 5637 2302 5690 2336
rect 5550 2268 5690 2302
rect 5550 2234 5603 2268
rect 5637 2234 5690 2268
rect 5550 2200 5690 2234
rect 5550 2166 5603 2200
rect 5637 2166 5690 2200
rect 5550 2132 5690 2166
rect 5550 2098 5603 2132
rect 5637 2098 5690 2132
rect 5550 2064 5690 2098
rect 5550 2030 5603 2064
rect 5637 2030 5690 2064
rect 5550 1996 5690 2030
rect 5550 1962 5603 1996
rect 5637 1962 5690 1996
rect 5550 1928 5690 1962
rect 5550 1894 5603 1928
rect 5637 1894 5690 1928
rect 5550 1860 5690 1894
rect 5550 1826 5603 1860
rect 5637 1826 5690 1860
rect 5550 1792 5690 1826
rect 5550 1758 5603 1792
rect 5637 1758 5690 1792
rect 5550 1724 5690 1758
rect 5550 1690 5603 1724
rect 5637 1690 5690 1724
rect 5550 1656 5690 1690
rect 5550 1622 5603 1656
rect 5637 1622 5690 1656
rect 5550 1552 5690 1622
rect 6542 2540 6682 2552
rect 6542 2506 6595 2540
rect 6629 2506 6682 2540
rect 6542 2472 6682 2506
rect 6542 2438 6595 2472
rect 6629 2438 6682 2472
rect 6542 2404 6682 2438
rect 6542 2370 6595 2404
rect 6629 2370 6682 2404
rect 6542 2336 6682 2370
rect 6542 2302 6595 2336
rect 6629 2302 6682 2336
rect 6542 2268 6682 2302
rect 6542 2234 6595 2268
rect 6629 2234 6682 2268
rect 6542 2200 6682 2234
rect 6542 2166 6595 2200
rect 6629 2166 6682 2200
rect 6542 2132 6682 2166
rect 6542 2098 6595 2132
rect 6629 2098 6682 2132
rect 6542 2064 6682 2098
rect 6542 2030 6595 2064
rect 6629 2030 6682 2064
rect 6542 1996 6682 2030
rect 6542 1962 6595 1996
rect 6629 1962 6682 1996
rect 6542 1928 6682 1962
rect 6542 1894 6595 1928
rect 6629 1894 6682 1928
rect 6542 1860 6682 1894
rect 6542 1826 6595 1860
rect 6629 1826 6682 1860
rect 6542 1792 6682 1826
rect 6542 1758 6595 1792
rect 6629 1758 6682 1792
rect 6542 1724 6682 1758
rect 6542 1690 6595 1724
rect 6629 1690 6682 1724
rect 6542 1656 6682 1690
rect 6542 1622 6595 1656
rect 6629 1622 6682 1656
rect 6542 1552 6682 1622
rect 7534 2540 7674 2552
rect 7534 2506 7587 2540
rect 7621 2506 7674 2540
rect 7534 2472 7674 2506
rect 7534 2438 7587 2472
rect 7621 2438 7674 2472
rect 7534 2404 7674 2438
rect 7534 2370 7587 2404
rect 7621 2370 7674 2404
rect 7534 2336 7674 2370
rect 7534 2302 7587 2336
rect 7621 2302 7674 2336
rect 7534 2268 7674 2302
rect 7534 2234 7587 2268
rect 7621 2234 7674 2268
rect 7534 2200 7674 2234
rect 7534 2166 7587 2200
rect 7621 2166 7674 2200
rect 7534 2132 7674 2166
rect 7534 2098 7587 2132
rect 7621 2098 7674 2132
rect 7534 2064 7674 2098
rect 7534 2030 7587 2064
rect 7621 2030 7674 2064
rect 7534 1996 7674 2030
rect 7534 1962 7587 1996
rect 7621 1962 7674 1996
rect 7534 1928 7674 1962
rect 7534 1894 7587 1928
rect 7621 1894 7674 1928
rect 7534 1860 7674 1894
rect 7534 1826 7587 1860
rect 7621 1826 7674 1860
rect 7534 1792 7674 1826
rect 7534 1758 7587 1792
rect 7621 1758 7674 1792
rect 7534 1724 7674 1758
rect 7534 1690 7587 1724
rect 7621 1690 7674 1724
rect 7534 1656 7674 1690
rect 7534 1622 7587 1656
rect 7621 1622 7674 1656
rect 7534 1552 7674 1622
rect 8526 2540 8666 2552
rect 8526 2506 8579 2540
rect 8613 2506 8666 2540
rect 8526 2472 8666 2506
rect 8526 2438 8579 2472
rect 8613 2438 8666 2472
rect 8526 2404 8666 2438
rect 8526 2370 8579 2404
rect 8613 2370 8666 2404
rect 8526 2336 8666 2370
rect 8526 2302 8579 2336
rect 8613 2302 8666 2336
rect 8526 2268 8666 2302
rect 8526 2234 8579 2268
rect 8613 2234 8666 2268
rect 8526 2200 8666 2234
rect 8526 2166 8579 2200
rect 8613 2166 8666 2200
rect 8526 2132 8666 2166
rect 8526 2098 8579 2132
rect 8613 2098 8666 2132
rect 8526 2064 8666 2098
rect 8526 2030 8579 2064
rect 8613 2030 8666 2064
rect 8526 1996 8666 2030
rect 8526 1962 8579 1996
rect 8613 1962 8666 1996
rect 8526 1928 8666 1962
rect 8526 1894 8579 1928
rect 8613 1894 8666 1928
rect 8526 1860 8666 1894
rect 8526 1826 8579 1860
rect 8613 1826 8666 1860
rect 8526 1792 8666 1826
rect 8526 1758 8579 1792
rect 8613 1758 8666 1792
rect 8526 1724 8666 1758
rect 8526 1690 8579 1724
rect 8613 1690 8666 1724
rect 8526 1656 8666 1690
rect 8526 1622 8579 1656
rect 8613 1622 8666 1656
rect 8526 1552 8666 1622
rect 9518 2540 9658 2552
rect 9518 2506 9571 2540
rect 9605 2506 9658 2540
rect 9518 2472 9658 2506
rect 9518 2438 9571 2472
rect 9605 2438 9658 2472
rect 9518 2404 9658 2438
rect 9518 2370 9571 2404
rect 9605 2370 9658 2404
rect 9518 2336 9658 2370
rect 9518 2302 9571 2336
rect 9605 2302 9658 2336
rect 9518 2268 9658 2302
rect 9518 2234 9571 2268
rect 9605 2234 9658 2268
rect 9518 2200 9658 2234
rect 9518 2166 9571 2200
rect 9605 2166 9658 2200
rect 9518 2132 9658 2166
rect 9518 2098 9571 2132
rect 9605 2098 9658 2132
rect 9518 2064 9658 2098
rect 9518 2030 9571 2064
rect 9605 2030 9658 2064
rect 9518 1996 9658 2030
rect 9518 1962 9571 1996
rect 9605 1962 9658 1996
rect 9518 1928 9658 1962
rect 9518 1894 9571 1928
rect 9605 1894 9658 1928
rect 9518 1860 9658 1894
rect 9518 1826 9571 1860
rect 9605 1826 9658 1860
rect 9518 1792 9658 1826
rect 9518 1758 9571 1792
rect 9605 1758 9658 1792
rect 9518 1724 9658 1758
rect 9518 1690 9571 1724
rect 9605 1690 9658 1724
rect 9518 1656 9658 1690
rect 9518 1622 9571 1656
rect 9605 1622 9658 1656
rect 9518 1552 9658 1622
rect 10510 2540 10650 2552
rect 10510 2506 10563 2540
rect 10597 2506 10650 2540
rect 10510 2472 10650 2506
rect 10510 2438 10563 2472
rect 10597 2438 10650 2472
rect 10510 2404 10650 2438
rect 10510 2370 10563 2404
rect 10597 2370 10650 2404
rect 10510 2336 10650 2370
rect 10510 2302 10563 2336
rect 10597 2302 10650 2336
rect 10510 2268 10650 2302
rect 10510 2234 10563 2268
rect 10597 2234 10650 2268
rect 10510 2200 10650 2234
rect 10510 2166 10563 2200
rect 10597 2166 10650 2200
rect 10510 2132 10650 2166
rect 10510 2098 10563 2132
rect 10597 2098 10650 2132
rect 10510 2064 10650 2098
rect 10510 2030 10563 2064
rect 10597 2030 10650 2064
rect 10510 1996 10650 2030
rect 10510 1962 10563 1996
rect 10597 1962 10650 1996
rect 10510 1928 10650 1962
rect 10510 1894 10563 1928
rect 10597 1894 10650 1928
rect 10510 1860 10650 1894
rect 10510 1826 10563 1860
rect 10597 1826 10650 1860
rect 10510 1792 10650 1826
rect 10510 1758 10563 1792
rect 10597 1758 10650 1792
rect 10510 1724 10650 1758
rect 10510 1690 10563 1724
rect 10597 1690 10650 1724
rect 10510 1656 10650 1690
rect 10510 1622 10563 1656
rect 10597 1622 10650 1656
rect 10510 1552 10650 1622
rect 11502 2540 11642 2552
rect 11502 2506 11555 2540
rect 11589 2506 11642 2540
rect 11502 2472 11642 2506
rect 11502 2438 11555 2472
rect 11589 2438 11642 2472
rect 11502 2404 11642 2438
rect 11502 2370 11555 2404
rect 11589 2370 11642 2404
rect 11502 2336 11642 2370
rect 11502 2302 11555 2336
rect 11589 2302 11642 2336
rect 11502 2268 11642 2302
rect 11502 2234 11555 2268
rect 11589 2234 11642 2268
rect 11502 2200 11642 2234
rect 11502 2166 11555 2200
rect 11589 2166 11642 2200
rect 11502 2132 11642 2166
rect 11502 2098 11555 2132
rect 11589 2098 11642 2132
rect 11502 2064 11642 2098
rect 11502 2030 11555 2064
rect 11589 2030 11642 2064
rect 11502 1996 11642 2030
rect 11502 1962 11555 1996
rect 11589 1962 11642 1996
rect 11502 1928 11642 1962
rect 11502 1894 11555 1928
rect 11589 1894 11642 1928
rect 11502 1860 11642 1894
rect 11502 1826 11555 1860
rect 11589 1826 11642 1860
rect 11502 1792 11642 1826
rect 11502 1758 11555 1792
rect 11589 1758 11642 1792
rect 11502 1724 11642 1758
rect 11502 1690 11555 1724
rect 11589 1690 11642 1724
rect 11502 1656 11642 1690
rect 11502 1622 11555 1656
rect 11589 1622 11642 1656
rect 11502 1552 11642 1622
rect 12494 2540 12634 2552
rect 12494 2506 12547 2540
rect 12581 2506 12634 2540
rect 12494 2472 12634 2506
rect 12494 2438 12547 2472
rect 12581 2438 12634 2472
rect 12494 2404 12634 2438
rect 12494 2370 12547 2404
rect 12581 2370 12634 2404
rect 12494 2336 12634 2370
rect 12494 2302 12547 2336
rect 12581 2302 12634 2336
rect 12494 2268 12634 2302
rect 12494 2234 12547 2268
rect 12581 2234 12634 2268
rect 12494 2200 12634 2234
rect 12494 2166 12547 2200
rect 12581 2166 12634 2200
rect 12494 2132 12634 2166
rect 12494 2098 12547 2132
rect 12581 2098 12634 2132
rect 12494 2064 12634 2098
rect 12494 2030 12547 2064
rect 12581 2030 12634 2064
rect 12494 1996 12634 2030
rect 12494 1962 12547 1996
rect 12581 1962 12634 1996
rect 12494 1928 12634 1962
rect 12494 1894 12547 1928
rect 12581 1894 12634 1928
rect 12494 1860 12634 1894
rect 12494 1826 12547 1860
rect 12581 1826 12634 1860
rect 12494 1792 12634 1826
rect 12494 1758 12547 1792
rect 12581 1758 12634 1792
rect 12494 1724 12634 1758
rect 12494 1690 12547 1724
rect 12581 1690 12634 1724
rect 12494 1656 12634 1690
rect 12494 1622 12547 1656
rect 12581 1622 12634 1656
rect 12494 1552 12634 1622
rect 13486 2540 13626 2552
rect 13486 2506 13539 2540
rect 13573 2506 13626 2540
rect 13486 2472 13626 2506
rect 13486 2438 13539 2472
rect 13573 2438 13626 2472
rect 13486 2404 13626 2438
rect 13486 2370 13539 2404
rect 13573 2370 13626 2404
rect 13486 2336 13626 2370
rect 13486 2302 13539 2336
rect 13573 2302 13626 2336
rect 13486 2268 13626 2302
rect 13486 2234 13539 2268
rect 13573 2234 13626 2268
rect 13486 2200 13626 2234
rect 13486 2166 13539 2200
rect 13573 2166 13626 2200
rect 13486 2132 13626 2166
rect 13486 2098 13539 2132
rect 13573 2098 13626 2132
rect 13486 2064 13626 2098
rect 13486 2030 13539 2064
rect 13573 2030 13626 2064
rect 13486 1996 13626 2030
rect 13486 1962 13539 1996
rect 13573 1962 13626 1996
rect 13486 1928 13626 1962
rect 13486 1894 13539 1928
rect 13573 1894 13626 1928
rect 13486 1860 13626 1894
rect 13486 1826 13539 1860
rect 13573 1826 13626 1860
rect 13486 1792 13626 1826
rect 13486 1758 13539 1792
rect 13573 1758 13626 1792
rect 13486 1724 13626 1758
rect 13486 1690 13539 1724
rect 13573 1690 13626 1724
rect 13486 1656 13626 1690
rect 13486 1622 13539 1656
rect 13573 1622 13626 1656
rect 13486 1552 13626 1622
rect 14427 2543 14468 2552
rect 14502 2544 14536 2577
rect 14570 2545 14604 2578
rect 14638 2545 14653 2579
rect 14570 2544 14653 2545
rect 14502 2543 14653 2544
rect 14427 2511 14653 2543
rect 14427 2509 14604 2511
rect 14427 2508 14536 2509
rect 14427 2474 14468 2508
rect 14502 2475 14536 2508
rect 14570 2477 14604 2509
rect 14638 2477 14653 2511
rect 14570 2475 14653 2477
rect 14502 2474 14653 2475
rect 14427 2443 14653 2474
rect 14427 2440 14604 2443
rect 14427 2439 14536 2440
rect 14427 2405 14468 2439
rect 14502 2406 14536 2439
rect 14570 2409 14604 2440
rect 14638 2409 14653 2443
rect 14570 2406 14653 2409
rect 14502 2405 14653 2406
rect 14427 2375 14653 2405
rect 14427 2371 14604 2375
rect 14427 2370 14536 2371
rect 14427 2336 14468 2370
rect 14502 2337 14536 2370
rect 14570 2341 14604 2371
rect 14638 2341 14653 2375
rect 14570 2337 14653 2341
rect 14502 2336 14653 2337
rect 14427 2307 14653 2336
rect 14427 2302 14604 2307
rect 14427 2301 14536 2302
rect 14427 2267 14468 2301
rect 14502 2268 14536 2301
rect 14570 2273 14604 2302
rect 14638 2273 14653 2307
rect 14570 2268 14653 2273
rect 14502 2267 14653 2268
rect 14427 2239 14653 2267
rect 14427 2233 14604 2239
rect 14427 2232 14536 2233
rect 14427 2198 14468 2232
rect 14502 2199 14536 2232
rect 14570 2205 14604 2233
rect 14638 2205 14653 2239
rect 14570 2199 14653 2205
rect 14502 2198 14653 2199
rect 14427 2171 14653 2198
rect 14427 2164 14604 2171
rect 14427 2163 14536 2164
rect 14427 2129 14468 2163
rect 14502 2130 14536 2163
rect 14570 2137 14604 2164
rect 14638 2137 14653 2171
rect 14570 2130 14653 2137
rect 14502 2129 14653 2130
rect 14427 2103 14653 2129
rect 14427 2095 14604 2103
rect 14427 2094 14536 2095
rect 14427 2060 14468 2094
rect 14502 2061 14536 2094
rect 14570 2069 14604 2095
rect 14638 2069 14653 2103
rect 14570 2061 14653 2069
rect 14502 2060 14653 2061
rect 14427 2035 14653 2060
rect 14427 2026 14604 2035
rect 14427 2025 14536 2026
rect 14427 1991 14468 2025
rect 14502 1992 14536 2025
rect 14570 2001 14604 2026
rect 14638 2001 14653 2035
rect 14570 1992 14653 2001
rect 14502 1991 14653 1992
rect 14427 1967 14653 1991
rect 14427 1957 14604 1967
rect 14427 1956 14536 1957
rect 14427 1922 14468 1956
rect 14502 1923 14536 1956
rect 14570 1933 14604 1957
rect 14638 1933 14653 1967
rect 14570 1923 14653 1933
rect 14502 1922 14653 1923
rect 14427 1899 14653 1922
rect 14427 1888 14604 1899
rect 14427 1887 14536 1888
rect 14427 1853 14468 1887
rect 14502 1854 14536 1887
rect 14570 1865 14604 1888
rect 14638 1865 14653 1899
rect 14570 1854 14653 1865
rect 14502 1853 14653 1854
rect 14427 1831 14653 1853
rect 14427 1819 14604 1831
rect 14427 1818 14536 1819
rect 14427 1784 14468 1818
rect 14502 1785 14536 1818
rect 14570 1797 14604 1819
rect 14638 1797 14653 1831
rect 14570 1785 14653 1797
rect 14502 1784 14653 1785
rect 14427 1763 14653 1784
rect 14427 1750 14604 1763
rect 14427 1749 14536 1750
rect 14427 1715 14468 1749
rect 14502 1716 14536 1749
rect 14570 1729 14604 1750
rect 14638 1729 14653 1763
rect 14570 1716 14653 1729
rect 14502 1715 14653 1716
rect 14427 1695 14653 1715
rect 14427 1681 14604 1695
rect 14427 1680 14536 1681
rect 14427 1646 14468 1680
rect 14502 1647 14536 1680
rect 14570 1661 14604 1681
rect 14638 1661 14653 1695
rect 14570 1647 14653 1661
rect 14502 1646 14653 1647
rect 14427 1627 14653 1646
rect 14427 1612 14604 1627
rect 14427 1611 14536 1612
rect 14427 1577 14468 1611
rect 14502 1578 14536 1611
rect 14570 1593 14604 1612
rect 14638 1593 14653 1627
rect 14570 1578 14653 1593
rect 14502 1577 14653 1578
rect 14427 1559 14653 1577
rect 14427 1552 14604 1559
rect 482 1551 682 1552
rect 482 1517 497 1551
rect 531 1541 682 1551
rect 531 1517 565 1541
rect 482 1507 565 1517
rect 599 1507 633 1541
rect 667 1507 682 1541
rect 482 1483 682 1507
rect 482 1449 497 1483
rect 531 1472 682 1483
rect 531 1449 565 1472
rect 482 1438 565 1449
rect 599 1438 633 1472
rect 667 1438 682 1472
rect 482 1415 682 1438
rect 482 1381 497 1415
rect 531 1403 682 1415
rect 531 1381 565 1403
rect 482 1369 565 1381
rect 599 1369 633 1403
rect 667 1369 682 1403
rect 14453 1543 14604 1552
rect 14453 1542 14536 1543
rect 14453 1508 14468 1542
rect 14502 1509 14536 1542
rect 14570 1525 14604 1543
rect 14638 1525 14653 1559
rect 14570 1509 14653 1525
rect 14502 1508 14653 1509
rect 14453 1491 14653 1508
rect 14453 1474 14604 1491
rect 14453 1473 14536 1474
rect 14453 1439 14468 1473
rect 14502 1440 14536 1473
rect 14570 1457 14604 1474
rect 14638 1457 14653 1491
rect 14570 1440 14653 1457
rect 14502 1439 14653 1440
rect 14453 1423 14653 1439
rect 14453 1405 14604 1423
rect 14453 1404 14536 1405
rect 482 1347 682 1369
rect 482 1313 497 1347
rect 531 1334 682 1347
rect 531 1313 565 1334
rect 482 1300 565 1313
rect 599 1300 633 1334
rect 667 1300 682 1334
rect 482 1279 682 1300
rect 482 1245 497 1279
rect 531 1265 682 1279
rect 531 1245 565 1265
rect 482 1231 565 1245
rect 599 1231 633 1265
rect 667 1231 682 1265
rect 482 1211 682 1231
rect 482 1177 497 1211
rect 531 1196 682 1211
rect 531 1177 565 1196
rect 482 1162 565 1177
rect 599 1162 633 1196
rect 667 1162 682 1196
rect 482 1143 682 1162
rect 482 1109 497 1143
rect 531 1127 682 1143
rect 531 1109 565 1127
rect 482 1093 565 1109
rect 599 1093 633 1127
rect 667 1093 682 1127
rect 482 1075 682 1093
rect 482 1041 497 1075
rect 531 1058 682 1075
rect 531 1041 565 1058
rect 482 1024 565 1041
rect 599 1024 633 1058
rect 667 1024 682 1058
rect 482 1007 682 1024
rect 482 973 497 1007
rect 531 989 682 1007
rect 531 973 565 989
rect 482 955 565 973
rect 599 955 633 989
rect 667 955 682 989
rect 482 939 682 955
rect 482 769 497 939
rect 531 920 682 939
rect 667 867 682 920
rect 14453 1370 14468 1404
rect 14502 1371 14536 1404
rect 14570 1389 14604 1405
rect 14638 1389 14653 1423
rect 14570 1371 14653 1389
rect 14502 1370 14653 1371
rect 14453 1355 14653 1370
rect 14453 1336 14604 1355
rect 14453 1335 14536 1336
rect 14453 1301 14468 1335
rect 14502 1302 14536 1335
rect 14570 1321 14604 1336
rect 14638 1321 14653 1355
rect 14570 1302 14653 1321
rect 14502 1301 14653 1302
rect 14453 1287 14653 1301
rect 14453 1267 14604 1287
rect 14453 1266 14536 1267
rect 14453 1232 14468 1266
rect 14502 1233 14536 1266
rect 14570 1253 14604 1267
rect 14638 1253 14653 1287
rect 14570 1233 14653 1253
rect 14502 1232 14653 1233
rect 14453 1218 14653 1232
rect 14453 1198 14604 1218
rect 14453 1197 14536 1198
rect 14453 1163 14468 1197
rect 14502 1164 14536 1197
rect 14570 1184 14604 1198
rect 14638 1184 14653 1218
rect 14570 1164 14653 1184
rect 14502 1163 14653 1164
rect 14453 1149 14653 1163
rect 14453 1129 14604 1149
rect 14453 1128 14536 1129
rect 14453 1094 14468 1128
rect 14502 1095 14536 1128
rect 14570 1115 14604 1129
rect 14638 1115 14653 1149
rect 14570 1095 14653 1115
rect 14502 1094 14653 1095
rect 14453 1080 14653 1094
rect 14453 1060 14604 1080
rect 14453 1059 14536 1060
rect 14453 1025 14468 1059
rect 14502 1026 14536 1059
rect 14570 1046 14604 1060
rect 14638 1046 14653 1080
rect 14570 1026 14653 1046
rect 14502 1025 14653 1026
rect 14453 1011 14653 1025
rect 14453 991 14604 1011
rect 14453 990 14536 991
rect 14453 956 14468 990
rect 14502 957 14536 990
rect 14570 977 14604 991
rect 14638 977 14653 1011
rect 14570 957 14653 977
rect 14502 956 14653 957
rect 14453 942 14653 956
rect 14453 922 14604 942
rect 14453 921 14536 922
rect 14453 887 14468 921
rect 14502 888 14536 921
rect 14570 908 14604 922
rect 14638 908 14653 942
rect 14570 888 14653 908
rect 14502 887 14653 888
rect 14453 873 14653 887
rect 14453 867 14604 873
rect 667 853 14604 867
rect 667 852 14536 853
rect 667 818 702 852
rect 736 818 771 852
rect 805 818 840 852
rect 874 818 909 852
rect 943 818 978 852
rect 1012 818 1047 852
rect 1081 818 1116 852
rect 1150 818 1185 852
rect 1219 818 1254 852
rect 1288 818 1323 852
rect 1357 818 1392 852
rect 1426 818 1461 852
rect 1495 818 1530 852
rect 1564 818 1599 852
rect 1633 818 1668 852
rect 1702 818 1737 852
rect 1771 818 1806 852
rect 1840 818 1875 852
rect 1909 818 1944 852
rect 1978 818 2013 852
rect 2047 818 2082 852
rect 2116 818 2151 852
rect 2185 818 2220 852
rect 2254 818 2289 852
rect 2323 818 2358 852
rect 2392 818 2427 852
rect 2461 818 2496 852
rect 2530 818 2565 852
rect 2599 818 2634 852
rect 2668 818 2703 852
rect 2737 818 2772 852
rect 599 784 2772 818
rect 14502 819 14536 852
rect 14570 839 14604 853
rect 14638 839 14653 873
rect 14570 819 14653 839
rect 14502 804 14653 819
rect 14502 784 14604 804
rect 482 750 565 769
rect 599 750 634 784
rect 668 750 703 784
rect 737 750 772 784
rect 806 750 841 784
rect 875 750 910 784
rect 944 750 979 784
rect 1013 750 1048 784
rect 1082 750 1117 784
rect 1151 750 1186 784
rect 1220 750 1255 784
rect 1289 750 1324 784
rect 1358 750 1393 784
rect 1427 750 1462 784
rect 1496 750 1531 784
rect 1565 750 1600 784
rect 1634 750 1669 784
rect 1703 750 1738 784
rect 1772 750 1807 784
rect 1841 750 1876 784
rect 1910 750 1945 784
rect 1979 750 2014 784
rect 2048 750 2083 784
rect 2117 750 2152 784
rect 2186 750 2221 784
rect 2255 750 2290 784
rect 2324 750 2359 784
rect 2393 750 2428 784
rect 2462 750 2497 784
rect 2531 750 2566 784
rect 2600 750 2635 784
rect 2669 750 2704 784
rect 2738 750 2772 784
rect 14570 770 14604 784
rect 14638 770 14653 804
rect 14570 750 14653 770
rect 482 716 4725 750
rect 482 682 516 716
rect 550 682 585 716
rect 619 682 654 716
rect 688 682 723 716
rect 757 682 792 716
rect 826 682 861 716
rect 895 682 930 716
rect 964 682 999 716
rect 1033 682 1068 716
rect 1102 682 1137 716
rect 1171 682 1206 716
rect 1240 682 1275 716
rect 1309 682 1344 716
rect 1378 682 1413 716
rect 1447 682 1482 716
rect 1516 682 1551 716
rect 1585 682 1620 716
rect 1654 682 1689 716
rect 1723 682 1758 716
rect 1792 682 1827 716
rect 1861 682 1896 716
rect 1930 682 1965 716
rect 1999 682 2034 716
rect 2068 682 2103 716
rect 2137 682 2172 716
rect 2206 682 2241 716
rect 2275 682 2310 716
rect 2344 682 2379 716
rect 2413 682 2448 716
rect 2482 682 2517 716
rect 2551 682 2586 716
rect 2620 682 2655 716
rect 2689 682 2724 716
rect 2758 682 2793 716
rect 2827 682 2862 716
rect 2896 682 2931 716
rect 2965 682 3000 716
rect 3034 682 3069 716
rect 3103 682 3138 716
rect 3172 682 3207 716
rect 3241 682 3276 716
rect 3310 682 3345 716
rect 3379 682 3414 716
rect 3448 682 3483 716
rect 3517 682 3552 716
rect 3586 682 3621 716
rect 3655 682 3690 716
rect 3724 682 3759 716
rect 3793 682 3828 716
rect 3862 682 3897 716
rect 3931 682 3966 716
rect 4000 682 4035 716
rect 4069 682 4104 716
rect 4138 682 4173 716
rect 4207 682 4242 716
rect 4276 682 4311 716
rect 4345 682 4380 716
rect 4414 682 4449 716
rect 4483 682 4518 716
rect 4552 682 4587 716
rect 4621 682 4656 716
rect 4690 682 4725 716
rect 14551 735 14653 750
rect 14551 701 14604 735
rect 14638 701 14653 735
rect 14551 682 14653 701
rect 482 667 14653 682
<< mvpsubdiffcont >>
rect 252 5048 286 5082
rect 320 5048 354 5082
rect 388 5048 422 5082
rect 456 5048 490 5082
rect 524 5048 558 5082
rect 592 5048 626 5082
rect 660 5048 694 5082
rect 728 5048 762 5082
rect 796 5048 830 5082
rect 864 5048 898 5082
rect 932 5048 966 5082
rect 1000 5048 1034 5082
rect 1068 5048 1102 5082
rect 1136 5048 1170 5082
rect 1204 5048 1238 5082
rect 1272 5048 1306 5082
rect 1340 5048 1374 5082
rect 1408 5048 1442 5082
rect 1476 5048 1510 5082
rect 1544 5048 1578 5082
rect 1612 5048 1646 5082
rect 1680 5048 1714 5082
rect 1748 5048 1782 5082
rect 1816 5048 1850 5082
rect 1884 5048 1918 5082
rect 1952 5048 1986 5082
rect 2020 5048 2054 5082
rect 2088 5048 2122 5082
rect 2156 5048 2190 5082
rect 2224 5048 2258 5082
rect 2292 5048 2326 5082
rect 2360 5048 2394 5082
rect 2428 5048 2462 5082
rect 2496 5048 2530 5082
rect 2564 5048 2598 5082
rect 2632 5048 2666 5082
rect 2700 5048 2734 5082
rect 2768 5048 2802 5082
rect 2836 5048 2870 5082
rect 2904 5048 2938 5082
rect 2972 5048 3006 5082
rect 3040 5048 3074 5082
rect 3108 5048 3142 5082
rect 3176 5048 3210 5082
rect 3244 5048 3278 5082
rect 3312 5048 3346 5082
rect 3380 5048 3414 5082
rect 3448 5048 3482 5082
rect 3516 5048 3550 5082
rect 3584 5048 3618 5082
rect 3652 5048 3686 5082
rect 3720 5048 3754 5082
rect 3788 5048 3822 5082
rect 3856 5048 3890 5082
rect 3924 5048 3958 5082
rect 3992 5048 4026 5082
rect 4060 5048 4094 5082
rect 4128 5048 4162 5082
rect 4196 5048 4230 5082
rect 4264 5048 4298 5082
rect 4332 5048 4366 5082
rect 4400 5048 4434 5082
rect 4468 5048 4502 5082
rect 4536 5048 4570 5082
rect 4604 5048 4638 5082
rect 4672 5048 4706 5082
rect 4740 5048 4774 5082
rect 4808 5048 4842 5082
rect 4876 5048 4910 5082
rect 4944 5048 4978 5082
rect 5012 5048 5046 5082
rect 5080 5048 5114 5082
rect 5148 5048 5182 5082
rect 5216 5048 5250 5082
rect 5284 5048 5318 5082
rect 5352 5048 5386 5082
rect 5420 5048 5454 5082
rect 5488 5048 5522 5082
rect 5556 5048 5590 5082
rect 5624 5048 5658 5082
rect 5692 5048 5726 5082
rect 5760 5048 5794 5082
rect 5828 5048 5862 5082
rect 5896 5048 5930 5082
rect 5964 5048 5998 5082
rect 6032 5048 6066 5082
rect 6100 5048 6134 5082
rect 6168 5048 6202 5082
rect 6236 5048 6270 5082
rect 6304 5048 6338 5082
rect 6372 5048 6406 5082
rect 6440 5048 6474 5082
rect 6508 5048 6542 5082
rect 6576 5048 6610 5082
rect 6644 5048 6678 5082
rect 6712 5048 6746 5082
rect 6780 5048 6814 5082
rect 6848 5048 6882 5082
rect 6916 5048 6950 5082
rect 6984 5048 7018 5082
rect 7052 5048 7086 5082
rect 7120 5048 7154 5082
rect 7188 5048 7222 5082
rect 7256 5048 7290 5082
rect 7324 5048 7358 5082
rect 7392 5048 7426 5082
rect 7460 5048 7494 5082
rect 7528 5048 7562 5082
rect 7596 5048 7630 5082
rect 7664 5048 7698 5082
rect 7732 5048 7766 5082
rect 7800 5048 7834 5082
rect 7868 5048 7902 5082
rect 7936 5048 7970 5082
rect 8004 5048 8038 5082
rect 8072 5048 8106 5082
rect 8140 5048 8174 5082
rect 8208 5048 8242 5082
rect 8276 5048 8310 5082
rect 8344 5048 8378 5082
rect 8412 5048 8446 5082
rect 8480 5048 8514 5082
rect 8548 5048 8582 5082
rect 8616 5048 8650 5082
rect 8684 5048 8718 5082
rect 8752 5048 8786 5082
rect 8820 5048 8854 5082
rect 8888 5048 8922 5082
rect 8956 5048 8990 5082
rect 9024 5048 9058 5082
rect 9092 5048 9126 5082
rect 9160 5048 9194 5082
rect 9228 5048 9262 5082
rect 9296 5048 9330 5082
rect 9364 5048 9398 5082
rect 9432 5048 9466 5082
rect 9500 5048 9534 5082
rect 9568 5048 9602 5082
rect 9636 5048 9670 5082
rect 9704 5048 9738 5082
rect 9772 5048 9806 5082
rect 9840 5048 9874 5082
rect 9908 5048 9942 5082
rect 9976 5048 10010 5082
rect 10044 5048 10078 5082
rect 10112 5048 10146 5082
rect 10180 5048 10214 5082
rect 10248 5048 10282 5082
rect 10316 5048 10350 5082
rect 10384 5048 10418 5082
rect 10452 5048 10486 5082
rect 10520 5048 10554 5082
rect 10588 5048 10622 5082
rect 10656 5048 10690 5082
rect 10724 5048 10758 5082
rect 10792 5048 10826 5082
rect 10860 5048 10894 5082
rect 10928 5048 10962 5082
rect 10996 5048 11030 5082
rect 11064 5048 11098 5082
rect 11132 5048 11166 5082
rect 11200 5048 11234 5082
rect 11268 5048 11302 5082
rect 11336 5048 11370 5082
rect 11404 5048 11438 5082
rect 11472 5048 11506 5082
rect 11540 5048 11574 5082
rect 11608 5048 11642 5082
rect 11676 5048 11710 5082
rect 11744 5048 11778 5082
rect 11812 5048 11846 5082
rect 11880 5048 11914 5082
rect 11948 5048 11982 5082
rect 12016 5048 12050 5082
rect 12084 5048 12118 5082
rect 12152 5048 12186 5082
rect 12220 5048 12254 5082
rect 12288 5048 12322 5082
rect 12356 5048 12390 5082
rect 12424 5048 12458 5082
rect 12492 5048 12526 5082
rect 12560 5048 12594 5082
rect 12628 5048 12662 5082
rect 12696 5048 12730 5082
rect 12764 5048 12798 5082
rect 12832 5048 12866 5082
rect 12900 5048 12934 5082
rect 12968 5048 13002 5082
rect 13036 5048 13070 5082
rect 13104 5048 13138 5082
rect 13172 5048 13206 5082
rect 13240 5048 13274 5082
rect 13308 5048 13342 5082
rect 13376 5048 13410 5082
rect 13444 5048 13478 5082
rect 13512 5048 13546 5082
rect 13580 5048 13614 5082
rect 13648 5048 13682 5082
rect 13716 5048 13750 5082
rect 13784 5048 13818 5082
rect 13852 5048 13886 5082
rect 13920 5048 13954 5082
rect 13988 5048 14022 5082
rect 14056 5048 14090 5082
rect 14124 5048 14158 5082
rect 14192 5048 14226 5082
rect 14260 5048 14294 5082
rect 14328 5048 14362 5082
rect 14396 5048 14430 5082
rect 14464 5048 14498 5082
rect 14532 5048 14566 5082
rect 14600 5048 14634 5082
rect 14668 5048 14702 5082
rect 14736 5048 14770 5082
rect 14804 5048 14838 5082
rect 14872 5048 14906 5082
rect 252 4966 286 5000
rect 320 4966 354 5000
rect 388 4966 422 5000
rect 456 4966 490 5000
rect 524 4966 558 5000
rect 592 4966 626 5000
rect 660 4966 694 5000
rect 728 4966 762 5000
rect 796 4966 830 5000
rect 864 4966 898 5000
rect 932 4966 966 5000
rect 1000 4966 1034 5000
rect 1068 4966 1102 5000
rect 1136 4966 1170 5000
rect 1204 4966 1238 5000
rect 1272 4966 1306 5000
rect 1340 4966 1374 5000
rect 1408 4966 1442 5000
rect 1476 4966 1510 5000
rect 1544 4966 1578 5000
rect 1612 4966 1646 5000
rect 1680 4966 1714 5000
rect 1748 4966 1782 5000
rect 1816 4966 1850 5000
rect 1884 4966 1918 5000
rect 1952 4966 1986 5000
rect 2020 4966 2054 5000
rect 2088 4966 2122 5000
rect 2156 4966 2190 5000
rect 2224 4966 2258 5000
rect 2292 4966 2326 5000
rect 2360 4966 2394 5000
rect 2428 4966 2462 5000
rect 2496 4966 2530 5000
rect 2564 4966 2598 5000
rect 2632 4966 2666 5000
rect 2700 4966 2734 5000
rect 2768 4966 2802 5000
rect 2836 4966 2870 5000
rect 2904 4966 2938 5000
rect 2972 4966 3006 5000
rect 3040 4966 3074 5000
rect 3108 4966 3142 5000
rect 3176 4966 3210 5000
rect 3244 4966 3278 5000
rect 3312 4966 3346 5000
rect 3380 4966 3414 5000
rect 3448 4966 3482 5000
rect 3516 4966 3550 5000
rect 3584 4966 3618 5000
rect 3652 4966 3686 5000
rect 3720 4966 3754 5000
rect 3788 4966 3822 5000
rect 3856 4966 3890 5000
rect 3924 4966 3958 5000
rect 3992 4966 4026 5000
rect 4060 4966 4094 5000
rect 4128 4966 4162 5000
rect 4196 4966 4230 5000
rect 4264 4966 4298 5000
rect 4332 4966 4366 5000
rect 4400 4966 4434 5000
rect 4468 4966 4502 5000
rect 4536 4966 4570 5000
rect 4604 4966 4638 5000
rect 4672 4966 4706 5000
rect 4740 4966 4774 5000
rect 4808 4966 4842 5000
rect 4876 4966 4910 5000
rect 4944 4966 4978 5000
rect 5012 4966 5046 5000
rect 5080 4966 5114 5000
rect 5148 4966 5182 5000
rect 5216 4966 5250 5000
rect 5284 4966 5318 5000
rect 5352 4966 5386 5000
rect 5420 4966 5454 5000
rect 5488 4966 5522 5000
rect 5556 4966 5590 5000
rect 5624 4966 5658 5000
rect 5692 4966 5726 5000
rect 5760 4966 5794 5000
rect 5828 4966 5862 5000
rect 5896 4966 5930 5000
rect 5964 4966 5998 5000
rect 6032 4966 6066 5000
rect 6100 4966 6134 5000
rect 6168 4966 6202 5000
rect 6236 4966 6270 5000
rect 6304 4966 6338 5000
rect 6372 4966 6406 5000
rect 6440 4966 6474 5000
rect 6508 4966 6542 5000
rect 6576 4966 6610 5000
rect 6644 4966 6678 5000
rect 6712 4966 6746 5000
rect 6780 4966 6814 5000
rect 6848 4966 6882 5000
rect 6916 4966 6950 5000
rect 6984 4966 7018 5000
rect 7052 4966 7086 5000
rect 7120 4966 7154 5000
rect 7188 4966 7222 5000
rect 7256 4966 7290 5000
rect 7324 4966 7358 5000
rect 7392 4966 7426 5000
rect 7460 4966 7494 5000
rect 7528 4966 7562 5000
rect 7596 4966 7630 5000
rect 7664 4966 7698 5000
rect 7732 4966 7766 5000
rect 7800 4966 7834 5000
rect 7868 4966 7902 5000
rect 7936 4966 7970 5000
rect 8004 4966 8038 5000
rect 8072 4966 8106 5000
rect 8140 4966 8174 5000
rect 8208 4966 8242 5000
rect 8276 4966 8310 5000
rect 8344 4966 8378 5000
rect 8412 4966 8446 5000
rect 8480 4966 8514 5000
rect 8548 4966 8582 5000
rect 8616 4966 8650 5000
rect 8684 4966 8718 5000
rect 8752 4966 8786 5000
rect 8820 4966 8854 5000
rect 8888 4966 8922 5000
rect 8956 4966 8990 5000
rect 9024 4966 9058 5000
rect 9092 4966 9126 5000
rect 9160 4966 9194 5000
rect 9228 4966 9262 5000
rect 9296 4966 9330 5000
rect 9364 4966 9398 5000
rect 9432 4966 9466 5000
rect 9500 4966 9534 5000
rect 9568 4966 9602 5000
rect 9636 4966 9670 5000
rect 9704 4966 9738 5000
rect 9772 4966 9806 5000
rect 9840 4966 9874 5000
rect 9908 4966 9942 5000
rect 9976 4966 10010 5000
rect 10044 4966 10078 5000
rect 10112 4966 10146 5000
rect 10180 4966 10214 5000
rect 10248 4966 10282 5000
rect 10316 4966 10350 5000
rect 10384 4966 10418 5000
rect 10452 4966 10486 5000
rect 10520 4966 10554 5000
rect 10588 4966 10622 5000
rect 10656 4966 10690 5000
rect 10724 4966 10758 5000
rect 10792 4966 10826 5000
rect 10860 4966 10894 5000
rect 10928 4966 10962 5000
rect 10996 4966 11030 5000
rect 11064 4966 11098 5000
rect 11132 4966 11166 5000
rect 11200 4966 11234 5000
rect 11268 4966 11302 5000
rect 11336 4966 11370 5000
rect 11404 4966 11438 5000
rect 11472 4966 11506 5000
rect 11540 4966 11574 5000
rect 11608 4966 11642 5000
rect 11676 4966 11710 5000
rect 11744 4966 11778 5000
rect 11812 4966 11846 5000
rect 11880 4966 11914 5000
rect 11948 4966 11982 5000
rect 12016 4966 12050 5000
rect 12084 4966 12118 5000
rect 12152 4966 12186 5000
rect 12220 4966 12254 5000
rect 12288 4966 12322 5000
rect 12356 4966 12390 5000
rect 12424 4966 12458 5000
rect 12492 4966 12526 5000
rect 12560 4966 12594 5000
rect 12628 4966 12662 5000
rect 12696 4966 12730 5000
rect 12764 4966 12798 5000
rect 12832 4966 12866 5000
rect 12900 4966 12934 5000
rect 12968 4966 13002 5000
rect 13036 4966 13070 5000
rect 13104 4966 13138 5000
rect 13172 4966 13206 5000
rect 13240 4966 13274 5000
rect 13308 4966 13342 5000
rect 13376 4966 13410 5000
rect 13444 4966 13478 5000
rect 13512 4966 13546 5000
rect 13580 4966 13614 5000
rect 13648 4966 13682 5000
rect 13716 4966 13750 5000
rect 13784 4966 13818 5000
rect 13852 4966 13886 5000
rect 13920 4966 13954 5000
rect 13988 4966 14022 5000
rect 14056 4966 14090 5000
rect 14124 4966 14158 5000
rect 14192 4966 14226 5000
rect 14260 4966 14294 5000
rect 14328 4966 14362 5000
rect 14396 4966 14430 5000
rect 14464 4966 14498 5000
rect 14532 4966 14566 5000
rect 14600 4966 14634 5000
rect 14668 4966 14702 5000
rect 14736 4966 14770 5000
rect 14804 4966 14838 5000
rect 14872 4966 14906 5000
rect 252 4884 286 4918
rect 320 4884 354 4918
rect 388 4884 422 4918
rect 456 4884 490 4918
rect 524 4884 558 4918
rect 592 4884 626 4918
rect 660 4884 694 4918
rect 728 4884 762 4918
rect 796 4884 830 4918
rect 864 4884 898 4918
rect 932 4884 966 4918
rect 1000 4884 1034 4918
rect 1068 4884 1102 4918
rect 1136 4884 1170 4918
rect 1204 4884 1238 4918
rect 1272 4884 1306 4918
rect 1340 4884 1374 4918
rect 1408 4884 1442 4918
rect 1476 4884 1510 4918
rect 1544 4884 1578 4918
rect 1612 4884 1646 4918
rect 1680 4884 1714 4918
rect 1748 4884 1782 4918
rect 1816 4884 1850 4918
rect 1884 4884 1918 4918
rect 1952 4884 1986 4918
rect 2020 4884 2054 4918
rect 2088 4884 2122 4918
rect 2156 4884 2190 4918
rect 2224 4884 2258 4918
rect 2292 4884 2326 4918
rect 2360 4884 2394 4918
rect 2428 4884 2462 4918
rect 2496 4884 2530 4918
rect 2564 4884 2598 4918
rect 2632 4884 2666 4918
rect 2700 4884 2734 4918
rect 2768 4884 2802 4918
rect 2836 4884 2870 4918
rect 2904 4884 2938 4918
rect 2972 4884 3006 4918
rect 3040 4884 3074 4918
rect 3108 4884 3142 4918
rect 3176 4884 3210 4918
rect 3244 4884 3278 4918
rect 3312 4884 3346 4918
rect 3380 4884 3414 4918
rect 3448 4884 3482 4918
rect 3516 4884 3550 4918
rect 3584 4884 3618 4918
rect 3652 4884 3686 4918
rect 3720 4884 3754 4918
rect 3788 4884 3822 4918
rect 3856 4884 3890 4918
rect 3924 4884 3958 4918
rect 3992 4884 4026 4918
rect 4060 4884 4094 4918
rect 4128 4884 4162 4918
rect 4196 4884 4230 4918
rect 4264 4884 4298 4918
rect 4332 4884 4366 4918
rect 4400 4884 4434 4918
rect 4468 4884 4502 4918
rect 4536 4884 4570 4918
rect 4604 4884 4638 4918
rect 4672 4884 4706 4918
rect 4740 4884 4774 4918
rect 4808 4884 4842 4918
rect 4876 4884 4910 4918
rect 4944 4884 4978 4918
rect 5012 4884 5046 4918
rect 5080 4884 5114 4918
rect 5148 4884 5182 4918
rect 5216 4884 5250 4918
rect 5284 4884 5318 4918
rect 5352 4884 5386 4918
rect 5420 4884 5454 4918
rect 5488 4884 5522 4918
rect 5556 4884 5590 4918
rect 5624 4884 5658 4918
rect 5692 4884 5726 4918
rect 5760 4884 5794 4918
rect 5828 4884 5862 4918
rect 5896 4884 5930 4918
rect 5964 4884 5998 4918
rect 6032 4884 6066 4918
rect 6100 4884 6134 4918
rect 6168 4884 6202 4918
rect 6236 4884 6270 4918
rect 6304 4884 6338 4918
rect 6372 4884 6406 4918
rect 6440 4884 6474 4918
rect 6508 4884 6542 4918
rect 6576 4884 6610 4918
rect 6644 4884 6678 4918
rect 6712 4884 6746 4918
rect 6780 4884 6814 4918
rect 6848 4884 6882 4918
rect 6916 4884 6950 4918
rect 6984 4884 7018 4918
rect 7052 4884 7086 4918
rect 7120 4884 7154 4918
rect 7188 4884 7222 4918
rect 7256 4884 7290 4918
rect 7324 4884 7358 4918
rect 7392 4884 7426 4918
rect 7460 4884 7494 4918
rect 7528 4884 7562 4918
rect 7596 4884 7630 4918
rect 7664 4884 7698 4918
rect 7732 4884 7766 4918
rect 7800 4884 7834 4918
rect 7868 4884 7902 4918
rect 7936 4884 7970 4918
rect 8004 4884 8038 4918
rect 8072 4884 8106 4918
rect 8140 4884 8174 4918
rect 8208 4884 8242 4918
rect 8276 4884 8310 4918
rect 8344 4884 8378 4918
rect 8412 4884 8446 4918
rect 8480 4884 8514 4918
rect 8548 4884 8582 4918
rect 8616 4884 8650 4918
rect 8684 4884 8718 4918
rect 8752 4884 8786 4918
rect 8820 4884 8854 4918
rect 8888 4884 8922 4918
rect 8956 4884 8990 4918
rect 9024 4884 9058 4918
rect 9092 4884 9126 4918
rect 9160 4884 9194 4918
rect 9228 4884 9262 4918
rect 9296 4884 9330 4918
rect 9364 4884 9398 4918
rect 9432 4884 9466 4918
rect 9500 4884 9534 4918
rect 9568 4884 9602 4918
rect 9636 4884 9670 4918
rect 9704 4884 9738 4918
rect 9772 4884 9806 4918
rect 9840 4884 9874 4918
rect 9908 4884 9942 4918
rect 9976 4884 10010 4918
rect 10044 4884 10078 4918
rect 10112 4884 10146 4918
rect 10180 4884 10214 4918
rect 10248 4884 10282 4918
rect 10316 4884 10350 4918
rect 10384 4884 10418 4918
rect 10452 4884 10486 4918
rect 10520 4884 10554 4918
rect 10588 4884 10622 4918
rect 10656 4884 10690 4918
rect 10724 4884 10758 4918
rect 10792 4884 10826 4918
rect 10860 4884 10894 4918
rect 10928 4884 10962 4918
rect 10996 4884 11030 4918
rect 11064 4884 11098 4918
rect 11132 4884 11166 4918
rect 11200 4884 11234 4918
rect 11268 4884 11302 4918
rect 11336 4884 11370 4918
rect 11404 4884 11438 4918
rect 11472 4884 11506 4918
rect 11540 4884 11574 4918
rect 11608 4884 11642 4918
rect 11676 4884 11710 4918
rect 11744 4884 11778 4918
rect 11812 4884 11846 4918
rect 11880 4884 11914 4918
rect 11948 4884 11982 4918
rect 12016 4884 12050 4918
rect 12084 4884 12118 4918
rect 12152 4884 12186 4918
rect 12220 4884 12254 4918
rect 12288 4884 12322 4918
rect 12356 4884 12390 4918
rect 12424 4884 12458 4918
rect 12492 4884 12526 4918
rect 12560 4884 12594 4918
rect 12628 4884 12662 4918
rect 12696 4884 12730 4918
rect 12764 4884 12798 4918
rect 12832 4884 12866 4918
rect 12900 4884 12934 4918
rect 12968 4884 13002 4918
rect 13036 4884 13070 4918
rect 13104 4884 13138 4918
rect 13172 4884 13206 4918
rect 13240 4884 13274 4918
rect 13308 4884 13342 4918
rect 13376 4884 13410 4918
rect 13444 4884 13478 4918
rect 13512 4884 13546 4918
rect 13580 4884 13614 4918
rect 13648 4884 13682 4918
rect 13716 4884 13750 4918
rect 13784 4884 13818 4918
rect 13852 4884 13886 4918
rect 13920 4884 13954 4918
rect 13988 4884 14022 4918
rect 14056 4884 14090 4918
rect 14124 4884 14158 4918
rect 14192 4884 14226 4918
rect 14260 4884 14294 4918
rect 14328 4884 14362 4918
rect 14396 4884 14430 4918
rect 14464 4884 14498 4918
rect 14532 4884 14566 4918
rect 14600 4884 14634 4918
rect 14668 4884 14702 4918
rect 14736 4884 14770 4918
rect 14804 4884 14838 4918
rect 14872 4884 14906 4918
rect 193 599 295 4849
rect 14806 4815 14840 4849
rect 14906 4815 14940 4849
rect 14806 4747 14840 4781
rect 14906 4747 14940 4781
rect 14806 4679 14840 4713
rect 14906 4679 14940 4713
rect 14806 4611 14840 4645
rect 14906 4611 14940 4645
rect 14806 4543 14840 4577
rect 14906 4543 14940 4577
rect 14806 4475 14840 4509
rect 14906 4475 14940 4509
rect 14806 4407 14840 4441
rect 14906 4407 14940 4441
rect 14806 4339 14840 4373
rect 14906 4339 14940 4373
rect 14806 4271 14840 4305
rect 14906 4271 14940 4305
rect 14806 4203 14840 4237
rect 14906 4203 14940 4237
rect 14806 4135 14840 4169
rect 14906 4135 14940 4169
rect 14806 4067 14840 4101
rect 14906 4067 14940 4101
rect 14806 3999 14840 4033
rect 14906 3999 14940 4033
rect 14806 3931 14840 3965
rect 14906 3931 14940 3965
rect 14806 3863 14840 3897
rect 14906 3863 14940 3897
rect 14806 3795 14840 3829
rect 14906 3795 14940 3829
rect 14806 3727 14840 3761
rect 14906 3727 14940 3761
rect 14806 3659 14840 3693
rect 14906 3659 14940 3693
rect 14806 3591 14840 3625
rect 14906 3591 14940 3625
rect 14806 3523 14840 3557
rect 14906 3523 14940 3557
rect 14806 3455 14840 3489
rect 14906 3455 14940 3489
rect 14806 3387 14840 3421
rect 14906 3387 14940 3421
rect 14806 3319 14840 3353
rect 14906 3319 14940 3353
rect 14806 3251 14840 3285
rect 14906 3251 14940 3285
rect 14806 3183 14840 3217
rect 14906 3183 14940 3217
rect 14806 3115 14840 3149
rect 14906 3115 14940 3149
rect 14806 3047 14840 3081
rect 14906 3047 14940 3081
rect 14806 2979 14840 3013
rect 14906 2979 14940 3013
rect 14806 2911 14840 2945
rect 14906 2911 14940 2945
rect 14806 2843 14840 2877
rect 14906 2843 14940 2877
rect 14806 2775 14840 2809
rect 14906 2775 14940 2809
rect 14806 2707 14840 2741
rect 14906 2707 14940 2741
rect 14806 2639 14840 2673
rect 14906 2639 14940 2673
rect 14806 2571 14840 2605
rect 14906 2571 14940 2605
rect 14806 2503 14840 2537
rect 14906 2503 14940 2537
rect 14806 2435 14840 2469
rect 14906 2435 14940 2469
rect 14806 2367 14840 2401
rect 14906 2367 14940 2401
rect 14806 2299 14840 2333
rect 14906 2299 14940 2333
rect 14806 2231 14840 2265
rect 14906 2231 14940 2265
rect 14806 2163 14840 2197
rect 14906 2163 14940 2197
rect 14806 2095 14840 2129
rect 14906 2095 14940 2129
rect 14806 2027 14840 2061
rect 14906 2027 14940 2061
rect 14806 1959 14840 1993
rect 14906 1959 14940 1993
rect 14806 1891 14840 1925
rect 14906 1891 14940 1925
rect 14806 1823 14840 1857
rect 14906 1823 14940 1857
rect 14806 1755 14840 1789
rect 14906 1755 14940 1789
rect 14806 1687 14840 1721
rect 14906 1687 14940 1721
rect 14806 1619 14840 1653
rect 14906 1619 14940 1653
rect 14806 1551 14840 1585
rect 14906 1551 14940 1585
rect 14806 1483 14840 1517
rect 14906 1483 14940 1517
rect 14806 1415 14840 1449
rect 14906 1415 14940 1449
rect 14806 1347 14840 1381
rect 14906 1347 14940 1381
rect 14806 1279 14840 1313
rect 14906 1279 14940 1313
rect 14806 1211 14840 1245
rect 14906 1211 14940 1245
rect 14806 1143 14840 1177
rect 14906 1143 14940 1177
rect 14806 1075 14840 1109
rect 14906 1075 14940 1109
rect 14806 1007 14840 1041
rect 14906 1007 14940 1041
rect 14806 939 14840 973
rect 14906 939 14940 973
rect 14806 871 14840 905
rect 14906 871 14940 905
rect 14806 803 14840 837
rect 14906 803 14940 837
rect 14806 735 14840 769
rect 14906 735 14940 769
rect 14806 667 14840 701
rect 14906 667 14940 701
rect 14806 599 14840 633
rect 14906 599 14940 633
rect 193 407 14847 509
<< mvnsubdiffcont >>
rect 497 4585 531 4619
rect 584 4570 10410 4638
rect 10445 4604 10479 4638
rect 10514 4604 10548 4638
rect 10583 4604 10617 4638
rect 10652 4604 10686 4638
rect 10721 4604 10755 4638
rect 10790 4604 10824 4638
rect 10859 4604 10893 4638
rect 10928 4604 10962 4638
rect 10997 4604 11031 4638
rect 11066 4604 11100 4638
rect 11135 4604 11169 4638
rect 11204 4604 11238 4638
rect 11273 4604 11307 4638
rect 11342 4604 11376 4638
rect 11411 4604 11445 4638
rect 11480 4604 11514 4638
rect 11549 4604 11583 4638
rect 11618 4604 11652 4638
rect 11687 4604 11721 4638
rect 11756 4604 11790 4638
rect 11825 4604 11859 4638
rect 11894 4604 11928 4638
rect 11963 4604 11997 4638
rect 12032 4604 12066 4638
rect 12101 4604 12135 4638
rect 12170 4604 12204 4638
rect 12239 4604 12273 4638
rect 12308 4604 12342 4638
rect 12377 4604 12411 4638
rect 12446 4604 12480 4638
rect 12515 4604 12549 4638
rect 12584 4604 12618 4638
rect 12653 4604 12687 4638
rect 12722 4604 12756 4638
rect 12791 4604 12825 4638
rect 12860 4604 12894 4638
rect 12929 4604 12963 4638
rect 12998 4604 13032 4638
rect 13067 4604 13101 4638
rect 13136 4604 13170 4638
rect 13205 4604 13239 4638
rect 13274 4604 13308 4638
rect 13343 4604 13377 4638
rect 13412 4604 13446 4638
rect 13481 4604 13515 4638
rect 13550 4604 13584 4638
rect 13619 4604 13653 4638
rect 13688 4604 13722 4638
rect 13757 4604 13791 4638
rect 13826 4604 13860 4638
rect 13895 4604 13929 4638
rect 13964 4604 13998 4638
rect 14033 4604 14067 4638
rect 14102 4604 14136 4638
rect 14171 4604 14205 4638
rect 14240 4604 14274 4638
rect 14309 4604 14343 4638
rect 14378 4604 14412 4638
rect 14447 4604 14481 4638
rect 14516 4604 14550 4638
rect 14585 4604 14619 4638
rect 497 4515 531 4549
rect 565 4536 12363 4570
rect 12397 4536 12431 4570
rect 12466 4536 12500 4570
rect 12535 4536 12569 4570
rect 12604 4536 12638 4570
rect 12673 4536 12707 4570
rect 12742 4536 12776 4570
rect 12811 4536 12845 4570
rect 12880 4536 12914 4570
rect 12949 4536 12983 4570
rect 13018 4536 13052 4570
rect 13087 4536 13121 4570
rect 13156 4536 13190 4570
rect 13225 4536 13259 4570
rect 13294 4536 13328 4570
rect 13363 4536 13397 4570
rect 13432 4536 13466 4570
rect 13501 4536 13535 4570
rect 13570 4536 13604 4570
rect 13639 4536 13673 4570
rect 13708 4536 13742 4570
rect 13777 4536 13811 4570
rect 13846 4536 13880 4570
rect 13915 4536 13949 4570
rect 13984 4536 14018 4570
rect 14053 4536 14087 4570
rect 14122 4536 14156 4570
rect 14191 4536 14225 4570
rect 14260 4536 14294 4570
rect 14329 4536 14363 4570
rect 14398 4536 14432 4570
rect 14467 4536 14501 4570
rect 14536 4551 14570 4570
rect 497 4445 531 4479
rect 565 4464 599 4498
rect 633 4468 12363 4536
rect 14536 4502 14638 4551
rect 12398 4468 12432 4502
rect 12467 4468 12501 4502
rect 12536 4468 12570 4502
rect 12605 4468 12639 4502
rect 12674 4468 12708 4502
rect 12743 4468 12777 4502
rect 12812 4468 12846 4502
rect 12881 4468 12915 4502
rect 12950 4468 12984 4502
rect 13019 4468 13053 4502
rect 13088 4468 13122 4502
rect 13157 4468 13191 4502
rect 13226 4468 13260 4502
rect 13295 4468 13329 4502
rect 13364 4468 13398 4502
rect 13433 4468 13467 4502
rect 13502 4468 13536 4502
rect 13571 4468 13605 4502
rect 13640 4468 13674 4502
rect 13709 4468 13743 4502
rect 13778 4468 13812 4502
rect 13847 4468 13881 4502
rect 13916 4468 13950 4502
rect 13985 4468 14019 4502
rect 14054 4468 14088 4502
rect 14123 4468 14157 4502
rect 14192 4468 14226 4502
rect 14261 4468 14295 4502
rect 14330 4468 14364 4502
rect 14399 4468 14433 4502
rect 497 4375 531 4409
rect 565 4392 599 4426
rect 633 4395 667 4429
rect 497 4305 531 4339
rect 565 4320 599 4354
rect 633 4322 667 4356
rect 497 4235 531 4269
rect 565 4248 599 4282
rect 633 4249 667 4283
rect 497 4165 531 4199
rect 565 4176 599 4210
rect 633 4177 667 4211
rect 497 4095 531 4129
rect 565 4104 599 4138
rect 633 4105 667 4139
rect 497 4025 531 4059
rect 565 4032 599 4066
rect 633 4033 667 4067
rect 497 3955 531 3989
rect 565 3960 599 3994
rect 633 3961 667 3995
rect 497 3886 531 3920
rect 565 3888 599 3922
rect 633 3889 667 3923
rect 497 3817 531 3851
rect 565 3817 599 3851
rect 633 3817 667 3851
rect 497 3715 531 3749
rect 565 3715 599 3749
rect 633 3715 667 3749
rect 497 3646 531 3680
rect 565 3646 599 3680
rect 633 3646 667 3680
rect 497 3577 531 3611
rect 565 3577 599 3611
rect 633 3577 667 3611
rect 497 3508 531 3542
rect 565 3508 599 3542
rect 633 3508 667 3542
rect 497 3439 531 3473
rect 565 3439 599 3473
rect 633 3439 667 3473
rect 497 3370 531 3404
rect 565 3370 599 3404
rect 633 3370 667 3404
rect 497 3301 531 3335
rect 565 3301 599 3335
rect 633 3301 667 3335
rect 497 3232 531 3266
rect 565 3232 599 3266
rect 633 3232 667 3266
rect 497 3163 531 3197
rect 565 3163 599 3197
rect 633 3163 667 3197
rect 1635 4048 1669 4082
rect 1635 3980 1669 4014
rect 1635 3912 1669 3946
rect 1635 3844 1669 3878
rect 1635 3776 1669 3810
rect 1635 3708 1669 3742
rect 1635 3640 1669 3674
rect 1635 3572 1669 3606
rect 1635 3504 1669 3538
rect 1635 3436 1669 3470
rect 1635 3368 1669 3402
rect 1635 3300 1669 3334
rect 1635 3232 1669 3266
rect 1635 3164 1669 3198
rect 2627 4048 2661 4082
rect 2627 3980 2661 4014
rect 2627 3912 2661 3946
rect 2627 3844 2661 3878
rect 2627 3776 2661 3810
rect 2627 3708 2661 3742
rect 2627 3640 2661 3674
rect 2627 3572 2661 3606
rect 2627 3504 2661 3538
rect 2627 3436 2661 3470
rect 2627 3368 2661 3402
rect 2627 3300 2661 3334
rect 2627 3232 2661 3266
rect 2627 3164 2661 3198
rect 3619 4048 3653 4082
rect 3619 3980 3653 4014
rect 3619 3912 3653 3946
rect 3619 3844 3653 3878
rect 3619 3776 3653 3810
rect 3619 3708 3653 3742
rect 3619 3640 3653 3674
rect 3619 3572 3653 3606
rect 3619 3504 3653 3538
rect 3619 3436 3653 3470
rect 3619 3368 3653 3402
rect 3619 3300 3653 3334
rect 3619 3232 3653 3266
rect 3619 3164 3653 3198
rect 4611 4048 4645 4082
rect 4611 3980 4645 4014
rect 4611 3912 4645 3946
rect 4611 3844 4645 3878
rect 4611 3776 4645 3810
rect 4611 3708 4645 3742
rect 4611 3640 4645 3674
rect 4611 3572 4645 3606
rect 4611 3504 4645 3538
rect 4611 3436 4645 3470
rect 4611 3368 4645 3402
rect 4611 3300 4645 3334
rect 4611 3232 4645 3266
rect 4611 3164 4645 3198
rect 5603 4048 5637 4082
rect 5603 3980 5637 4014
rect 5603 3912 5637 3946
rect 5603 3844 5637 3878
rect 5603 3776 5637 3810
rect 5603 3708 5637 3742
rect 5603 3640 5637 3674
rect 5603 3572 5637 3606
rect 5603 3504 5637 3538
rect 5603 3436 5637 3470
rect 5603 3368 5637 3402
rect 5603 3300 5637 3334
rect 5603 3232 5637 3266
rect 5603 3164 5637 3198
rect 6595 4048 6629 4082
rect 6595 3980 6629 4014
rect 6595 3912 6629 3946
rect 6595 3844 6629 3878
rect 6595 3776 6629 3810
rect 6595 3708 6629 3742
rect 6595 3640 6629 3674
rect 6595 3572 6629 3606
rect 6595 3504 6629 3538
rect 6595 3436 6629 3470
rect 6595 3368 6629 3402
rect 6595 3300 6629 3334
rect 6595 3232 6629 3266
rect 6595 3164 6629 3198
rect 7587 4048 7621 4082
rect 7587 3980 7621 4014
rect 7587 3912 7621 3946
rect 7587 3844 7621 3878
rect 7587 3776 7621 3810
rect 7587 3708 7621 3742
rect 7587 3640 7621 3674
rect 7587 3572 7621 3606
rect 7587 3504 7621 3538
rect 7587 3436 7621 3470
rect 7587 3368 7621 3402
rect 7587 3300 7621 3334
rect 7587 3232 7621 3266
rect 7587 3164 7621 3198
rect 8579 4048 8613 4082
rect 8579 3980 8613 4014
rect 8579 3912 8613 3946
rect 8579 3844 8613 3878
rect 8579 3776 8613 3810
rect 8579 3708 8613 3742
rect 8579 3640 8613 3674
rect 8579 3572 8613 3606
rect 8579 3504 8613 3538
rect 8579 3436 8613 3470
rect 8579 3368 8613 3402
rect 8579 3300 8613 3334
rect 8579 3232 8613 3266
rect 8579 3164 8613 3198
rect 9571 4048 9605 4082
rect 9571 3980 9605 4014
rect 9571 3912 9605 3946
rect 9571 3844 9605 3878
rect 9571 3776 9605 3810
rect 9571 3708 9605 3742
rect 9571 3640 9605 3674
rect 9571 3572 9605 3606
rect 9571 3504 9605 3538
rect 9571 3436 9605 3470
rect 9571 3368 9605 3402
rect 9571 3300 9605 3334
rect 9571 3232 9605 3266
rect 9571 3164 9605 3198
rect 10563 4048 10597 4082
rect 10563 3980 10597 4014
rect 10563 3912 10597 3946
rect 10563 3844 10597 3878
rect 10563 3776 10597 3810
rect 10563 3708 10597 3742
rect 10563 3640 10597 3674
rect 10563 3572 10597 3606
rect 10563 3504 10597 3538
rect 10563 3436 10597 3470
rect 10563 3368 10597 3402
rect 10563 3300 10597 3334
rect 10563 3232 10597 3266
rect 10563 3164 10597 3198
rect 11555 4048 11589 4082
rect 11555 3980 11589 4014
rect 11555 3912 11589 3946
rect 11555 3844 11589 3878
rect 11555 3776 11589 3810
rect 11555 3708 11589 3742
rect 11555 3640 11589 3674
rect 11555 3572 11589 3606
rect 11555 3504 11589 3538
rect 11555 3436 11589 3470
rect 11555 3368 11589 3402
rect 11555 3300 11589 3334
rect 11555 3232 11589 3266
rect 11555 3164 11589 3198
rect 12547 4048 12581 4082
rect 12547 3980 12581 4014
rect 12547 3912 12581 3946
rect 12547 3844 12581 3878
rect 12547 3776 12581 3810
rect 12547 3708 12581 3742
rect 12547 3640 12581 3674
rect 12547 3572 12581 3606
rect 12547 3504 12581 3538
rect 12547 3436 12581 3470
rect 12547 3368 12581 3402
rect 12547 3300 12581 3334
rect 12547 3232 12581 3266
rect 12547 3164 12581 3198
rect 13539 4048 13573 4082
rect 13539 3980 13573 4014
rect 13539 3912 13573 3946
rect 13539 3844 13573 3878
rect 13539 3776 13573 3810
rect 13539 3708 13573 3742
rect 13539 3640 13573 3674
rect 13539 3572 13573 3606
rect 13539 3504 13573 3538
rect 13539 3436 13573 3470
rect 13539 3368 13573 3402
rect 13539 3300 13573 3334
rect 13539 3232 13573 3266
rect 13539 3164 13573 3198
rect 14468 3992 14638 4502
rect 14468 3923 14502 3957
rect 14536 3924 14638 3992
rect 14604 3905 14638 3924
rect 14468 3854 14502 3888
rect 14536 3855 14570 3889
rect 14604 3837 14638 3871
rect 14468 3785 14502 3819
rect 14536 3786 14570 3820
rect 14604 3769 14638 3803
rect 14468 3716 14502 3750
rect 14536 3717 14570 3751
rect 14604 3701 14638 3735
rect 14468 3647 14502 3681
rect 14536 3648 14570 3682
rect 14604 3633 14638 3667
rect 14468 3578 14502 3612
rect 14536 3579 14570 3613
rect 14604 3565 14638 3599
rect 14468 3509 14502 3543
rect 14536 3510 14570 3544
rect 14604 3497 14638 3531
rect 14468 3440 14502 3474
rect 14536 3441 14570 3475
rect 14604 3429 14638 3463
rect 14468 3371 14502 3405
rect 14536 3372 14570 3406
rect 14604 3361 14638 3395
rect 14468 3302 14502 3336
rect 14536 3303 14570 3337
rect 14604 3293 14638 3327
rect 14468 3233 14502 3267
rect 14536 3234 14570 3268
rect 14604 3225 14638 3259
rect 14468 3164 14502 3198
rect 14536 3165 14570 3199
rect 14604 3157 14638 3191
rect 497 3094 531 3128
rect 565 3094 599 3128
rect 633 3094 667 3128
rect 497 3025 531 3059
rect 565 3025 599 3059
rect 633 3025 667 3059
rect 497 2956 531 2990
rect 565 2956 599 2990
rect 633 2956 667 2990
rect 497 2887 531 2921
rect 565 2887 599 2921
rect 633 2887 667 2921
rect 497 2818 531 2852
rect 565 2818 599 2852
rect 633 2818 667 2852
rect 497 2749 531 2783
rect 565 2749 599 2783
rect 633 2749 667 2783
rect 497 2680 531 2714
rect 565 2680 599 2714
rect 633 2680 667 2714
rect 497 2611 531 2645
rect 565 2611 599 2645
rect 633 2611 667 2645
rect 497 2542 531 2576
rect 565 2542 599 2576
rect 633 2542 667 2576
rect 1601 3010 1635 3044
rect 1669 3010 1703 3044
rect 1601 2940 1635 2974
rect 1669 2940 1703 2974
rect 1601 2870 1635 2904
rect 1669 2870 1703 2904
rect 1601 2800 1635 2834
rect 1669 2800 1703 2834
rect 1601 2730 1635 2764
rect 1669 2730 1703 2764
rect 1601 2660 1635 2694
rect 1669 2660 1703 2694
rect 2593 3010 2627 3044
rect 2661 3010 2695 3044
rect 2593 2940 2627 2974
rect 2661 2940 2695 2974
rect 2593 2870 2627 2904
rect 2661 2870 2695 2904
rect 2593 2800 2627 2834
rect 2661 2800 2695 2834
rect 2593 2730 2627 2764
rect 2661 2730 2695 2764
rect 2593 2660 2627 2694
rect 2661 2660 2695 2694
rect 3585 3010 3619 3044
rect 3653 3010 3687 3044
rect 3585 2940 3619 2974
rect 3653 2940 3687 2974
rect 3585 2870 3619 2904
rect 3653 2870 3687 2904
rect 3585 2800 3619 2834
rect 3653 2800 3687 2834
rect 3585 2730 3619 2764
rect 3653 2730 3687 2764
rect 3585 2660 3619 2694
rect 3653 2660 3687 2694
rect 4577 3010 4611 3044
rect 4645 3010 4679 3044
rect 4577 2940 4611 2974
rect 4645 2940 4679 2974
rect 4577 2870 4611 2904
rect 4645 2870 4679 2904
rect 4577 2800 4611 2834
rect 4645 2800 4679 2834
rect 4577 2730 4611 2764
rect 4645 2730 4679 2764
rect 4577 2660 4611 2694
rect 4645 2660 4679 2694
rect 5569 3010 5603 3044
rect 5637 3010 5671 3044
rect 5569 2940 5603 2974
rect 5637 2940 5671 2974
rect 5569 2870 5603 2904
rect 5637 2870 5671 2904
rect 5569 2800 5603 2834
rect 5637 2800 5671 2834
rect 5569 2730 5603 2764
rect 5637 2730 5671 2764
rect 5569 2660 5603 2694
rect 5637 2660 5671 2694
rect 6561 3010 6595 3044
rect 6629 3010 6663 3044
rect 6561 2940 6595 2974
rect 6629 2940 6663 2974
rect 6561 2870 6595 2904
rect 6629 2870 6663 2904
rect 6561 2800 6595 2834
rect 6629 2800 6663 2834
rect 6561 2730 6595 2764
rect 6629 2730 6663 2764
rect 6561 2660 6595 2694
rect 6629 2660 6663 2694
rect 7553 3010 7587 3044
rect 7621 3010 7655 3044
rect 7553 2940 7587 2974
rect 7621 2940 7655 2974
rect 7553 2870 7587 2904
rect 7621 2870 7655 2904
rect 7553 2800 7587 2834
rect 7621 2800 7655 2834
rect 7553 2730 7587 2764
rect 7621 2730 7655 2764
rect 7553 2660 7587 2694
rect 7621 2660 7655 2694
rect 8545 3010 8579 3044
rect 8613 3010 8647 3044
rect 8545 2940 8579 2974
rect 8613 2940 8647 2974
rect 8545 2870 8579 2904
rect 8613 2870 8647 2904
rect 8545 2800 8579 2834
rect 8613 2800 8647 2834
rect 8545 2730 8579 2764
rect 8613 2730 8647 2764
rect 8545 2660 8579 2694
rect 8613 2660 8647 2694
rect 9537 3010 9571 3044
rect 9605 3010 9639 3044
rect 9537 2940 9571 2974
rect 9605 2940 9639 2974
rect 9537 2870 9571 2904
rect 9605 2870 9639 2904
rect 9537 2800 9571 2834
rect 9605 2800 9639 2834
rect 9537 2730 9571 2764
rect 9605 2730 9639 2764
rect 9537 2660 9571 2694
rect 9605 2660 9639 2694
rect 10529 3010 10563 3044
rect 10597 3010 10631 3044
rect 10529 2940 10563 2974
rect 10597 2940 10631 2974
rect 10529 2870 10563 2904
rect 10597 2870 10631 2904
rect 10529 2800 10563 2834
rect 10597 2800 10631 2834
rect 10529 2730 10563 2764
rect 10597 2730 10631 2764
rect 10529 2660 10563 2694
rect 10597 2660 10631 2694
rect 11521 3010 11555 3044
rect 11589 3010 11623 3044
rect 11521 2940 11555 2974
rect 11589 2940 11623 2974
rect 11521 2870 11555 2904
rect 11589 2870 11623 2904
rect 11521 2800 11555 2834
rect 11589 2800 11623 2834
rect 11521 2730 11555 2764
rect 11589 2730 11623 2764
rect 11521 2660 11555 2694
rect 11589 2660 11623 2694
rect 12513 3010 12547 3044
rect 12581 3010 12615 3044
rect 12513 2940 12547 2974
rect 12581 2940 12615 2974
rect 12513 2870 12547 2904
rect 12581 2870 12615 2904
rect 12513 2800 12547 2834
rect 12581 2800 12615 2834
rect 12513 2730 12547 2764
rect 12581 2730 12615 2764
rect 12513 2660 12547 2694
rect 12581 2660 12615 2694
rect 13505 3010 13539 3044
rect 13573 3010 13607 3044
rect 13505 2940 13539 2974
rect 13573 2940 13607 2974
rect 13505 2870 13539 2904
rect 13573 2870 13607 2904
rect 13505 2800 13539 2834
rect 13573 2800 13607 2834
rect 13505 2730 13539 2764
rect 13573 2730 13607 2764
rect 13505 2660 13539 2694
rect 13573 2660 13607 2694
rect 14468 3095 14502 3129
rect 14536 3096 14570 3130
rect 14604 3089 14638 3123
rect 14468 3026 14502 3060
rect 14536 3027 14570 3061
rect 14604 3021 14638 3055
rect 14468 2957 14502 2991
rect 14536 2958 14570 2992
rect 14604 2953 14638 2987
rect 14468 2888 14502 2922
rect 14536 2889 14570 2923
rect 14604 2885 14638 2919
rect 14468 2819 14502 2853
rect 14536 2820 14570 2854
rect 14604 2817 14638 2851
rect 14468 2750 14502 2784
rect 14536 2751 14570 2785
rect 14604 2749 14638 2783
rect 14468 2681 14502 2715
rect 14536 2682 14570 2716
rect 14604 2681 14638 2715
rect 14468 2612 14502 2646
rect 14536 2613 14570 2647
rect 14604 2613 14638 2647
rect 497 2473 531 2507
rect 565 2473 599 2507
rect 633 2473 667 2507
rect 497 2404 531 2438
rect 565 2404 599 2438
rect 633 2404 667 2438
rect 497 2335 531 2369
rect 565 2335 599 2369
rect 633 2335 667 2369
rect 497 2266 531 2300
rect 565 2266 599 2300
rect 633 2266 667 2300
rect 497 2197 531 2231
rect 565 2197 599 2231
rect 633 2197 667 2231
rect 497 2129 531 2163
rect 565 2128 599 2162
rect 633 2128 667 2162
rect 497 2061 531 2095
rect 565 2059 599 2093
rect 633 2059 667 2093
rect 497 1993 531 2027
rect 565 1990 599 2024
rect 633 1990 667 2024
rect 497 1925 531 1959
rect 565 1921 599 1955
rect 633 1921 667 1955
rect 497 1857 531 1891
rect 565 1852 599 1886
rect 633 1852 667 1886
rect 497 1789 531 1823
rect 565 1783 599 1817
rect 633 1783 667 1817
rect 497 1721 531 1755
rect 565 1714 599 1748
rect 633 1714 667 1748
rect 497 1653 531 1687
rect 565 1645 599 1679
rect 633 1645 667 1679
rect 497 1585 531 1619
rect 565 1576 599 1610
rect 633 1576 667 1610
rect 1635 2506 1669 2540
rect 1635 2438 1669 2472
rect 1635 2370 1669 2404
rect 1635 2302 1669 2336
rect 1635 2234 1669 2268
rect 1635 2166 1669 2200
rect 1635 2098 1669 2132
rect 1635 2030 1669 2064
rect 1635 1962 1669 1996
rect 1635 1894 1669 1928
rect 1635 1826 1669 1860
rect 1635 1758 1669 1792
rect 1635 1690 1669 1724
rect 1635 1622 1669 1656
rect 2627 2506 2661 2540
rect 2627 2438 2661 2472
rect 2627 2370 2661 2404
rect 2627 2302 2661 2336
rect 2627 2234 2661 2268
rect 2627 2166 2661 2200
rect 2627 2098 2661 2132
rect 2627 2030 2661 2064
rect 2627 1962 2661 1996
rect 2627 1894 2661 1928
rect 2627 1826 2661 1860
rect 2627 1758 2661 1792
rect 2627 1690 2661 1724
rect 2627 1622 2661 1656
rect 3619 2506 3653 2540
rect 3619 2438 3653 2472
rect 3619 2370 3653 2404
rect 3619 2302 3653 2336
rect 3619 2234 3653 2268
rect 3619 2166 3653 2200
rect 3619 2098 3653 2132
rect 3619 2030 3653 2064
rect 3619 1962 3653 1996
rect 3619 1894 3653 1928
rect 3619 1826 3653 1860
rect 3619 1758 3653 1792
rect 3619 1690 3653 1724
rect 3619 1622 3653 1656
rect 4611 2506 4645 2540
rect 4611 2438 4645 2472
rect 4611 2370 4645 2404
rect 4611 2302 4645 2336
rect 4611 2234 4645 2268
rect 4611 2166 4645 2200
rect 4611 2098 4645 2132
rect 4611 2030 4645 2064
rect 4611 1962 4645 1996
rect 4611 1894 4645 1928
rect 4611 1826 4645 1860
rect 4611 1758 4645 1792
rect 4611 1690 4645 1724
rect 4611 1622 4645 1656
rect 5603 2506 5637 2540
rect 5603 2438 5637 2472
rect 5603 2370 5637 2404
rect 5603 2302 5637 2336
rect 5603 2234 5637 2268
rect 5603 2166 5637 2200
rect 5603 2098 5637 2132
rect 5603 2030 5637 2064
rect 5603 1962 5637 1996
rect 5603 1894 5637 1928
rect 5603 1826 5637 1860
rect 5603 1758 5637 1792
rect 5603 1690 5637 1724
rect 5603 1622 5637 1656
rect 6595 2506 6629 2540
rect 6595 2438 6629 2472
rect 6595 2370 6629 2404
rect 6595 2302 6629 2336
rect 6595 2234 6629 2268
rect 6595 2166 6629 2200
rect 6595 2098 6629 2132
rect 6595 2030 6629 2064
rect 6595 1962 6629 1996
rect 6595 1894 6629 1928
rect 6595 1826 6629 1860
rect 6595 1758 6629 1792
rect 6595 1690 6629 1724
rect 6595 1622 6629 1656
rect 7587 2506 7621 2540
rect 7587 2438 7621 2472
rect 7587 2370 7621 2404
rect 7587 2302 7621 2336
rect 7587 2234 7621 2268
rect 7587 2166 7621 2200
rect 7587 2098 7621 2132
rect 7587 2030 7621 2064
rect 7587 1962 7621 1996
rect 7587 1894 7621 1928
rect 7587 1826 7621 1860
rect 7587 1758 7621 1792
rect 7587 1690 7621 1724
rect 7587 1622 7621 1656
rect 8579 2506 8613 2540
rect 8579 2438 8613 2472
rect 8579 2370 8613 2404
rect 8579 2302 8613 2336
rect 8579 2234 8613 2268
rect 8579 2166 8613 2200
rect 8579 2098 8613 2132
rect 8579 2030 8613 2064
rect 8579 1962 8613 1996
rect 8579 1894 8613 1928
rect 8579 1826 8613 1860
rect 8579 1758 8613 1792
rect 8579 1690 8613 1724
rect 8579 1622 8613 1656
rect 9571 2506 9605 2540
rect 9571 2438 9605 2472
rect 9571 2370 9605 2404
rect 9571 2302 9605 2336
rect 9571 2234 9605 2268
rect 9571 2166 9605 2200
rect 9571 2098 9605 2132
rect 9571 2030 9605 2064
rect 9571 1962 9605 1996
rect 9571 1894 9605 1928
rect 9571 1826 9605 1860
rect 9571 1758 9605 1792
rect 9571 1690 9605 1724
rect 9571 1622 9605 1656
rect 10563 2506 10597 2540
rect 10563 2438 10597 2472
rect 10563 2370 10597 2404
rect 10563 2302 10597 2336
rect 10563 2234 10597 2268
rect 10563 2166 10597 2200
rect 10563 2098 10597 2132
rect 10563 2030 10597 2064
rect 10563 1962 10597 1996
rect 10563 1894 10597 1928
rect 10563 1826 10597 1860
rect 10563 1758 10597 1792
rect 10563 1690 10597 1724
rect 10563 1622 10597 1656
rect 11555 2506 11589 2540
rect 11555 2438 11589 2472
rect 11555 2370 11589 2404
rect 11555 2302 11589 2336
rect 11555 2234 11589 2268
rect 11555 2166 11589 2200
rect 11555 2098 11589 2132
rect 11555 2030 11589 2064
rect 11555 1962 11589 1996
rect 11555 1894 11589 1928
rect 11555 1826 11589 1860
rect 11555 1758 11589 1792
rect 11555 1690 11589 1724
rect 11555 1622 11589 1656
rect 12547 2506 12581 2540
rect 12547 2438 12581 2472
rect 12547 2370 12581 2404
rect 12547 2302 12581 2336
rect 12547 2234 12581 2268
rect 12547 2166 12581 2200
rect 12547 2098 12581 2132
rect 12547 2030 12581 2064
rect 12547 1962 12581 1996
rect 12547 1894 12581 1928
rect 12547 1826 12581 1860
rect 12547 1758 12581 1792
rect 12547 1690 12581 1724
rect 12547 1622 12581 1656
rect 13539 2506 13573 2540
rect 13539 2438 13573 2472
rect 13539 2370 13573 2404
rect 13539 2302 13573 2336
rect 13539 2234 13573 2268
rect 13539 2166 13573 2200
rect 13539 2098 13573 2132
rect 13539 2030 13573 2064
rect 13539 1962 13573 1996
rect 13539 1894 13573 1928
rect 13539 1826 13573 1860
rect 13539 1758 13573 1792
rect 13539 1690 13573 1724
rect 13539 1622 13573 1656
rect 14468 2543 14502 2577
rect 14536 2544 14570 2578
rect 14604 2545 14638 2579
rect 14468 2474 14502 2508
rect 14536 2475 14570 2509
rect 14604 2477 14638 2511
rect 14468 2405 14502 2439
rect 14536 2406 14570 2440
rect 14604 2409 14638 2443
rect 14468 2336 14502 2370
rect 14536 2337 14570 2371
rect 14604 2341 14638 2375
rect 14468 2267 14502 2301
rect 14536 2268 14570 2302
rect 14604 2273 14638 2307
rect 14468 2198 14502 2232
rect 14536 2199 14570 2233
rect 14604 2205 14638 2239
rect 14468 2129 14502 2163
rect 14536 2130 14570 2164
rect 14604 2137 14638 2171
rect 14468 2060 14502 2094
rect 14536 2061 14570 2095
rect 14604 2069 14638 2103
rect 14468 1991 14502 2025
rect 14536 1992 14570 2026
rect 14604 2001 14638 2035
rect 14468 1922 14502 1956
rect 14536 1923 14570 1957
rect 14604 1933 14638 1967
rect 14468 1853 14502 1887
rect 14536 1854 14570 1888
rect 14604 1865 14638 1899
rect 14468 1784 14502 1818
rect 14536 1785 14570 1819
rect 14604 1797 14638 1831
rect 14468 1715 14502 1749
rect 14536 1716 14570 1750
rect 14604 1729 14638 1763
rect 14468 1646 14502 1680
rect 14536 1647 14570 1681
rect 14604 1661 14638 1695
rect 14468 1577 14502 1611
rect 14536 1578 14570 1612
rect 14604 1593 14638 1627
rect 497 1517 531 1551
rect 565 1507 599 1541
rect 633 1507 667 1541
rect 497 1449 531 1483
rect 565 1438 599 1472
rect 633 1438 667 1472
rect 497 1381 531 1415
rect 565 1369 599 1403
rect 633 1369 667 1403
rect 14468 1508 14502 1542
rect 14536 1509 14570 1543
rect 14604 1525 14638 1559
rect 14468 1439 14502 1473
rect 14536 1440 14570 1474
rect 14604 1457 14638 1491
rect 497 1313 531 1347
rect 565 1300 599 1334
rect 633 1300 667 1334
rect 497 1245 531 1279
rect 565 1231 599 1265
rect 633 1231 667 1265
rect 497 1177 531 1211
rect 565 1162 599 1196
rect 633 1162 667 1196
rect 497 1109 531 1143
rect 565 1093 599 1127
rect 633 1093 667 1127
rect 497 1041 531 1075
rect 565 1024 599 1058
rect 633 1024 667 1058
rect 497 973 531 1007
rect 565 955 599 989
rect 633 955 667 989
rect 497 920 531 939
rect 497 818 667 920
rect 14468 1370 14502 1404
rect 14536 1371 14570 1405
rect 14604 1389 14638 1423
rect 14468 1301 14502 1335
rect 14536 1302 14570 1336
rect 14604 1321 14638 1355
rect 14468 1232 14502 1266
rect 14536 1233 14570 1267
rect 14604 1253 14638 1287
rect 14468 1163 14502 1197
rect 14536 1164 14570 1198
rect 14604 1184 14638 1218
rect 14468 1094 14502 1128
rect 14536 1095 14570 1129
rect 14604 1115 14638 1149
rect 14468 1025 14502 1059
rect 14536 1026 14570 1060
rect 14604 1046 14638 1080
rect 14468 956 14502 990
rect 14536 957 14570 991
rect 14604 977 14638 1011
rect 14468 887 14502 921
rect 14536 888 14570 922
rect 14604 908 14638 942
rect 702 818 736 852
rect 771 818 805 852
rect 840 818 874 852
rect 909 818 943 852
rect 978 818 1012 852
rect 1047 818 1081 852
rect 1116 818 1150 852
rect 1185 818 1219 852
rect 1254 818 1288 852
rect 1323 818 1357 852
rect 1392 818 1426 852
rect 1461 818 1495 852
rect 1530 818 1564 852
rect 1599 818 1633 852
rect 1668 818 1702 852
rect 1737 818 1771 852
rect 1806 818 1840 852
rect 1875 818 1909 852
rect 1944 818 1978 852
rect 2013 818 2047 852
rect 2082 818 2116 852
rect 2151 818 2185 852
rect 2220 818 2254 852
rect 2289 818 2323 852
rect 2358 818 2392 852
rect 2427 818 2461 852
rect 2496 818 2530 852
rect 2565 818 2599 852
rect 2634 818 2668 852
rect 2703 818 2737 852
rect 497 769 599 818
rect 2772 784 14502 852
rect 14536 819 14570 853
rect 14604 839 14638 873
rect 565 750 599 769
rect 634 750 668 784
rect 703 750 737 784
rect 772 750 806 784
rect 841 750 875 784
rect 910 750 944 784
rect 979 750 1013 784
rect 1048 750 1082 784
rect 1117 750 1151 784
rect 1186 750 1220 784
rect 1255 750 1289 784
rect 1324 750 1358 784
rect 1393 750 1427 784
rect 1462 750 1496 784
rect 1531 750 1565 784
rect 1600 750 1634 784
rect 1669 750 1703 784
rect 1738 750 1772 784
rect 1807 750 1841 784
rect 1876 750 1910 784
rect 1945 750 1979 784
rect 2014 750 2048 784
rect 2083 750 2117 784
rect 2152 750 2186 784
rect 2221 750 2255 784
rect 2290 750 2324 784
rect 2359 750 2393 784
rect 2428 750 2462 784
rect 2497 750 2531 784
rect 2566 750 2600 784
rect 2635 750 2669 784
rect 2704 750 2738 784
rect 2772 750 14570 784
rect 14604 770 14638 804
rect 516 682 550 716
rect 585 682 619 716
rect 654 682 688 716
rect 723 682 757 716
rect 792 682 826 716
rect 861 682 895 716
rect 930 682 964 716
rect 999 682 1033 716
rect 1068 682 1102 716
rect 1137 682 1171 716
rect 1206 682 1240 716
rect 1275 682 1309 716
rect 1344 682 1378 716
rect 1413 682 1447 716
rect 1482 682 1516 716
rect 1551 682 1585 716
rect 1620 682 1654 716
rect 1689 682 1723 716
rect 1758 682 1792 716
rect 1827 682 1861 716
rect 1896 682 1930 716
rect 1965 682 1999 716
rect 2034 682 2068 716
rect 2103 682 2137 716
rect 2172 682 2206 716
rect 2241 682 2275 716
rect 2310 682 2344 716
rect 2379 682 2413 716
rect 2448 682 2482 716
rect 2517 682 2551 716
rect 2586 682 2620 716
rect 2655 682 2689 716
rect 2724 682 2758 716
rect 2793 682 2827 716
rect 2862 682 2896 716
rect 2931 682 2965 716
rect 3000 682 3034 716
rect 3069 682 3103 716
rect 3138 682 3172 716
rect 3207 682 3241 716
rect 3276 682 3310 716
rect 3345 682 3379 716
rect 3414 682 3448 716
rect 3483 682 3517 716
rect 3552 682 3586 716
rect 3621 682 3655 716
rect 3690 682 3724 716
rect 3759 682 3793 716
rect 3828 682 3862 716
rect 3897 682 3931 716
rect 3966 682 4000 716
rect 4035 682 4069 716
rect 4104 682 4138 716
rect 4173 682 4207 716
rect 4242 682 4276 716
rect 4311 682 4345 716
rect 4380 682 4414 716
rect 4449 682 4483 716
rect 4518 682 4552 716
rect 4587 682 4621 716
rect 4656 682 4690 716
rect 4725 682 14551 750
rect 14604 701 14638 735
<< poly >>
rect 881 4308 1001 4324
rect 881 4274 924 4308
rect 958 4274 1001 4308
rect 881 4234 1001 4274
rect 881 4200 924 4234
rect 958 4200 1001 4234
rect 881 4152 1001 4200
rect 1311 4308 1431 4324
rect 1311 4274 1354 4308
rect 1388 4274 1431 4308
rect 1311 4234 1431 4274
rect 1311 4200 1354 4234
rect 1388 4200 1431 4234
rect 1311 4152 1431 4200
rect 1873 4308 1993 4324
rect 1873 4274 1916 4308
rect 1950 4274 1993 4308
rect 1873 4234 1993 4274
rect 1873 4200 1916 4234
rect 1950 4200 1993 4234
rect 1873 4152 1993 4200
rect 2303 4308 2423 4324
rect 2303 4274 2346 4308
rect 2380 4274 2423 4308
rect 2303 4234 2423 4274
rect 2303 4200 2346 4234
rect 2380 4200 2423 4234
rect 2303 4152 2423 4200
rect 2865 4308 2985 4324
rect 2865 4274 2908 4308
rect 2942 4274 2985 4308
rect 2865 4234 2985 4274
rect 2865 4200 2908 4234
rect 2942 4200 2985 4234
rect 2865 4152 2985 4200
rect 3295 4308 3415 4324
rect 3295 4274 3338 4308
rect 3372 4274 3415 4308
rect 3295 4234 3415 4274
rect 3295 4200 3338 4234
rect 3372 4200 3415 4234
rect 3295 4152 3415 4200
rect 3857 4308 3977 4324
rect 3857 4274 3900 4308
rect 3934 4274 3977 4308
rect 3857 4234 3977 4274
rect 3857 4200 3900 4234
rect 3934 4200 3977 4234
rect 3857 4152 3977 4200
rect 4287 4308 4407 4324
rect 4287 4274 4330 4308
rect 4364 4274 4407 4308
rect 4287 4234 4407 4274
rect 4287 4200 4330 4234
rect 4364 4200 4407 4234
rect 4287 4152 4407 4200
rect 4849 4308 4969 4324
rect 4849 4274 4892 4308
rect 4926 4274 4969 4308
rect 4849 4234 4969 4274
rect 4849 4200 4892 4234
rect 4926 4200 4969 4234
rect 4849 4152 4969 4200
rect 5279 4308 5399 4324
rect 5279 4274 5322 4308
rect 5356 4274 5399 4308
rect 5279 4234 5399 4274
rect 5279 4200 5322 4234
rect 5356 4200 5399 4234
rect 5279 4152 5399 4200
rect 5841 4308 5961 4324
rect 5841 4274 5884 4308
rect 5918 4274 5961 4308
rect 5841 4234 5961 4274
rect 5841 4200 5884 4234
rect 5918 4200 5961 4234
rect 5841 4152 5961 4200
rect 6271 4308 6391 4324
rect 6271 4274 6314 4308
rect 6348 4274 6391 4308
rect 6271 4234 6391 4274
rect 6271 4200 6314 4234
rect 6348 4200 6391 4234
rect 6271 4152 6391 4200
rect 6833 4308 6953 4324
rect 6833 4274 6876 4308
rect 6910 4274 6953 4308
rect 6833 4234 6953 4274
rect 6833 4200 6876 4234
rect 6910 4200 6953 4234
rect 6833 4152 6953 4200
rect 7263 4308 7383 4324
rect 7263 4274 7306 4308
rect 7340 4274 7383 4308
rect 7263 4234 7383 4274
rect 7263 4200 7306 4234
rect 7340 4200 7383 4234
rect 7263 4152 7383 4200
rect 7825 4308 7945 4324
rect 7825 4274 7868 4308
rect 7902 4274 7945 4308
rect 7825 4234 7945 4274
rect 7825 4200 7868 4234
rect 7902 4200 7945 4234
rect 7825 4152 7945 4200
rect 8255 4308 8375 4324
rect 8255 4274 8298 4308
rect 8332 4274 8375 4308
rect 8255 4234 8375 4274
rect 8255 4200 8298 4234
rect 8332 4200 8375 4234
rect 8255 4152 8375 4200
rect 8817 4308 8937 4324
rect 8817 4274 8860 4308
rect 8894 4274 8937 4308
rect 8817 4234 8937 4274
rect 8817 4200 8860 4234
rect 8894 4200 8937 4234
rect 8817 4152 8937 4200
rect 9247 4308 9367 4324
rect 9247 4274 9290 4308
rect 9324 4274 9367 4308
rect 9247 4234 9367 4274
rect 9247 4200 9290 4234
rect 9324 4200 9367 4234
rect 9247 4152 9367 4200
rect 9809 4308 9929 4324
rect 9809 4274 9852 4308
rect 9886 4274 9929 4308
rect 9809 4234 9929 4274
rect 9809 4200 9852 4234
rect 9886 4200 9929 4234
rect 9809 4152 9929 4200
rect 10239 4308 10359 4324
rect 10239 4274 10282 4308
rect 10316 4274 10359 4308
rect 10239 4234 10359 4274
rect 10239 4200 10282 4234
rect 10316 4200 10359 4234
rect 10239 4152 10359 4200
rect 10801 4308 10921 4324
rect 10801 4274 10844 4308
rect 10878 4274 10921 4308
rect 10801 4234 10921 4274
rect 10801 4200 10844 4234
rect 10878 4200 10921 4234
rect 10801 4152 10921 4200
rect 11231 4308 11351 4324
rect 11231 4274 11274 4308
rect 11308 4274 11351 4308
rect 11231 4234 11351 4274
rect 11231 4200 11274 4234
rect 11308 4200 11351 4234
rect 11231 4152 11351 4200
rect 11793 4308 11913 4324
rect 11793 4274 11836 4308
rect 11870 4274 11913 4308
rect 11793 4234 11913 4274
rect 11793 4200 11836 4234
rect 11870 4200 11913 4234
rect 11793 4152 11913 4200
rect 12223 4308 12343 4324
rect 12223 4274 12266 4308
rect 12300 4274 12343 4308
rect 12223 4234 12343 4274
rect 12223 4200 12266 4234
rect 12300 4200 12343 4234
rect 12223 4152 12343 4200
rect 12785 4308 12905 4324
rect 12785 4274 12828 4308
rect 12862 4274 12905 4308
rect 12785 4234 12905 4274
rect 12785 4200 12828 4234
rect 12862 4200 12905 4234
rect 12785 4152 12905 4200
rect 13215 4308 13335 4324
rect 13215 4274 13258 4308
rect 13292 4274 13335 4308
rect 13215 4234 13335 4274
rect 13215 4200 13258 4234
rect 13292 4200 13335 4234
rect 13215 4152 13335 4200
rect 13777 4308 13897 4324
rect 13777 4274 13820 4308
rect 13854 4274 13897 4308
rect 13777 4234 13897 4274
rect 13777 4200 13820 4234
rect 13854 4200 13897 4234
rect 13777 4152 13897 4200
rect 14135 4308 14255 4324
rect 14135 4274 14178 4308
rect 14212 4274 14255 4308
rect 14135 4234 14255 4274
rect 14135 4200 14178 4234
rect 14212 4200 14255 4234
rect 14135 4152 14255 4200
rect 881 3104 1001 3152
rect 881 3070 924 3104
rect 958 3070 1001 3104
rect 881 3026 1001 3070
rect 881 2992 924 3026
rect 958 2992 1001 3026
rect 881 2948 1001 2992
rect 881 2914 924 2948
rect 958 2914 1001 2948
rect 881 2870 1001 2914
rect 881 2836 924 2870
rect 958 2836 1001 2870
rect 881 2792 1001 2836
rect 881 2758 924 2792
rect 958 2758 1001 2792
rect 881 2713 1001 2758
rect 881 2679 924 2713
rect 958 2679 1001 2713
rect 881 2634 1001 2679
rect 881 2600 924 2634
rect 958 2600 1001 2634
rect 881 2552 1001 2600
rect 1311 3104 1431 3152
rect 1311 3070 1354 3104
rect 1388 3070 1431 3104
rect 1873 3104 1993 3152
rect 1311 3026 1431 3070
rect 1311 2992 1354 3026
rect 1388 2992 1431 3026
rect 1311 2948 1431 2992
rect 1311 2914 1354 2948
rect 1388 2914 1431 2948
rect 1311 2870 1431 2914
rect 1311 2836 1354 2870
rect 1388 2836 1431 2870
rect 1311 2792 1431 2836
rect 1311 2758 1354 2792
rect 1388 2758 1431 2792
rect 1311 2713 1431 2758
rect 1311 2679 1354 2713
rect 1388 2679 1431 2713
rect 1311 2634 1431 2679
rect 1311 2600 1354 2634
rect 1388 2600 1431 2634
rect 1873 3070 1916 3104
rect 1950 3070 1993 3104
rect 1873 3026 1993 3070
rect 1873 2992 1916 3026
rect 1950 2992 1993 3026
rect 1873 2948 1993 2992
rect 1873 2914 1916 2948
rect 1950 2914 1993 2948
rect 1873 2870 1993 2914
rect 1873 2836 1916 2870
rect 1950 2836 1993 2870
rect 1873 2792 1993 2836
rect 1873 2758 1916 2792
rect 1950 2758 1993 2792
rect 1873 2713 1993 2758
rect 1873 2679 1916 2713
rect 1950 2679 1993 2713
rect 1873 2634 1993 2679
rect 1311 2552 1431 2600
rect 1873 2600 1916 2634
rect 1950 2600 1993 2634
rect 1873 2552 1993 2600
rect 2303 3104 2423 3152
rect 2303 3070 2346 3104
rect 2380 3070 2423 3104
rect 2865 3104 2985 3152
rect 2303 3026 2423 3070
rect 2303 2992 2346 3026
rect 2380 2992 2423 3026
rect 2303 2948 2423 2992
rect 2303 2914 2346 2948
rect 2380 2914 2423 2948
rect 2303 2870 2423 2914
rect 2303 2836 2346 2870
rect 2380 2836 2423 2870
rect 2303 2792 2423 2836
rect 2303 2758 2346 2792
rect 2380 2758 2423 2792
rect 2303 2713 2423 2758
rect 2303 2679 2346 2713
rect 2380 2679 2423 2713
rect 2303 2634 2423 2679
rect 2303 2600 2346 2634
rect 2380 2600 2423 2634
rect 2865 3070 2908 3104
rect 2942 3070 2985 3104
rect 2865 3026 2985 3070
rect 2865 2992 2908 3026
rect 2942 2992 2985 3026
rect 2865 2948 2985 2992
rect 2865 2914 2908 2948
rect 2942 2914 2985 2948
rect 2865 2870 2985 2914
rect 2865 2836 2908 2870
rect 2942 2836 2985 2870
rect 2865 2792 2985 2836
rect 2865 2758 2908 2792
rect 2942 2758 2985 2792
rect 2865 2713 2985 2758
rect 2865 2679 2908 2713
rect 2942 2679 2985 2713
rect 2865 2634 2985 2679
rect 2303 2552 2423 2600
rect 2865 2600 2908 2634
rect 2942 2600 2985 2634
rect 2865 2552 2985 2600
rect 3295 3104 3415 3152
rect 3295 3070 3338 3104
rect 3372 3070 3415 3104
rect 3857 3104 3977 3152
rect 3295 3026 3415 3070
rect 3295 2992 3338 3026
rect 3372 2992 3415 3026
rect 3295 2948 3415 2992
rect 3295 2914 3338 2948
rect 3372 2914 3415 2948
rect 3295 2870 3415 2914
rect 3295 2836 3338 2870
rect 3372 2836 3415 2870
rect 3295 2792 3415 2836
rect 3295 2758 3338 2792
rect 3372 2758 3415 2792
rect 3295 2713 3415 2758
rect 3295 2679 3338 2713
rect 3372 2679 3415 2713
rect 3295 2634 3415 2679
rect 3295 2600 3338 2634
rect 3372 2600 3415 2634
rect 3857 3070 3900 3104
rect 3934 3070 3977 3104
rect 3857 3026 3977 3070
rect 3857 2992 3900 3026
rect 3934 2992 3977 3026
rect 3857 2948 3977 2992
rect 3857 2914 3900 2948
rect 3934 2914 3977 2948
rect 3857 2870 3977 2914
rect 3857 2836 3900 2870
rect 3934 2836 3977 2870
rect 3857 2792 3977 2836
rect 3857 2758 3900 2792
rect 3934 2758 3977 2792
rect 3857 2713 3977 2758
rect 3857 2679 3900 2713
rect 3934 2679 3977 2713
rect 3857 2634 3977 2679
rect 3295 2552 3415 2600
rect 3857 2600 3900 2634
rect 3934 2600 3977 2634
rect 3857 2552 3977 2600
rect 4287 3104 4407 3152
rect 4287 3070 4330 3104
rect 4364 3070 4407 3104
rect 4849 3104 4969 3152
rect 4287 3026 4407 3070
rect 4287 2992 4330 3026
rect 4364 2992 4407 3026
rect 4287 2948 4407 2992
rect 4287 2914 4330 2948
rect 4364 2914 4407 2948
rect 4287 2870 4407 2914
rect 4287 2836 4330 2870
rect 4364 2836 4407 2870
rect 4287 2792 4407 2836
rect 4287 2758 4330 2792
rect 4364 2758 4407 2792
rect 4287 2713 4407 2758
rect 4287 2679 4330 2713
rect 4364 2679 4407 2713
rect 4287 2634 4407 2679
rect 4287 2600 4330 2634
rect 4364 2600 4407 2634
rect 4849 3070 4892 3104
rect 4926 3070 4969 3104
rect 4849 3026 4969 3070
rect 4849 2992 4892 3026
rect 4926 2992 4969 3026
rect 4849 2948 4969 2992
rect 4849 2914 4892 2948
rect 4926 2914 4969 2948
rect 4849 2870 4969 2914
rect 4849 2836 4892 2870
rect 4926 2836 4969 2870
rect 4849 2792 4969 2836
rect 4849 2758 4892 2792
rect 4926 2758 4969 2792
rect 4849 2713 4969 2758
rect 4849 2679 4892 2713
rect 4926 2679 4969 2713
rect 4849 2634 4969 2679
rect 4287 2552 4407 2600
rect 4849 2600 4892 2634
rect 4926 2600 4969 2634
rect 4849 2552 4969 2600
rect 5279 3104 5399 3152
rect 5279 3070 5322 3104
rect 5356 3070 5399 3104
rect 5841 3104 5961 3152
rect 5279 3026 5399 3070
rect 5279 2992 5322 3026
rect 5356 2992 5399 3026
rect 5279 2948 5399 2992
rect 5279 2914 5322 2948
rect 5356 2914 5399 2948
rect 5279 2870 5399 2914
rect 5279 2836 5322 2870
rect 5356 2836 5399 2870
rect 5279 2792 5399 2836
rect 5279 2758 5322 2792
rect 5356 2758 5399 2792
rect 5279 2713 5399 2758
rect 5279 2679 5322 2713
rect 5356 2679 5399 2713
rect 5279 2634 5399 2679
rect 5279 2600 5322 2634
rect 5356 2600 5399 2634
rect 5841 3070 5884 3104
rect 5918 3070 5961 3104
rect 5841 3026 5961 3070
rect 5841 2992 5884 3026
rect 5918 2992 5961 3026
rect 5841 2948 5961 2992
rect 5841 2914 5884 2948
rect 5918 2914 5961 2948
rect 5841 2870 5961 2914
rect 5841 2836 5884 2870
rect 5918 2836 5961 2870
rect 5841 2792 5961 2836
rect 5841 2758 5884 2792
rect 5918 2758 5961 2792
rect 5841 2713 5961 2758
rect 5841 2679 5884 2713
rect 5918 2679 5961 2713
rect 5841 2634 5961 2679
rect 5279 2552 5399 2600
rect 5841 2600 5884 2634
rect 5918 2600 5961 2634
rect 5841 2552 5961 2600
rect 6271 3104 6391 3152
rect 6271 3070 6314 3104
rect 6348 3070 6391 3104
rect 6833 3104 6953 3152
rect 6271 3026 6391 3070
rect 6271 2992 6314 3026
rect 6348 2992 6391 3026
rect 6271 2948 6391 2992
rect 6271 2914 6314 2948
rect 6348 2914 6391 2948
rect 6271 2870 6391 2914
rect 6271 2836 6314 2870
rect 6348 2836 6391 2870
rect 6271 2792 6391 2836
rect 6271 2758 6314 2792
rect 6348 2758 6391 2792
rect 6271 2713 6391 2758
rect 6271 2679 6314 2713
rect 6348 2679 6391 2713
rect 6271 2634 6391 2679
rect 6271 2600 6314 2634
rect 6348 2600 6391 2634
rect 6833 3070 6876 3104
rect 6910 3070 6953 3104
rect 6833 3026 6953 3070
rect 6833 2992 6876 3026
rect 6910 2992 6953 3026
rect 6833 2948 6953 2992
rect 6833 2914 6876 2948
rect 6910 2914 6953 2948
rect 6833 2870 6953 2914
rect 6833 2836 6876 2870
rect 6910 2836 6953 2870
rect 6833 2792 6953 2836
rect 6833 2758 6876 2792
rect 6910 2758 6953 2792
rect 6833 2713 6953 2758
rect 6833 2679 6876 2713
rect 6910 2679 6953 2713
rect 6833 2634 6953 2679
rect 6271 2552 6391 2600
rect 6833 2600 6876 2634
rect 6910 2600 6953 2634
rect 6833 2552 6953 2600
rect 7263 3104 7383 3152
rect 7263 3070 7306 3104
rect 7340 3070 7383 3104
rect 7825 3104 7945 3152
rect 7263 3026 7383 3070
rect 7263 2992 7306 3026
rect 7340 2992 7383 3026
rect 7263 2948 7383 2992
rect 7263 2914 7306 2948
rect 7340 2914 7383 2948
rect 7263 2870 7383 2914
rect 7263 2836 7306 2870
rect 7340 2836 7383 2870
rect 7263 2792 7383 2836
rect 7263 2758 7306 2792
rect 7340 2758 7383 2792
rect 7263 2713 7383 2758
rect 7263 2679 7306 2713
rect 7340 2679 7383 2713
rect 7263 2634 7383 2679
rect 7263 2600 7306 2634
rect 7340 2600 7383 2634
rect 7825 3070 7868 3104
rect 7902 3070 7945 3104
rect 7825 3026 7945 3070
rect 7825 2992 7868 3026
rect 7902 2992 7945 3026
rect 7825 2948 7945 2992
rect 7825 2914 7868 2948
rect 7902 2914 7945 2948
rect 7825 2870 7945 2914
rect 7825 2836 7868 2870
rect 7902 2836 7945 2870
rect 7825 2792 7945 2836
rect 7825 2758 7868 2792
rect 7902 2758 7945 2792
rect 7825 2713 7945 2758
rect 7825 2679 7868 2713
rect 7902 2679 7945 2713
rect 7825 2634 7945 2679
rect 7263 2552 7383 2600
rect 7825 2600 7868 2634
rect 7902 2600 7945 2634
rect 7825 2552 7945 2600
rect 8255 3104 8375 3152
rect 8255 3070 8298 3104
rect 8332 3070 8375 3104
rect 8817 3104 8937 3152
rect 8255 3026 8375 3070
rect 8255 2992 8298 3026
rect 8332 2992 8375 3026
rect 8255 2948 8375 2992
rect 8255 2914 8298 2948
rect 8332 2914 8375 2948
rect 8255 2870 8375 2914
rect 8255 2836 8298 2870
rect 8332 2836 8375 2870
rect 8255 2792 8375 2836
rect 8255 2758 8298 2792
rect 8332 2758 8375 2792
rect 8255 2713 8375 2758
rect 8255 2679 8298 2713
rect 8332 2679 8375 2713
rect 8255 2634 8375 2679
rect 8255 2600 8298 2634
rect 8332 2600 8375 2634
rect 8817 3070 8860 3104
rect 8894 3070 8937 3104
rect 8817 3026 8937 3070
rect 8817 2992 8860 3026
rect 8894 2992 8937 3026
rect 8817 2948 8937 2992
rect 8817 2914 8860 2948
rect 8894 2914 8937 2948
rect 8817 2870 8937 2914
rect 8817 2836 8860 2870
rect 8894 2836 8937 2870
rect 8817 2792 8937 2836
rect 8817 2758 8860 2792
rect 8894 2758 8937 2792
rect 8817 2713 8937 2758
rect 8817 2679 8860 2713
rect 8894 2679 8937 2713
rect 8817 2634 8937 2679
rect 8255 2552 8375 2600
rect 8817 2600 8860 2634
rect 8894 2600 8937 2634
rect 8817 2552 8937 2600
rect 9247 3104 9367 3152
rect 9247 3070 9290 3104
rect 9324 3070 9367 3104
rect 9809 3104 9929 3152
rect 9247 3026 9367 3070
rect 9247 2992 9290 3026
rect 9324 2992 9367 3026
rect 9247 2948 9367 2992
rect 9247 2914 9290 2948
rect 9324 2914 9367 2948
rect 9247 2870 9367 2914
rect 9247 2836 9290 2870
rect 9324 2836 9367 2870
rect 9247 2792 9367 2836
rect 9247 2758 9290 2792
rect 9324 2758 9367 2792
rect 9247 2713 9367 2758
rect 9247 2679 9290 2713
rect 9324 2679 9367 2713
rect 9247 2634 9367 2679
rect 9247 2600 9290 2634
rect 9324 2600 9367 2634
rect 9809 3070 9852 3104
rect 9886 3070 9929 3104
rect 9809 3026 9929 3070
rect 9809 2992 9852 3026
rect 9886 2992 9929 3026
rect 9809 2948 9929 2992
rect 9809 2914 9852 2948
rect 9886 2914 9929 2948
rect 9809 2870 9929 2914
rect 9809 2836 9852 2870
rect 9886 2836 9929 2870
rect 9809 2792 9929 2836
rect 9809 2758 9852 2792
rect 9886 2758 9929 2792
rect 9809 2713 9929 2758
rect 9809 2679 9852 2713
rect 9886 2679 9929 2713
rect 9809 2634 9929 2679
rect 9247 2552 9367 2600
rect 9809 2600 9852 2634
rect 9886 2600 9929 2634
rect 9809 2552 9929 2600
rect 10239 3104 10359 3152
rect 10239 3070 10282 3104
rect 10316 3070 10359 3104
rect 10801 3104 10921 3152
rect 10239 3026 10359 3070
rect 10239 2992 10282 3026
rect 10316 2992 10359 3026
rect 10239 2948 10359 2992
rect 10239 2914 10282 2948
rect 10316 2914 10359 2948
rect 10239 2870 10359 2914
rect 10239 2836 10282 2870
rect 10316 2836 10359 2870
rect 10239 2792 10359 2836
rect 10239 2758 10282 2792
rect 10316 2758 10359 2792
rect 10239 2713 10359 2758
rect 10239 2679 10282 2713
rect 10316 2679 10359 2713
rect 10239 2634 10359 2679
rect 10239 2600 10282 2634
rect 10316 2600 10359 2634
rect 10801 3070 10844 3104
rect 10878 3070 10921 3104
rect 10801 3026 10921 3070
rect 10801 2992 10844 3026
rect 10878 2992 10921 3026
rect 10801 2948 10921 2992
rect 10801 2914 10844 2948
rect 10878 2914 10921 2948
rect 10801 2870 10921 2914
rect 10801 2836 10844 2870
rect 10878 2836 10921 2870
rect 10801 2792 10921 2836
rect 10801 2758 10844 2792
rect 10878 2758 10921 2792
rect 10801 2713 10921 2758
rect 10801 2679 10844 2713
rect 10878 2679 10921 2713
rect 10801 2634 10921 2679
rect 10239 2552 10359 2600
rect 10801 2600 10844 2634
rect 10878 2600 10921 2634
rect 10801 2552 10921 2600
rect 11231 3104 11351 3152
rect 11231 3070 11274 3104
rect 11308 3070 11351 3104
rect 11793 3104 11913 3152
rect 11231 3026 11351 3070
rect 11231 2992 11274 3026
rect 11308 2992 11351 3026
rect 11231 2948 11351 2992
rect 11231 2914 11274 2948
rect 11308 2914 11351 2948
rect 11231 2870 11351 2914
rect 11231 2836 11274 2870
rect 11308 2836 11351 2870
rect 11231 2792 11351 2836
rect 11231 2758 11274 2792
rect 11308 2758 11351 2792
rect 11231 2713 11351 2758
rect 11231 2679 11274 2713
rect 11308 2679 11351 2713
rect 11231 2634 11351 2679
rect 11231 2600 11274 2634
rect 11308 2600 11351 2634
rect 11793 3070 11836 3104
rect 11870 3070 11913 3104
rect 11793 3026 11913 3070
rect 11793 2992 11836 3026
rect 11870 2992 11913 3026
rect 11793 2948 11913 2992
rect 11793 2914 11836 2948
rect 11870 2914 11913 2948
rect 11793 2870 11913 2914
rect 11793 2836 11836 2870
rect 11870 2836 11913 2870
rect 11793 2792 11913 2836
rect 11793 2758 11836 2792
rect 11870 2758 11913 2792
rect 11793 2713 11913 2758
rect 11793 2679 11836 2713
rect 11870 2679 11913 2713
rect 11793 2634 11913 2679
rect 11231 2552 11351 2600
rect 11793 2600 11836 2634
rect 11870 2600 11913 2634
rect 11793 2552 11913 2600
rect 12223 3104 12343 3152
rect 12223 3070 12266 3104
rect 12300 3070 12343 3104
rect 12785 3104 12905 3152
rect 12223 3026 12343 3070
rect 12223 2992 12266 3026
rect 12300 2992 12343 3026
rect 12223 2948 12343 2992
rect 12223 2914 12266 2948
rect 12300 2914 12343 2948
rect 12223 2870 12343 2914
rect 12223 2836 12266 2870
rect 12300 2836 12343 2870
rect 12223 2792 12343 2836
rect 12223 2758 12266 2792
rect 12300 2758 12343 2792
rect 12223 2713 12343 2758
rect 12223 2679 12266 2713
rect 12300 2679 12343 2713
rect 12223 2634 12343 2679
rect 12223 2600 12266 2634
rect 12300 2600 12343 2634
rect 12785 3070 12828 3104
rect 12862 3070 12905 3104
rect 12785 3026 12905 3070
rect 12785 2992 12828 3026
rect 12862 2992 12905 3026
rect 12785 2948 12905 2992
rect 12785 2914 12828 2948
rect 12862 2914 12905 2948
rect 12785 2870 12905 2914
rect 12785 2836 12828 2870
rect 12862 2836 12905 2870
rect 12785 2792 12905 2836
rect 12785 2758 12828 2792
rect 12862 2758 12905 2792
rect 12785 2713 12905 2758
rect 12785 2679 12828 2713
rect 12862 2679 12905 2713
rect 12785 2634 12905 2679
rect 12223 2552 12343 2600
rect 12785 2600 12828 2634
rect 12862 2600 12905 2634
rect 12785 2552 12905 2600
rect 13215 3104 13335 3152
rect 13215 3070 13258 3104
rect 13292 3070 13335 3104
rect 13777 3104 13897 3152
rect 13215 3026 13335 3070
rect 13215 2992 13258 3026
rect 13292 2992 13335 3026
rect 13215 2948 13335 2992
rect 13215 2914 13258 2948
rect 13292 2914 13335 2948
rect 13215 2870 13335 2914
rect 13215 2836 13258 2870
rect 13292 2836 13335 2870
rect 13215 2792 13335 2836
rect 13215 2758 13258 2792
rect 13292 2758 13335 2792
rect 13215 2713 13335 2758
rect 13215 2679 13258 2713
rect 13292 2679 13335 2713
rect 13215 2634 13335 2679
rect 13215 2600 13258 2634
rect 13292 2600 13335 2634
rect 13777 3070 13820 3104
rect 13854 3070 13897 3104
rect 13777 3026 13897 3070
rect 13777 2992 13820 3026
rect 13854 2992 13897 3026
rect 13777 2948 13897 2992
rect 13777 2914 13820 2948
rect 13854 2914 13897 2948
rect 13777 2870 13897 2914
rect 13777 2836 13820 2870
rect 13854 2836 13897 2870
rect 13777 2792 13897 2836
rect 13777 2758 13820 2792
rect 13854 2758 13897 2792
rect 13777 2713 13897 2758
rect 13777 2679 13820 2713
rect 13854 2679 13897 2713
rect 13777 2634 13897 2679
rect 13215 2552 13335 2600
rect 13777 2600 13820 2634
rect 13854 2600 13897 2634
rect 13777 2552 13897 2600
rect 14135 3104 14255 3152
rect 14135 3070 14178 3104
rect 14212 3070 14255 3104
rect 14135 3026 14255 3070
rect 14135 2992 14178 3026
rect 14212 2992 14255 3026
rect 14135 2948 14255 2992
rect 14135 2914 14178 2948
rect 14212 2914 14255 2948
rect 14135 2870 14255 2914
rect 14135 2836 14178 2870
rect 14212 2836 14255 2870
rect 14135 2792 14255 2836
rect 14135 2758 14178 2792
rect 14212 2758 14255 2792
rect 14135 2713 14255 2758
rect 14135 2679 14178 2713
rect 14212 2679 14255 2713
rect 14135 2634 14255 2679
rect 14135 2600 14178 2634
rect 14212 2600 14255 2634
rect 14135 2552 14255 2600
rect 881 1504 1001 1552
rect 881 1470 924 1504
rect 958 1470 1001 1504
rect 881 1430 1001 1470
rect 881 1396 924 1430
rect 958 1396 1001 1430
rect 881 1380 1001 1396
rect 1311 1504 1431 1552
rect 1311 1470 1354 1504
rect 1388 1470 1431 1504
rect 1311 1430 1431 1470
rect 1311 1396 1354 1430
rect 1388 1396 1431 1430
rect 1311 1380 1431 1396
rect 1873 1504 1993 1552
rect 1873 1470 1916 1504
rect 1950 1470 1993 1504
rect 1873 1430 1993 1470
rect 1873 1396 1916 1430
rect 1950 1396 1993 1430
rect 1873 1380 1993 1396
rect 2303 1504 2423 1552
rect 2303 1470 2346 1504
rect 2380 1470 2423 1504
rect 2303 1430 2423 1470
rect 2303 1396 2346 1430
rect 2380 1396 2423 1430
rect 2303 1380 2423 1396
rect 2865 1504 2985 1552
rect 2865 1470 2908 1504
rect 2942 1470 2985 1504
rect 2865 1430 2985 1470
rect 2865 1396 2908 1430
rect 2942 1396 2985 1430
rect 2865 1380 2985 1396
rect 3295 1504 3415 1552
rect 3295 1470 3338 1504
rect 3372 1470 3415 1504
rect 3295 1430 3415 1470
rect 3295 1396 3338 1430
rect 3372 1396 3415 1430
rect 3295 1380 3415 1396
rect 3857 1504 3977 1552
rect 3857 1470 3900 1504
rect 3934 1470 3977 1504
rect 3857 1430 3977 1470
rect 3857 1396 3900 1430
rect 3934 1396 3977 1430
rect 3857 1380 3977 1396
rect 4287 1504 4407 1552
rect 4287 1470 4330 1504
rect 4364 1470 4407 1504
rect 4287 1430 4407 1470
rect 4287 1396 4330 1430
rect 4364 1396 4407 1430
rect 4287 1380 4407 1396
rect 4849 1504 4969 1552
rect 4849 1470 4892 1504
rect 4926 1470 4969 1504
rect 4849 1430 4969 1470
rect 4849 1396 4892 1430
rect 4926 1396 4969 1430
rect 4849 1380 4969 1396
rect 5279 1504 5399 1552
rect 5279 1470 5322 1504
rect 5356 1470 5399 1504
rect 5279 1430 5399 1470
rect 5279 1396 5322 1430
rect 5356 1396 5399 1430
rect 5279 1380 5399 1396
rect 5841 1504 5961 1552
rect 5841 1470 5884 1504
rect 5918 1470 5961 1504
rect 5841 1430 5961 1470
rect 5841 1396 5884 1430
rect 5918 1396 5961 1430
rect 5841 1380 5961 1396
rect 6271 1504 6391 1552
rect 6271 1470 6314 1504
rect 6348 1470 6391 1504
rect 6271 1430 6391 1470
rect 6271 1396 6314 1430
rect 6348 1396 6391 1430
rect 6271 1380 6391 1396
rect 6833 1504 6953 1552
rect 6833 1470 6876 1504
rect 6910 1470 6953 1504
rect 6833 1430 6953 1470
rect 6833 1396 6876 1430
rect 6910 1396 6953 1430
rect 6833 1380 6953 1396
rect 7263 1504 7383 1552
rect 7263 1470 7306 1504
rect 7340 1470 7383 1504
rect 7263 1430 7383 1470
rect 7263 1396 7306 1430
rect 7340 1396 7383 1430
rect 7263 1380 7383 1396
rect 7825 1504 7945 1552
rect 7825 1470 7868 1504
rect 7902 1470 7945 1504
rect 7825 1430 7945 1470
rect 7825 1396 7868 1430
rect 7902 1396 7945 1430
rect 7825 1380 7945 1396
rect 8255 1504 8375 1552
rect 8255 1470 8298 1504
rect 8332 1470 8375 1504
rect 8255 1430 8375 1470
rect 8255 1396 8298 1430
rect 8332 1396 8375 1430
rect 8255 1380 8375 1396
rect 8817 1504 8937 1552
rect 8817 1470 8860 1504
rect 8894 1470 8937 1504
rect 8817 1430 8937 1470
rect 8817 1396 8860 1430
rect 8894 1396 8937 1430
rect 8817 1380 8937 1396
rect 9247 1504 9367 1552
rect 9247 1470 9290 1504
rect 9324 1470 9367 1504
rect 9247 1430 9367 1470
rect 9247 1396 9290 1430
rect 9324 1396 9367 1430
rect 9247 1380 9367 1396
rect 9809 1504 9929 1552
rect 9809 1470 9852 1504
rect 9886 1470 9929 1504
rect 9809 1430 9929 1470
rect 9809 1396 9852 1430
rect 9886 1396 9929 1430
rect 9809 1380 9929 1396
rect 10239 1504 10359 1552
rect 10239 1470 10282 1504
rect 10316 1470 10359 1504
rect 10239 1430 10359 1470
rect 10239 1396 10282 1430
rect 10316 1396 10359 1430
rect 10239 1380 10359 1396
rect 10801 1504 10921 1552
rect 10801 1470 10844 1504
rect 10878 1470 10921 1504
rect 10801 1430 10921 1470
rect 10801 1396 10844 1430
rect 10878 1396 10921 1430
rect 10801 1380 10921 1396
rect 11231 1504 11351 1552
rect 11231 1470 11274 1504
rect 11308 1470 11351 1504
rect 11231 1430 11351 1470
rect 11231 1396 11274 1430
rect 11308 1396 11351 1430
rect 11231 1380 11351 1396
rect 11793 1504 11913 1552
rect 11793 1470 11836 1504
rect 11870 1470 11913 1504
rect 11793 1430 11913 1470
rect 11793 1396 11836 1430
rect 11870 1396 11913 1430
rect 11793 1380 11913 1396
rect 12223 1504 12343 1552
rect 12223 1470 12266 1504
rect 12300 1470 12343 1504
rect 12223 1430 12343 1470
rect 12223 1396 12266 1430
rect 12300 1396 12343 1430
rect 12223 1380 12343 1396
rect 12785 1504 12905 1552
rect 12785 1470 12828 1504
rect 12862 1470 12905 1504
rect 12785 1430 12905 1470
rect 12785 1396 12828 1430
rect 12862 1396 12905 1430
rect 12785 1380 12905 1396
rect 13215 1504 13335 1552
rect 13215 1470 13258 1504
rect 13292 1470 13335 1504
rect 13215 1430 13335 1470
rect 13215 1396 13258 1430
rect 13292 1396 13335 1430
rect 13215 1380 13335 1396
rect 13777 1504 13897 1552
rect 13777 1470 13820 1504
rect 13854 1470 13897 1504
rect 13777 1430 13897 1470
rect 13777 1396 13820 1430
rect 13854 1396 13897 1430
rect 13777 1380 13897 1396
rect 14135 1504 14255 1552
rect 14135 1470 14178 1504
rect 14212 1470 14255 1504
rect 14135 1430 14255 1470
rect 14135 1396 14178 1430
rect 14212 1396 14255 1430
rect 14135 1380 14255 1396
<< polycont >>
rect 924 4274 958 4308
rect 924 4200 958 4234
rect 1354 4274 1388 4308
rect 1354 4200 1388 4234
rect 1916 4274 1950 4308
rect 1916 4200 1950 4234
rect 2346 4274 2380 4308
rect 2346 4200 2380 4234
rect 2908 4274 2942 4308
rect 2908 4200 2942 4234
rect 3338 4274 3372 4308
rect 3338 4200 3372 4234
rect 3900 4274 3934 4308
rect 3900 4200 3934 4234
rect 4330 4274 4364 4308
rect 4330 4200 4364 4234
rect 4892 4274 4926 4308
rect 4892 4200 4926 4234
rect 5322 4274 5356 4308
rect 5322 4200 5356 4234
rect 5884 4274 5918 4308
rect 5884 4200 5918 4234
rect 6314 4274 6348 4308
rect 6314 4200 6348 4234
rect 6876 4274 6910 4308
rect 6876 4200 6910 4234
rect 7306 4274 7340 4308
rect 7306 4200 7340 4234
rect 7868 4274 7902 4308
rect 7868 4200 7902 4234
rect 8298 4274 8332 4308
rect 8298 4200 8332 4234
rect 8860 4274 8894 4308
rect 8860 4200 8894 4234
rect 9290 4274 9324 4308
rect 9290 4200 9324 4234
rect 9852 4274 9886 4308
rect 9852 4200 9886 4234
rect 10282 4274 10316 4308
rect 10282 4200 10316 4234
rect 10844 4274 10878 4308
rect 10844 4200 10878 4234
rect 11274 4274 11308 4308
rect 11274 4200 11308 4234
rect 11836 4274 11870 4308
rect 11836 4200 11870 4234
rect 12266 4274 12300 4308
rect 12266 4200 12300 4234
rect 12828 4274 12862 4308
rect 12828 4200 12862 4234
rect 13258 4274 13292 4308
rect 13258 4200 13292 4234
rect 13820 4274 13854 4308
rect 13820 4200 13854 4234
rect 14178 4274 14212 4308
rect 14178 4200 14212 4234
rect 924 3070 958 3104
rect 924 2992 958 3026
rect 924 2914 958 2948
rect 924 2836 958 2870
rect 924 2758 958 2792
rect 924 2679 958 2713
rect 924 2600 958 2634
rect 1354 3070 1388 3104
rect 1354 2992 1388 3026
rect 1354 2914 1388 2948
rect 1354 2836 1388 2870
rect 1354 2758 1388 2792
rect 1354 2679 1388 2713
rect 1354 2600 1388 2634
rect 1916 3070 1950 3104
rect 1916 2992 1950 3026
rect 1916 2914 1950 2948
rect 1916 2836 1950 2870
rect 1916 2758 1950 2792
rect 1916 2679 1950 2713
rect 1916 2600 1950 2634
rect 2346 3070 2380 3104
rect 2346 2992 2380 3026
rect 2346 2914 2380 2948
rect 2346 2836 2380 2870
rect 2346 2758 2380 2792
rect 2346 2679 2380 2713
rect 2346 2600 2380 2634
rect 2908 3070 2942 3104
rect 2908 2992 2942 3026
rect 2908 2914 2942 2948
rect 2908 2836 2942 2870
rect 2908 2758 2942 2792
rect 2908 2679 2942 2713
rect 2908 2600 2942 2634
rect 3338 3070 3372 3104
rect 3338 2992 3372 3026
rect 3338 2914 3372 2948
rect 3338 2836 3372 2870
rect 3338 2758 3372 2792
rect 3338 2679 3372 2713
rect 3338 2600 3372 2634
rect 3900 3070 3934 3104
rect 3900 2992 3934 3026
rect 3900 2914 3934 2948
rect 3900 2836 3934 2870
rect 3900 2758 3934 2792
rect 3900 2679 3934 2713
rect 3900 2600 3934 2634
rect 4330 3070 4364 3104
rect 4330 2992 4364 3026
rect 4330 2914 4364 2948
rect 4330 2836 4364 2870
rect 4330 2758 4364 2792
rect 4330 2679 4364 2713
rect 4330 2600 4364 2634
rect 4892 3070 4926 3104
rect 4892 2992 4926 3026
rect 4892 2914 4926 2948
rect 4892 2836 4926 2870
rect 4892 2758 4926 2792
rect 4892 2679 4926 2713
rect 4892 2600 4926 2634
rect 5322 3070 5356 3104
rect 5322 2992 5356 3026
rect 5322 2914 5356 2948
rect 5322 2836 5356 2870
rect 5322 2758 5356 2792
rect 5322 2679 5356 2713
rect 5322 2600 5356 2634
rect 5884 3070 5918 3104
rect 5884 2992 5918 3026
rect 5884 2914 5918 2948
rect 5884 2836 5918 2870
rect 5884 2758 5918 2792
rect 5884 2679 5918 2713
rect 5884 2600 5918 2634
rect 6314 3070 6348 3104
rect 6314 2992 6348 3026
rect 6314 2914 6348 2948
rect 6314 2836 6348 2870
rect 6314 2758 6348 2792
rect 6314 2679 6348 2713
rect 6314 2600 6348 2634
rect 6876 3070 6910 3104
rect 6876 2992 6910 3026
rect 6876 2914 6910 2948
rect 6876 2836 6910 2870
rect 6876 2758 6910 2792
rect 6876 2679 6910 2713
rect 6876 2600 6910 2634
rect 7306 3070 7340 3104
rect 7306 2992 7340 3026
rect 7306 2914 7340 2948
rect 7306 2836 7340 2870
rect 7306 2758 7340 2792
rect 7306 2679 7340 2713
rect 7306 2600 7340 2634
rect 7868 3070 7902 3104
rect 7868 2992 7902 3026
rect 7868 2914 7902 2948
rect 7868 2836 7902 2870
rect 7868 2758 7902 2792
rect 7868 2679 7902 2713
rect 7868 2600 7902 2634
rect 8298 3070 8332 3104
rect 8298 2992 8332 3026
rect 8298 2914 8332 2948
rect 8298 2836 8332 2870
rect 8298 2758 8332 2792
rect 8298 2679 8332 2713
rect 8298 2600 8332 2634
rect 8860 3070 8894 3104
rect 8860 2992 8894 3026
rect 8860 2914 8894 2948
rect 8860 2836 8894 2870
rect 8860 2758 8894 2792
rect 8860 2679 8894 2713
rect 8860 2600 8894 2634
rect 9290 3070 9324 3104
rect 9290 2992 9324 3026
rect 9290 2914 9324 2948
rect 9290 2836 9324 2870
rect 9290 2758 9324 2792
rect 9290 2679 9324 2713
rect 9290 2600 9324 2634
rect 9852 3070 9886 3104
rect 9852 2992 9886 3026
rect 9852 2914 9886 2948
rect 9852 2836 9886 2870
rect 9852 2758 9886 2792
rect 9852 2679 9886 2713
rect 9852 2600 9886 2634
rect 10282 3070 10316 3104
rect 10282 2992 10316 3026
rect 10282 2914 10316 2948
rect 10282 2836 10316 2870
rect 10282 2758 10316 2792
rect 10282 2679 10316 2713
rect 10282 2600 10316 2634
rect 10844 3070 10878 3104
rect 10844 2992 10878 3026
rect 10844 2914 10878 2948
rect 10844 2836 10878 2870
rect 10844 2758 10878 2792
rect 10844 2679 10878 2713
rect 10844 2600 10878 2634
rect 11274 3070 11308 3104
rect 11274 2992 11308 3026
rect 11274 2914 11308 2948
rect 11274 2836 11308 2870
rect 11274 2758 11308 2792
rect 11274 2679 11308 2713
rect 11274 2600 11308 2634
rect 11836 3070 11870 3104
rect 11836 2992 11870 3026
rect 11836 2914 11870 2948
rect 11836 2836 11870 2870
rect 11836 2758 11870 2792
rect 11836 2679 11870 2713
rect 11836 2600 11870 2634
rect 12266 3070 12300 3104
rect 12266 2992 12300 3026
rect 12266 2914 12300 2948
rect 12266 2836 12300 2870
rect 12266 2758 12300 2792
rect 12266 2679 12300 2713
rect 12266 2600 12300 2634
rect 12828 3070 12862 3104
rect 12828 2992 12862 3026
rect 12828 2914 12862 2948
rect 12828 2836 12862 2870
rect 12828 2758 12862 2792
rect 12828 2679 12862 2713
rect 12828 2600 12862 2634
rect 13258 3070 13292 3104
rect 13258 2992 13292 3026
rect 13258 2914 13292 2948
rect 13258 2836 13292 2870
rect 13258 2758 13292 2792
rect 13258 2679 13292 2713
rect 13258 2600 13292 2634
rect 13820 3070 13854 3104
rect 13820 2992 13854 3026
rect 13820 2914 13854 2948
rect 13820 2836 13854 2870
rect 13820 2758 13854 2792
rect 13820 2679 13854 2713
rect 13820 2600 13854 2634
rect 14178 3070 14212 3104
rect 14178 2992 14212 3026
rect 14178 2914 14212 2948
rect 14178 2836 14212 2870
rect 14178 2758 14212 2792
rect 14178 2679 14212 2713
rect 14178 2600 14212 2634
rect 924 1470 958 1504
rect 924 1396 958 1430
rect 1354 1470 1388 1504
rect 1354 1396 1388 1430
rect 1916 1470 1950 1504
rect 1916 1396 1950 1430
rect 2346 1470 2380 1504
rect 2346 1396 2380 1430
rect 2908 1470 2942 1504
rect 2908 1396 2942 1430
rect 3338 1470 3372 1504
rect 3338 1396 3372 1430
rect 3900 1470 3934 1504
rect 3900 1396 3934 1430
rect 4330 1470 4364 1504
rect 4330 1396 4364 1430
rect 4892 1470 4926 1504
rect 4892 1396 4926 1430
rect 5322 1470 5356 1504
rect 5322 1396 5356 1430
rect 5884 1470 5918 1504
rect 5884 1396 5918 1430
rect 6314 1470 6348 1504
rect 6314 1396 6348 1430
rect 6876 1470 6910 1504
rect 6876 1396 6910 1430
rect 7306 1470 7340 1504
rect 7306 1396 7340 1430
rect 7868 1470 7902 1504
rect 7868 1396 7902 1430
rect 8298 1470 8332 1504
rect 8298 1396 8332 1430
rect 8860 1470 8894 1504
rect 8860 1396 8894 1430
rect 9290 1470 9324 1504
rect 9290 1396 9324 1430
rect 9852 1470 9886 1504
rect 9852 1396 9886 1430
rect 10282 1470 10316 1504
rect 10282 1396 10316 1430
rect 10844 1470 10878 1504
rect 10844 1396 10878 1430
rect 11274 1470 11308 1504
rect 11274 1396 11308 1430
rect 11836 1470 11870 1504
rect 11836 1396 11870 1430
rect 12266 1470 12300 1504
rect 12266 1396 12300 1430
rect 12828 1470 12862 1504
rect 12828 1396 12862 1430
rect 13258 1470 13292 1504
rect 13258 1396 13292 1430
rect 13820 1470 13854 1504
rect 13820 1396 13854 1430
rect 14178 1470 14212 1504
rect 14178 1396 14212 1430
<< locali >>
rect 100 5118 329 5148
rect 14807 5118 15013 5150
rect 100 5111 15013 5118
rect 100 5083 361 5111
rect 15 5082 361 5083
rect 395 5082 434 5111
rect 468 5082 507 5111
rect 541 5082 580 5111
rect 614 5082 653 5111
rect 687 5082 726 5111
rect 760 5082 799 5111
rect 833 5082 872 5111
rect 906 5082 945 5111
rect 979 5082 1018 5111
rect 1052 5082 1091 5111
rect 1125 5082 1164 5111
rect 1198 5082 1237 5111
rect 1271 5082 1310 5111
rect 1344 5082 1383 5111
rect 1417 5082 1456 5111
rect 1490 5082 1529 5111
rect 1563 5082 1602 5111
rect 1636 5082 1675 5111
rect 1709 5082 1748 5111
rect 1782 5082 1821 5111
rect 1855 5082 1894 5111
rect 1928 5082 1967 5111
rect 2001 5082 2040 5111
rect 2074 5082 2113 5111
rect 2147 5082 2186 5111
rect 2220 5082 2259 5111
rect 2293 5082 2332 5111
rect 2366 5082 2405 5111
rect 2439 5082 2478 5111
rect 2512 5082 2551 5111
rect 2585 5082 2624 5111
rect 2658 5082 2697 5111
rect 2731 5082 2770 5111
rect 2804 5082 2843 5111
rect 2877 5082 2916 5111
rect 2950 5082 2989 5111
rect 3023 5082 3062 5111
rect 3096 5082 3135 5111
rect 3169 5082 3208 5111
rect 3242 5082 3281 5111
rect 3315 5082 3354 5111
rect 3388 5082 3427 5111
rect 3461 5082 3500 5111
rect 3534 5082 3573 5111
rect 3607 5082 3646 5111
rect 3680 5082 3719 5111
rect 3753 5082 3792 5111
rect 3826 5082 3865 5111
rect 3899 5082 3938 5111
rect 3972 5082 4011 5111
rect 4045 5082 4084 5111
rect 4118 5082 4157 5111
rect 4191 5082 4229 5111
rect 4263 5082 4301 5111
rect 4335 5082 4373 5111
rect 4407 5082 4445 5111
rect 4479 5082 4517 5111
rect 4551 5082 4589 5111
rect 4623 5082 4661 5111
rect 4695 5082 4733 5111
rect 4767 5082 4805 5111
rect 4839 5082 4877 5111
rect 4911 5082 4949 5111
rect 4983 5082 5021 5111
rect 5055 5082 5093 5111
rect 5127 5082 5165 5111
rect 5199 5082 5237 5111
rect 5271 5082 5309 5111
rect 5343 5082 5381 5111
rect 5415 5082 5453 5111
rect 5487 5082 5525 5111
rect 5559 5082 5597 5111
rect 5631 5082 5669 5111
rect 5703 5082 5741 5111
rect 5775 5082 5813 5111
rect 5847 5082 5885 5111
rect 5919 5082 5957 5111
rect 5991 5082 6029 5111
rect 6063 5082 6101 5111
rect 6135 5082 6173 5111
rect 6207 5082 6245 5111
rect 6279 5082 6317 5111
rect 6351 5082 6389 5111
rect 6423 5082 6461 5111
rect 6495 5082 6533 5111
rect 6567 5082 6605 5111
rect 6639 5082 6677 5111
rect 6711 5082 6749 5111
rect 6783 5082 6821 5111
rect 6855 5082 6893 5111
rect 6927 5082 6965 5111
rect 6999 5082 7037 5111
rect 7071 5082 7109 5111
rect 7143 5082 7181 5111
rect 7215 5082 7253 5111
rect 7287 5082 7325 5111
rect 7359 5082 7397 5111
rect 7431 5082 7469 5111
rect 7503 5082 7541 5111
rect 7575 5082 7613 5111
rect 7647 5082 7685 5111
rect 7719 5082 7757 5111
rect 7791 5082 7829 5111
rect 7863 5082 7901 5111
rect 7935 5082 7973 5111
rect 8007 5082 8045 5111
rect 8079 5082 8117 5111
rect 8151 5082 8189 5111
rect 8223 5082 8261 5111
rect 8295 5082 8333 5111
rect 8367 5082 8405 5111
rect 8439 5082 8477 5111
rect 8511 5082 8549 5111
rect 8583 5082 8621 5111
rect 8655 5082 8693 5111
rect 8727 5082 8765 5111
rect 8799 5082 8837 5111
rect 8871 5082 8909 5111
rect 8943 5082 8981 5111
rect 9015 5082 9053 5111
rect 9087 5082 9125 5111
rect 9159 5082 9197 5111
rect 9231 5082 9269 5111
rect 9303 5082 9341 5111
rect 9375 5082 9413 5111
rect 9447 5082 9485 5111
rect 9519 5082 9557 5111
rect 9591 5082 9629 5111
rect 9663 5082 9701 5111
rect 9735 5082 9773 5111
rect 9807 5082 9845 5111
rect 9879 5082 9917 5111
rect 9951 5082 9989 5111
rect 10023 5082 10061 5111
rect 10095 5082 10133 5111
rect 10167 5082 10205 5111
rect 10239 5082 10277 5111
rect 10311 5082 10349 5111
rect 10383 5082 10421 5111
rect 10455 5082 10493 5111
rect 10527 5082 10565 5111
rect 10599 5082 10637 5111
rect 10671 5082 10709 5111
rect 10743 5082 10781 5111
rect 10815 5082 10853 5111
rect 10887 5082 10925 5111
rect 10959 5082 10997 5111
rect 11031 5082 11069 5111
rect 11103 5082 11141 5111
rect 11175 5082 11213 5111
rect 11247 5082 11285 5111
rect 11319 5082 11357 5111
rect 11391 5082 11429 5111
rect 11463 5082 11501 5111
rect 11535 5082 11573 5111
rect 11607 5082 11645 5111
rect 11679 5082 11717 5111
rect 11751 5082 11789 5111
rect 11823 5082 11861 5111
rect 11895 5082 11933 5111
rect 11967 5082 12005 5111
rect 12039 5082 12077 5111
rect 12111 5082 12149 5111
rect 12183 5082 12221 5111
rect 12255 5082 12293 5111
rect 12327 5082 12365 5111
rect 12399 5082 12437 5111
rect 12471 5082 12509 5111
rect 12543 5082 12581 5111
rect 12615 5082 12653 5111
rect 12687 5082 12725 5111
rect 12759 5082 12797 5111
rect 12831 5082 12869 5111
rect 12903 5082 12941 5111
rect 12975 5082 13013 5111
rect 13047 5082 13085 5111
rect 13119 5082 13157 5111
rect 13191 5082 13229 5111
rect 13263 5082 13301 5111
rect 13335 5082 13373 5111
rect 13407 5082 13445 5111
rect 13479 5082 13517 5111
rect 13551 5082 13589 5111
rect 13623 5082 13661 5111
rect 13695 5082 13733 5111
rect 13767 5082 13805 5111
rect 13839 5082 13877 5111
rect 13911 5082 13949 5111
rect 13983 5082 14021 5111
rect 14055 5082 14093 5111
rect 14127 5082 14165 5111
rect 14199 5082 14237 5111
rect 14271 5082 14309 5111
rect 14343 5082 14381 5111
rect 14415 5082 14453 5111
rect 14487 5082 14525 5111
rect 14559 5082 14597 5111
rect 14631 5082 14669 5111
rect 14703 5082 14741 5111
rect 14775 5082 15013 5111
rect 15 5048 252 5082
rect 286 5048 320 5082
rect 354 5077 361 5082
rect 422 5077 434 5082
rect 490 5077 507 5082
rect 558 5077 580 5082
rect 626 5077 653 5082
rect 694 5077 726 5082
rect 354 5048 388 5077
rect 422 5048 456 5077
rect 490 5048 524 5077
rect 558 5048 592 5077
rect 626 5048 660 5077
rect 694 5048 728 5077
rect 762 5048 796 5082
rect 833 5077 864 5082
rect 906 5077 932 5082
rect 979 5077 1000 5082
rect 1052 5077 1068 5082
rect 1125 5077 1136 5082
rect 1198 5077 1204 5082
rect 1271 5077 1272 5082
rect 830 5048 864 5077
rect 898 5048 932 5077
rect 966 5048 1000 5077
rect 1034 5048 1068 5077
rect 1102 5048 1136 5077
rect 1170 5048 1204 5077
rect 1238 5048 1272 5077
rect 1306 5077 1310 5082
rect 1374 5077 1383 5082
rect 1442 5077 1456 5082
rect 1510 5077 1529 5082
rect 1578 5077 1602 5082
rect 1646 5077 1675 5082
rect 1306 5048 1340 5077
rect 1374 5048 1408 5077
rect 1442 5048 1476 5077
rect 1510 5048 1544 5077
rect 1578 5048 1612 5077
rect 1646 5048 1680 5077
rect 1714 5048 1748 5082
rect 1782 5048 1816 5082
rect 1855 5077 1884 5082
rect 1928 5077 1952 5082
rect 2001 5077 2020 5082
rect 2074 5077 2088 5082
rect 2147 5077 2156 5082
rect 2220 5077 2224 5082
rect 1850 5048 1884 5077
rect 1918 5048 1952 5077
rect 1986 5048 2020 5077
rect 2054 5048 2088 5077
rect 2122 5048 2156 5077
rect 2190 5048 2224 5077
rect 2258 5077 2259 5082
rect 2326 5077 2332 5082
rect 2394 5077 2405 5082
rect 2462 5077 2478 5082
rect 2530 5077 2551 5082
rect 2598 5077 2624 5082
rect 2666 5077 2697 5082
rect 2258 5048 2292 5077
rect 2326 5048 2360 5077
rect 2394 5048 2428 5077
rect 2462 5048 2496 5077
rect 2530 5048 2564 5077
rect 2598 5048 2632 5077
rect 2666 5048 2700 5077
rect 2734 5048 2768 5082
rect 2804 5077 2836 5082
rect 2877 5077 2904 5082
rect 2950 5077 2972 5082
rect 3023 5077 3040 5082
rect 3096 5077 3108 5082
rect 3169 5077 3176 5082
rect 3242 5077 3244 5082
rect 2802 5048 2836 5077
rect 2870 5048 2904 5077
rect 2938 5048 2972 5077
rect 3006 5048 3040 5077
rect 3074 5048 3108 5077
rect 3142 5048 3176 5077
rect 3210 5048 3244 5077
rect 3278 5077 3281 5082
rect 3346 5077 3354 5082
rect 3414 5077 3427 5082
rect 3482 5077 3500 5082
rect 3550 5077 3573 5082
rect 3618 5077 3646 5082
rect 3686 5077 3719 5082
rect 3278 5048 3312 5077
rect 3346 5048 3380 5077
rect 3414 5048 3448 5077
rect 3482 5048 3516 5077
rect 3550 5048 3584 5077
rect 3618 5048 3652 5077
rect 3686 5048 3720 5077
rect 3754 5048 3788 5082
rect 3826 5077 3856 5082
rect 3899 5077 3924 5082
rect 3972 5077 3992 5082
rect 4045 5077 4060 5082
rect 4118 5077 4128 5082
rect 4191 5077 4196 5082
rect 4263 5077 4264 5082
rect 3822 5048 3856 5077
rect 3890 5048 3924 5077
rect 3958 5048 3992 5077
rect 4026 5048 4060 5077
rect 4094 5048 4128 5077
rect 4162 5048 4196 5077
rect 4230 5048 4264 5077
rect 4298 5077 4301 5082
rect 4366 5077 4373 5082
rect 4434 5077 4445 5082
rect 4502 5077 4517 5082
rect 4570 5077 4589 5082
rect 4638 5077 4661 5082
rect 4706 5077 4733 5082
rect 4774 5077 4805 5082
rect 4298 5048 4332 5077
rect 4366 5048 4400 5077
rect 4434 5048 4468 5077
rect 4502 5048 4536 5077
rect 4570 5048 4604 5077
rect 4638 5048 4672 5077
rect 4706 5048 4740 5077
rect 4774 5048 4808 5077
rect 4842 5048 4876 5082
rect 4911 5077 4944 5082
rect 4983 5077 5012 5082
rect 5055 5077 5080 5082
rect 5127 5077 5148 5082
rect 5199 5077 5216 5082
rect 5271 5077 5284 5082
rect 5343 5077 5352 5082
rect 5415 5077 5420 5082
rect 5487 5077 5488 5082
rect 4910 5048 4944 5077
rect 4978 5048 5012 5077
rect 5046 5048 5080 5077
rect 5114 5048 5148 5077
rect 5182 5048 5216 5077
rect 5250 5048 5284 5077
rect 5318 5048 5352 5077
rect 5386 5048 5420 5077
rect 5454 5048 5488 5077
rect 5522 5077 5525 5082
rect 5590 5077 5597 5082
rect 5658 5077 5669 5082
rect 5726 5077 5741 5082
rect 5794 5077 5813 5082
rect 5862 5077 5885 5082
rect 5930 5077 5957 5082
rect 5998 5077 6029 5082
rect 5522 5048 5556 5077
rect 5590 5048 5624 5077
rect 5658 5048 5692 5077
rect 5726 5048 5760 5077
rect 5794 5048 5828 5077
rect 5862 5048 5896 5077
rect 5930 5048 5964 5077
rect 5998 5048 6032 5077
rect 6066 5048 6100 5082
rect 6135 5077 6168 5082
rect 6207 5077 6236 5082
rect 6279 5077 6304 5082
rect 6351 5077 6372 5082
rect 6423 5077 6440 5082
rect 6495 5077 6508 5082
rect 6567 5077 6576 5082
rect 6639 5077 6644 5082
rect 6711 5077 6712 5082
rect 6134 5048 6168 5077
rect 6202 5048 6236 5077
rect 6270 5048 6304 5077
rect 6338 5048 6372 5077
rect 6406 5048 6440 5077
rect 6474 5048 6508 5077
rect 6542 5048 6576 5077
rect 6610 5048 6644 5077
rect 6678 5048 6712 5077
rect 6746 5077 6749 5082
rect 6814 5077 6821 5082
rect 6882 5077 6893 5082
rect 6950 5077 6965 5082
rect 7018 5077 7037 5082
rect 7086 5077 7109 5082
rect 7154 5077 7181 5082
rect 7222 5077 7253 5082
rect 6746 5048 6780 5077
rect 6814 5048 6848 5077
rect 6882 5048 6916 5077
rect 6950 5048 6984 5077
rect 7018 5048 7052 5077
rect 7086 5048 7120 5077
rect 7154 5048 7188 5077
rect 7222 5048 7256 5077
rect 7290 5048 7324 5082
rect 7359 5077 7392 5082
rect 7431 5077 7460 5082
rect 7503 5077 7528 5082
rect 7575 5077 7596 5082
rect 7647 5077 7664 5082
rect 7719 5077 7732 5082
rect 7791 5077 7800 5082
rect 7863 5077 7868 5082
rect 7935 5077 7936 5082
rect 7358 5048 7392 5077
rect 7426 5048 7460 5077
rect 7494 5048 7528 5077
rect 7562 5048 7596 5077
rect 7630 5048 7664 5077
rect 7698 5048 7732 5077
rect 7766 5048 7800 5077
rect 7834 5048 7868 5077
rect 7902 5048 7936 5077
rect 7970 5077 7973 5082
rect 8038 5077 8045 5082
rect 8106 5077 8117 5082
rect 8174 5077 8189 5082
rect 8242 5077 8261 5082
rect 8310 5077 8333 5082
rect 8378 5077 8405 5082
rect 8446 5077 8477 5082
rect 7970 5048 8004 5077
rect 8038 5048 8072 5077
rect 8106 5048 8140 5077
rect 8174 5048 8208 5077
rect 8242 5048 8276 5077
rect 8310 5048 8344 5077
rect 8378 5048 8412 5077
rect 8446 5048 8480 5077
rect 8514 5048 8548 5082
rect 8583 5077 8616 5082
rect 8655 5077 8684 5082
rect 8727 5077 8752 5082
rect 8799 5077 8820 5082
rect 8871 5077 8888 5082
rect 8943 5077 8956 5082
rect 9015 5077 9024 5082
rect 9087 5077 9092 5082
rect 9159 5077 9160 5082
rect 8582 5048 8616 5077
rect 8650 5048 8684 5077
rect 8718 5048 8752 5077
rect 8786 5048 8820 5077
rect 8854 5048 8888 5077
rect 8922 5048 8956 5077
rect 8990 5048 9024 5077
rect 9058 5048 9092 5077
rect 9126 5048 9160 5077
rect 9194 5077 9197 5082
rect 9262 5077 9269 5082
rect 9330 5077 9341 5082
rect 9398 5077 9413 5082
rect 9466 5077 9485 5082
rect 9534 5077 9557 5082
rect 9602 5077 9629 5082
rect 9670 5077 9701 5082
rect 9194 5048 9228 5077
rect 9262 5048 9296 5077
rect 9330 5048 9364 5077
rect 9398 5048 9432 5077
rect 9466 5048 9500 5077
rect 9534 5048 9568 5077
rect 9602 5048 9636 5077
rect 9670 5048 9704 5077
rect 9738 5048 9772 5082
rect 9807 5077 9840 5082
rect 9879 5077 9908 5082
rect 9951 5077 9976 5082
rect 10023 5077 10044 5082
rect 10095 5077 10112 5082
rect 10167 5077 10180 5082
rect 10239 5077 10248 5082
rect 10311 5077 10316 5082
rect 10383 5077 10384 5082
rect 9806 5048 9840 5077
rect 9874 5048 9908 5077
rect 9942 5048 9976 5077
rect 10010 5048 10044 5077
rect 10078 5048 10112 5077
rect 10146 5048 10180 5077
rect 10214 5048 10248 5077
rect 10282 5048 10316 5077
rect 10350 5048 10384 5077
rect 10418 5077 10421 5082
rect 10486 5077 10493 5082
rect 10554 5077 10565 5082
rect 10622 5077 10637 5082
rect 10690 5077 10709 5082
rect 10758 5077 10781 5082
rect 10826 5077 10853 5082
rect 10894 5077 10925 5082
rect 10418 5048 10452 5077
rect 10486 5048 10520 5077
rect 10554 5048 10588 5077
rect 10622 5048 10656 5077
rect 10690 5048 10724 5077
rect 10758 5048 10792 5077
rect 10826 5048 10860 5077
rect 10894 5048 10928 5077
rect 10962 5048 10996 5082
rect 11031 5077 11064 5082
rect 11103 5077 11132 5082
rect 11175 5077 11200 5082
rect 11247 5077 11268 5082
rect 11319 5077 11336 5082
rect 11391 5077 11404 5082
rect 11463 5077 11472 5082
rect 11535 5077 11540 5082
rect 11607 5077 11608 5082
rect 11030 5048 11064 5077
rect 11098 5048 11132 5077
rect 11166 5048 11200 5077
rect 11234 5048 11268 5077
rect 11302 5048 11336 5077
rect 11370 5048 11404 5077
rect 11438 5048 11472 5077
rect 11506 5048 11540 5077
rect 11574 5048 11608 5077
rect 11642 5077 11645 5082
rect 11710 5077 11717 5082
rect 11778 5077 11789 5082
rect 11846 5077 11861 5082
rect 11914 5077 11933 5082
rect 11982 5077 12005 5082
rect 12050 5077 12077 5082
rect 12118 5077 12149 5082
rect 11642 5048 11676 5077
rect 11710 5048 11744 5077
rect 11778 5048 11812 5077
rect 11846 5048 11880 5077
rect 11914 5048 11948 5077
rect 11982 5048 12016 5077
rect 12050 5048 12084 5077
rect 12118 5048 12152 5077
rect 12186 5048 12220 5082
rect 12255 5077 12288 5082
rect 12327 5077 12356 5082
rect 12399 5077 12424 5082
rect 12471 5077 12492 5082
rect 12543 5077 12560 5082
rect 12615 5077 12628 5082
rect 12687 5077 12696 5082
rect 12759 5077 12764 5082
rect 12831 5077 12832 5082
rect 12254 5048 12288 5077
rect 12322 5048 12356 5077
rect 12390 5048 12424 5077
rect 12458 5048 12492 5077
rect 12526 5048 12560 5077
rect 12594 5048 12628 5077
rect 12662 5048 12696 5077
rect 12730 5048 12764 5077
rect 12798 5048 12832 5077
rect 12866 5077 12869 5082
rect 12934 5077 12941 5082
rect 13002 5077 13013 5082
rect 13070 5077 13085 5082
rect 13138 5077 13157 5082
rect 13206 5077 13229 5082
rect 13274 5077 13301 5082
rect 13342 5077 13373 5082
rect 12866 5048 12900 5077
rect 12934 5048 12968 5077
rect 13002 5048 13036 5077
rect 13070 5048 13104 5077
rect 13138 5048 13172 5077
rect 13206 5048 13240 5077
rect 13274 5048 13308 5077
rect 13342 5048 13376 5077
rect 13410 5048 13444 5082
rect 13479 5077 13512 5082
rect 13551 5077 13580 5082
rect 13623 5077 13648 5082
rect 13695 5077 13716 5082
rect 13767 5077 13784 5082
rect 13839 5077 13852 5082
rect 13911 5077 13920 5082
rect 13983 5077 13988 5082
rect 14055 5077 14056 5082
rect 13478 5048 13512 5077
rect 13546 5048 13580 5077
rect 13614 5048 13648 5077
rect 13682 5048 13716 5077
rect 13750 5048 13784 5077
rect 13818 5048 13852 5077
rect 13886 5048 13920 5077
rect 13954 5048 13988 5077
rect 14022 5048 14056 5077
rect 14090 5077 14093 5082
rect 14158 5077 14165 5082
rect 14226 5077 14237 5082
rect 14294 5077 14309 5082
rect 14362 5077 14381 5082
rect 14430 5077 14453 5082
rect 14498 5077 14525 5082
rect 14566 5077 14597 5082
rect 14090 5048 14124 5077
rect 14158 5048 14192 5077
rect 14226 5048 14260 5077
rect 14294 5048 14328 5077
rect 14362 5048 14396 5077
rect 14430 5048 14464 5077
rect 14498 5048 14532 5077
rect 14566 5048 14600 5077
rect 14634 5048 14668 5082
rect 14703 5077 14736 5082
rect 14775 5077 14804 5082
rect 14702 5048 14736 5077
rect 14770 5048 14804 5077
rect 14838 5048 14872 5082
rect 14906 5062 15013 5082
rect 14906 5048 14907 5062
rect 15 5045 14907 5048
rect 15 331 125 5045
rect 231 5035 14907 5045
rect 231 5029 361 5035
rect 231 5000 269 5029
rect 303 5001 361 5029
rect 395 5001 434 5035
rect 468 5001 507 5035
rect 541 5001 580 5035
rect 614 5001 653 5035
rect 687 5001 726 5035
rect 760 5001 799 5035
rect 833 5001 872 5035
rect 906 5001 945 5035
rect 979 5001 1018 5035
rect 1052 5001 1091 5035
rect 1125 5001 1164 5035
rect 1198 5001 1237 5035
rect 1271 5001 1310 5035
rect 1344 5001 1383 5035
rect 1417 5001 1456 5035
rect 1490 5001 1529 5035
rect 1563 5001 1602 5035
rect 1636 5001 1675 5035
rect 1709 5001 1748 5035
rect 1782 5001 1821 5035
rect 1855 5001 1894 5035
rect 1928 5001 1967 5035
rect 2001 5001 2040 5035
rect 2074 5001 2113 5035
rect 2147 5001 2186 5035
rect 2220 5001 2259 5035
rect 2293 5001 2332 5035
rect 2366 5001 2405 5035
rect 2439 5001 2478 5035
rect 2512 5001 2551 5035
rect 2585 5001 2624 5035
rect 2658 5001 2697 5035
rect 2731 5001 2770 5035
rect 2804 5001 2843 5035
rect 2877 5001 2916 5035
rect 2950 5001 2989 5035
rect 3023 5001 3062 5035
rect 3096 5001 3135 5035
rect 3169 5001 3208 5035
rect 3242 5001 3281 5035
rect 3315 5001 3354 5035
rect 3388 5001 3427 5035
rect 3461 5001 3500 5035
rect 3534 5001 3573 5035
rect 3607 5001 3646 5035
rect 3680 5001 3719 5035
rect 3753 5001 3792 5035
rect 3826 5001 3865 5035
rect 3899 5001 3938 5035
rect 3972 5001 4011 5035
rect 4045 5001 4084 5035
rect 4118 5001 4157 5035
rect 4191 5001 4229 5035
rect 4263 5001 4301 5035
rect 4335 5001 4373 5035
rect 4407 5001 4445 5035
rect 4479 5001 4517 5035
rect 4551 5001 4589 5035
rect 4623 5001 4661 5035
rect 4695 5001 4733 5035
rect 4767 5001 4805 5035
rect 4839 5001 4877 5035
rect 4911 5001 4949 5035
rect 4983 5001 5021 5035
rect 5055 5001 5093 5035
rect 5127 5001 5165 5035
rect 5199 5001 5237 5035
rect 5271 5001 5309 5035
rect 5343 5001 5381 5035
rect 5415 5001 5453 5035
rect 5487 5001 5525 5035
rect 5559 5001 5597 5035
rect 5631 5001 5669 5035
rect 5703 5001 5741 5035
rect 5775 5001 5813 5035
rect 5847 5001 5885 5035
rect 5919 5001 5957 5035
rect 5991 5001 6029 5035
rect 6063 5001 6101 5035
rect 6135 5001 6173 5035
rect 6207 5001 6245 5035
rect 6279 5001 6317 5035
rect 6351 5001 6389 5035
rect 6423 5001 6461 5035
rect 6495 5001 6533 5035
rect 6567 5001 6605 5035
rect 6639 5001 6677 5035
rect 6711 5001 6749 5035
rect 6783 5001 6821 5035
rect 6855 5001 6893 5035
rect 6927 5001 6965 5035
rect 6999 5001 7037 5035
rect 7071 5001 7109 5035
rect 7143 5001 7181 5035
rect 7215 5001 7253 5035
rect 7287 5001 7325 5035
rect 7359 5001 7397 5035
rect 7431 5001 7469 5035
rect 7503 5001 7541 5035
rect 7575 5001 7613 5035
rect 7647 5001 7685 5035
rect 7719 5001 7757 5035
rect 7791 5001 7829 5035
rect 7863 5001 7901 5035
rect 7935 5001 7973 5035
rect 8007 5001 8045 5035
rect 8079 5001 8117 5035
rect 8151 5001 8189 5035
rect 8223 5001 8261 5035
rect 8295 5001 8333 5035
rect 8367 5001 8405 5035
rect 8439 5001 8477 5035
rect 8511 5001 8549 5035
rect 8583 5001 8621 5035
rect 8655 5001 8693 5035
rect 8727 5001 8765 5035
rect 8799 5001 8837 5035
rect 8871 5001 8909 5035
rect 8943 5001 8981 5035
rect 9015 5001 9053 5035
rect 9087 5001 9125 5035
rect 9159 5001 9197 5035
rect 9231 5001 9269 5035
rect 9303 5001 9341 5035
rect 9375 5001 9413 5035
rect 9447 5001 9485 5035
rect 9519 5001 9557 5035
rect 9591 5001 9629 5035
rect 9663 5001 9701 5035
rect 9735 5001 9773 5035
rect 9807 5001 9845 5035
rect 9879 5001 9917 5035
rect 9951 5001 9989 5035
rect 10023 5001 10061 5035
rect 10095 5001 10133 5035
rect 10167 5001 10205 5035
rect 10239 5001 10277 5035
rect 10311 5001 10349 5035
rect 10383 5001 10421 5035
rect 10455 5001 10493 5035
rect 10527 5001 10565 5035
rect 10599 5001 10637 5035
rect 10671 5001 10709 5035
rect 10743 5001 10781 5035
rect 10815 5001 10853 5035
rect 10887 5001 10925 5035
rect 10959 5001 10997 5035
rect 11031 5001 11069 5035
rect 11103 5001 11141 5035
rect 11175 5001 11213 5035
rect 11247 5001 11285 5035
rect 11319 5001 11357 5035
rect 11391 5001 11429 5035
rect 11463 5001 11501 5035
rect 11535 5001 11573 5035
rect 11607 5001 11645 5035
rect 11679 5001 11717 5035
rect 11751 5001 11789 5035
rect 11823 5001 11861 5035
rect 11895 5001 11933 5035
rect 11967 5001 12005 5035
rect 12039 5001 12077 5035
rect 12111 5001 12149 5035
rect 12183 5001 12221 5035
rect 12255 5001 12293 5035
rect 12327 5001 12365 5035
rect 12399 5001 12437 5035
rect 12471 5001 12509 5035
rect 12543 5001 12581 5035
rect 12615 5001 12653 5035
rect 12687 5001 12725 5035
rect 12759 5001 12797 5035
rect 12831 5001 12869 5035
rect 12903 5001 12941 5035
rect 12975 5001 13013 5035
rect 13047 5001 13085 5035
rect 13119 5001 13157 5035
rect 13191 5001 13229 5035
rect 13263 5001 13301 5035
rect 13335 5001 13373 5035
rect 13407 5001 13445 5035
rect 13479 5001 13517 5035
rect 13551 5001 13589 5035
rect 13623 5001 13661 5035
rect 13695 5001 13733 5035
rect 13767 5001 13805 5035
rect 13839 5001 13877 5035
rect 13911 5001 13949 5035
rect 13983 5001 14021 5035
rect 14055 5001 14093 5035
rect 14127 5001 14165 5035
rect 14199 5001 14237 5035
rect 14271 5001 14309 5035
rect 14343 5001 14381 5035
rect 14415 5001 14453 5035
rect 14487 5001 14525 5035
rect 14559 5001 14597 5035
rect 14631 5001 14669 5035
rect 14703 5001 14741 5035
rect 14775 5030 14907 5035
rect 14775 5001 14835 5030
rect 303 5000 14835 5001
rect 231 4966 252 5000
rect 303 4995 320 5000
rect 286 4966 320 4995
rect 354 4966 388 5000
rect 422 4966 456 5000
rect 490 4966 524 5000
rect 558 4966 592 5000
rect 626 4966 660 5000
rect 694 4966 728 5000
rect 762 4966 796 5000
rect 830 4966 864 5000
rect 898 4966 932 5000
rect 966 4966 1000 5000
rect 1034 4966 1068 5000
rect 1102 4966 1136 5000
rect 1170 4966 1204 5000
rect 1238 4966 1272 5000
rect 1306 4966 1340 5000
rect 1374 4966 1408 5000
rect 1442 4966 1476 5000
rect 1510 4966 1544 5000
rect 1578 4966 1612 5000
rect 1646 4966 1680 5000
rect 1714 4966 1748 5000
rect 1782 4966 1816 5000
rect 1850 4966 1884 5000
rect 1918 4966 1952 5000
rect 1986 4966 2020 5000
rect 2054 4966 2088 5000
rect 2122 4966 2156 5000
rect 2190 4966 2224 5000
rect 2258 4966 2292 5000
rect 2326 4966 2360 5000
rect 2394 4966 2428 5000
rect 2462 4966 2496 5000
rect 2530 4966 2564 5000
rect 2598 4966 2632 5000
rect 2666 4966 2700 5000
rect 2734 4966 2768 5000
rect 2802 4966 2836 5000
rect 2870 4966 2904 5000
rect 2938 4966 2972 5000
rect 3006 4966 3040 5000
rect 3074 4966 3108 5000
rect 3142 4966 3176 5000
rect 3210 4966 3244 5000
rect 3278 4966 3312 5000
rect 3346 4966 3380 5000
rect 3414 4966 3448 5000
rect 3482 4966 3516 5000
rect 3550 4966 3584 5000
rect 3618 4966 3652 5000
rect 3686 4966 3720 5000
rect 3754 4966 3788 5000
rect 3822 4966 3856 5000
rect 3890 4966 3924 5000
rect 3958 4966 3992 5000
rect 4026 4966 4060 5000
rect 4094 4966 4128 5000
rect 4162 4966 4196 5000
rect 4230 4966 4264 5000
rect 4298 4966 4332 5000
rect 4366 4966 4400 5000
rect 4434 4966 4468 5000
rect 4502 4966 4536 5000
rect 4570 4966 4604 5000
rect 4638 4966 4672 5000
rect 4706 4966 4740 5000
rect 4774 4966 4808 5000
rect 4842 4966 4876 5000
rect 4910 4966 4944 5000
rect 4978 4966 5012 5000
rect 5046 4966 5080 5000
rect 5114 4966 5148 5000
rect 5182 4966 5216 5000
rect 5250 4966 5284 5000
rect 5318 4966 5352 5000
rect 5386 4966 5420 5000
rect 5454 4966 5488 5000
rect 5522 4966 5556 5000
rect 5590 4966 5624 5000
rect 5658 4966 5692 5000
rect 5726 4966 5760 5000
rect 5794 4966 5828 5000
rect 5862 4966 5896 5000
rect 5930 4966 5964 5000
rect 5998 4966 6032 5000
rect 6066 4966 6100 5000
rect 6134 4966 6168 5000
rect 6202 4966 6236 5000
rect 6270 4966 6304 5000
rect 6338 4966 6372 5000
rect 6406 4966 6440 5000
rect 6474 4966 6508 5000
rect 6542 4966 6576 5000
rect 6610 4966 6644 5000
rect 6678 4966 6712 5000
rect 6746 4966 6780 5000
rect 6814 4966 6848 5000
rect 6882 4966 6916 5000
rect 6950 4966 6984 5000
rect 7018 4966 7052 5000
rect 7086 4966 7120 5000
rect 7154 4966 7188 5000
rect 7222 4966 7256 5000
rect 7290 4966 7324 5000
rect 7358 4966 7392 5000
rect 7426 4966 7460 5000
rect 7494 4966 7528 5000
rect 7562 4966 7596 5000
rect 7630 4966 7664 5000
rect 7698 4966 7732 5000
rect 7766 4966 7800 5000
rect 7834 4966 7868 5000
rect 7902 4966 7936 5000
rect 7970 4966 8004 5000
rect 8038 4966 8072 5000
rect 8106 4966 8140 5000
rect 8174 4966 8208 5000
rect 8242 4966 8276 5000
rect 8310 4966 8344 5000
rect 8378 4966 8412 5000
rect 8446 4966 8480 5000
rect 8514 4966 8548 5000
rect 8582 4966 8616 5000
rect 8650 4966 8684 5000
rect 8718 4966 8752 5000
rect 8786 4966 8820 5000
rect 8854 4966 8888 5000
rect 8922 4966 8956 5000
rect 8990 4966 9024 5000
rect 9058 4966 9092 5000
rect 9126 4966 9160 5000
rect 9194 4966 9228 5000
rect 9262 4966 9296 5000
rect 9330 4966 9364 5000
rect 9398 4966 9432 5000
rect 9466 4966 9500 5000
rect 9534 4966 9568 5000
rect 9602 4966 9636 5000
rect 9670 4966 9704 5000
rect 9738 4966 9772 5000
rect 9806 4966 9840 5000
rect 9874 4966 9908 5000
rect 9942 4966 9976 5000
rect 10010 4966 10044 5000
rect 10078 4966 10112 5000
rect 10146 4966 10180 5000
rect 10214 4966 10248 5000
rect 10282 4966 10316 5000
rect 10350 4966 10384 5000
rect 10418 4966 10452 5000
rect 10486 4966 10520 5000
rect 10554 4966 10588 5000
rect 10622 4966 10656 5000
rect 10690 4966 10724 5000
rect 10758 4966 10792 5000
rect 10826 4966 10860 5000
rect 10894 4966 10928 5000
rect 10962 4966 10996 5000
rect 11030 4966 11064 5000
rect 11098 4966 11132 5000
rect 11166 4966 11200 5000
rect 11234 4966 11268 5000
rect 11302 4966 11336 5000
rect 11370 4966 11404 5000
rect 11438 4966 11472 5000
rect 11506 4966 11540 5000
rect 11574 4966 11608 5000
rect 11642 4966 11676 5000
rect 11710 4966 11744 5000
rect 11778 4966 11812 5000
rect 11846 4966 11880 5000
rect 11914 4966 11948 5000
rect 11982 4966 12016 5000
rect 12050 4966 12084 5000
rect 12118 4966 12152 5000
rect 12186 4966 12220 5000
rect 12254 4966 12288 5000
rect 12322 4966 12356 5000
rect 12390 4966 12424 5000
rect 12458 4966 12492 5000
rect 12526 4966 12560 5000
rect 12594 4966 12628 5000
rect 12662 4966 12696 5000
rect 12730 4966 12764 5000
rect 12798 4966 12832 5000
rect 12866 4966 12900 5000
rect 12934 4966 12968 5000
rect 13002 4966 13036 5000
rect 13070 4966 13104 5000
rect 13138 4966 13172 5000
rect 13206 4966 13240 5000
rect 13274 4966 13308 5000
rect 13342 4966 13376 5000
rect 13410 4966 13444 5000
rect 13478 4966 13512 5000
rect 13546 4966 13580 5000
rect 13614 4966 13648 5000
rect 13682 4966 13716 5000
rect 13750 4966 13784 5000
rect 13818 4966 13852 5000
rect 13886 4966 13920 5000
rect 13954 4966 13988 5000
rect 14022 4966 14056 5000
rect 14090 4966 14124 5000
rect 14158 4966 14192 5000
rect 14226 4966 14260 5000
rect 14294 4966 14328 5000
rect 14362 4966 14396 5000
rect 14430 4966 14464 5000
rect 14498 4966 14532 5000
rect 14566 4966 14600 5000
rect 14634 4966 14668 5000
rect 14702 4966 14736 5000
rect 14770 4966 14804 5000
rect 231 4959 14835 4966
rect 231 4956 361 4959
rect 231 4922 269 4956
rect 303 4925 361 4956
rect 395 4925 434 4959
rect 468 4925 507 4959
rect 541 4925 580 4959
rect 614 4925 653 4959
rect 687 4925 726 4959
rect 760 4925 799 4959
rect 833 4925 872 4959
rect 906 4925 945 4959
rect 979 4925 1018 4959
rect 1052 4925 1091 4959
rect 1125 4925 1164 4959
rect 1198 4925 1237 4959
rect 1271 4925 1310 4959
rect 1344 4925 1383 4959
rect 1417 4925 1456 4959
rect 1490 4925 1529 4959
rect 1563 4925 1602 4959
rect 1636 4925 1675 4959
rect 1709 4925 1748 4959
rect 1782 4925 1821 4959
rect 1855 4925 1894 4959
rect 1928 4925 1967 4959
rect 2001 4925 2040 4959
rect 2074 4925 2113 4959
rect 2147 4925 2186 4959
rect 2220 4925 2259 4959
rect 2293 4925 2332 4959
rect 2366 4925 2405 4959
rect 2439 4925 2478 4959
rect 2512 4925 2551 4959
rect 2585 4925 2624 4959
rect 2658 4925 2697 4959
rect 2731 4925 2770 4959
rect 2804 4925 2843 4959
rect 2877 4925 2916 4959
rect 2950 4925 2989 4959
rect 3023 4925 3062 4959
rect 3096 4925 3135 4959
rect 3169 4925 3208 4959
rect 3242 4925 3281 4959
rect 3315 4925 3354 4959
rect 3388 4925 3427 4959
rect 3461 4925 3500 4959
rect 3534 4925 3573 4959
rect 3607 4925 3646 4959
rect 3680 4925 3719 4959
rect 3753 4925 3792 4959
rect 3826 4925 3865 4959
rect 3899 4925 3938 4959
rect 3972 4925 4011 4959
rect 4045 4925 4084 4959
rect 4118 4925 4157 4959
rect 4191 4925 4229 4959
rect 4263 4925 4301 4959
rect 4335 4925 4373 4959
rect 4407 4925 4445 4959
rect 4479 4925 4517 4959
rect 4551 4925 4589 4959
rect 4623 4925 4661 4959
rect 4695 4925 4733 4959
rect 4767 4925 4805 4959
rect 4839 4925 4877 4959
rect 4911 4925 4949 4959
rect 4983 4925 5021 4959
rect 5055 4925 5093 4959
rect 5127 4925 5165 4959
rect 5199 4925 5237 4959
rect 5271 4925 5309 4959
rect 5343 4925 5381 4959
rect 5415 4925 5453 4959
rect 5487 4925 5525 4959
rect 5559 4925 5597 4959
rect 5631 4925 5669 4959
rect 5703 4925 5741 4959
rect 5775 4925 5813 4959
rect 5847 4925 5885 4959
rect 5919 4925 5957 4959
rect 5991 4925 6029 4959
rect 6063 4925 6101 4959
rect 6135 4925 6173 4959
rect 6207 4925 6245 4959
rect 6279 4925 6317 4959
rect 6351 4925 6389 4959
rect 6423 4925 6461 4959
rect 6495 4925 6533 4959
rect 6567 4925 6605 4959
rect 6639 4925 6677 4959
rect 6711 4925 6749 4959
rect 6783 4925 6821 4959
rect 6855 4925 6893 4959
rect 6927 4925 6965 4959
rect 6999 4925 7037 4959
rect 7071 4925 7109 4959
rect 7143 4925 7181 4959
rect 7215 4925 7253 4959
rect 7287 4925 7325 4959
rect 7359 4925 7397 4959
rect 7431 4925 7469 4959
rect 7503 4925 7541 4959
rect 7575 4925 7613 4959
rect 7647 4925 7685 4959
rect 7719 4925 7757 4959
rect 7791 4925 7829 4959
rect 7863 4925 7901 4959
rect 7935 4925 7973 4959
rect 8007 4925 8045 4959
rect 8079 4925 8117 4959
rect 8151 4925 8189 4959
rect 8223 4925 8261 4959
rect 8295 4925 8333 4959
rect 8367 4925 8405 4959
rect 8439 4925 8477 4959
rect 8511 4925 8549 4959
rect 8583 4925 8621 4959
rect 8655 4925 8693 4959
rect 8727 4925 8765 4959
rect 8799 4925 8837 4959
rect 8871 4925 8909 4959
rect 8943 4925 8981 4959
rect 9015 4925 9053 4959
rect 9087 4925 9125 4959
rect 9159 4925 9197 4959
rect 9231 4925 9269 4959
rect 9303 4925 9341 4959
rect 9375 4925 9413 4959
rect 9447 4925 9485 4959
rect 9519 4925 9557 4959
rect 9591 4925 9629 4959
rect 9663 4925 9701 4959
rect 9735 4925 9773 4959
rect 9807 4925 9845 4959
rect 9879 4925 9917 4959
rect 9951 4925 9989 4959
rect 10023 4925 10061 4959
rect 10095 4925 10133 4959
rect 10167 4925 10205 4959
rect 10239 4925 10277 4959
rect 10311 4925 10349 4959
rect 10383 4925 10421 4959
rect 10455 4925 10493 4959
rect 10527 4925 10565 4959
rect 10599 4925 10637 4959
rect 10671 4925 10709 4959
rect 10743 4925 10781 4959
rect 10815 4925 10853 4959
rect 10887 4925 10925 4959
rect 10959 4925 10997 4959
rect 11031 4925 11069 4959
rect 11103 4925 11141 4959
rect 11175 4925 11213 4959
rect 11247 4925 11285 4959
rect 11319 4925 11357 4959
rect 11391 4925 11429 4959
rect 11463 4925 11501 4959
rect 11535 4925 11573 4959
rect 11607 4925 11645 4959
rect 11679 4925 11717 4959
rect 11751 4925 11789 4959
rect 11823 4925 11861 4959
rect 11895 4925 11933 4959
rect 11967 4925 12005 4959
rect 12039 4925 12077 4959
rect 12111 4925 12149 4959
rect 12183 4925 12221 4959
rect 12255 4925 12293 4959
rect 12327 4925 12365 4959
rect 12399 4925 12437 4959
rect 12471 4925 12509 4959
rect 12543 4925 12581 4959
rect 12615 4925 12653 4959
rect 12687 4925 12725 4959
rect 12759 4925 12797 4959
rect 12831 4925 12869 4959
rect 12903 4925 12941 4959
rect 12975 4925 13013 4959
rect 13047 4925 13085 4959
rect 13119 4925 13157 4959
rect 13191 4925 13229 4959
rect 13263 4925 13301 4959
rect 13335 4925 13373 4959
rect 13407 4925 13445 4959
rect 13479 4925 13517 4959
rect 13551 4925 13589 4959
rect 13623 4925 13661 4959
rect 13695 4925 13733 4959
rect 13767 4925 13805 4959
rect 13839 4925 13877 4959
rect 13911 4925 13949 4959
rect 13983 4925 14021 4959
rect 14055 4925 14093 4959
rect 14127 4925 14165 4959
rect 14199 4925 14237 4959
rect 14271 4925 14309 4959
rect 14343 4925 14381 4959
rect 14415 4925 14453 4959
rect 14487 4925 14525 4959
rect 14559 4925 14597 4959
rect 14631 4925 14669 4959
rect 14703 4925 14741 4959
rect 14775 4925 14835 4959
rect 303 4922 14835 4925
rect 231 4918 14835 4922
rect 231 4884 252 4918
rect 286 4884 320 4918
rect 354 4884 388 4918
rect 422 4884 456 4918
rect 490 4884 524 4918
rect 558 4884 592 4918
rect 626 4884 660 4918
rect 694 4884 728 4918
rect 762 4884 796 4918
rect 830 4884 864 4918
rect 898 4884 932 4918
rect 966 4884 1000 4918
rect 1034 4884 1068 4918
rect 1102 4884 1136 4918
rect 1170 4884 1204 4918
rect 1238 4884 1272 4918
rect 1306 4884 1340 4918
rect 1374 4884 1408 4918
rect 1442 4884 1476 4918
rect 1510 4884 1544 4918
rect 1578 4884 1612 4918
rect 1646 4884 1680 4918
rect 1714 4884 1748 4918
rect 1782 4884 1816 4918
rect 1850 4884 1884 4918
rect 1918 4884 1952 4918
rect 1986 4884 2020 4918
rect 2054 4884 2088 4918
rect 2122 4884 2156 4918
rect 2190 4884 2224 4918
rect 2258 4884 2292 4918
rect 2326 4884 2360 4918
rect 2394 4884 2428 4918
rect 2462 4884 2496 4918
rect 2530 4884 2564 4918
rect 2598 4884 2632 4918
rect 2666 4884 2700 4918
rect 2734 4884 2768 4918
rect 2802 4884 2836 4918
rect 2870 4884 2904 4918
rect 2938 4884 2972 4918
rect 3006 4884 3040 4918
rect 3074 4884 3108 4918
rect 3142 4884 3176 4918
rect 3210 4884 3244 4918
rect 3278 4884 3312 4918
rect 3346 4884 3380 4918
rect 3414 4884 3448 4918
rect 3482 4884 3516 4918
rect 3550 4884 3584 4918
rect 3618 4884 3652 4918
rect 3686 4884 3720 4918
rect 3754 4884 3788 4918
rect 3822 4884 3856 4918
rect 3890 4884 3924 4918
rect 3958 4884 3992 4918
rect 4026 4884 4060 4918
rect 4094 4884 4128 4918
rect 4162 4884 4196 4918
rect 4230 4884 4264 4918
rect 4298 4884 4332 4918
rect 4366 4884 4400 4918
rect 4434 4884 4468 4918
rect 4502 4884 4536 4918
rect 4570 4884 4604 4918
rect 4638 4884 4672 4918
rect 4706 4884 4740 4918
rect 4774 4884 4808 4918
rect 4842 4884 4876 4918
rect 4910 4884 4944 4918
rect 4978 4884 5012 4918
rect 5046 4884 5080 4918
rect 5114 4884 5148 4918
rect 5182 4884 5216 4918
rect 5250 4884 5284 4918
rect 5318 4884 5352 4918
rect 5386 4884 5420 4918
rect 5454 4884 5488 4918
rect 5522 4884 5556 4918
rect 5590 4884 5624 4918
rect 5658 4884 5692 4918
rect 5726 4884 5760 4918
rect 5794 4884 5828 4918
rect 5862 4884 5896 4918
rect 5930 4884 5964 4918
rect 5998 4884 6032 4918
rect 6066 4884 6100 4918
rect 6134 4884 6168 4918
rect 6202 4884 6236 4918
rect 6270 4884 6304 4918
rect 6338 4884 6372 4918
rect 6406 4884 6440 4918
rect 6474 4884 6508 4918
rect 6542 4884 6576 4918
rect 6610 4884 6644 4918
rect 6678 4884 6712 4918
rect 6746 4884 6780 4918
rect 6814 4884 6848 4918
rect 6882 4884 6916 4918
rect 6950 4884 6984 4918
rect 7018 4884 7052 4918
rect 7086 4884 7120 4918
rect 7154 4884 7188 4918
rect 7222 4884 7256 4918
rect 7290 4884 7324 4918
rect 7358 4884 7392 4918
rect 7426 4884 7460 4918
rect 7494 4884 7528 4918
rect 7562 4884 7596 4918
rect 7630 4884 7664 4918
rect 7698 4884 7732 4918
rect 7766 4884 7800 4918
rect 7834 4884 7868 4918
rect 7902 4884 7936 4918
rect 7970 4884 8004 4918
rect 8038 4884 8072 4918
rect 8106 4884 8140 4918
rect 8174 4884 8208 4918
rect 8242 4884 8276 4918
rect 8310 4884 8344 4918
rect 8378 4884 8412 4918
rect 8446 4884 8480 4918
rect 8514 4884 8548 4918
rect 8582 4884 8616 4918
rect 8650 4884 8684 4918
rect 8718 4884 8752 4918
rect 8786 4884 8820 4918
rect 8854 4884 8888 4918
rect 8922 4884 8956 4918
rect 8990 4884 9024 4918
rect 9058 4884 9092 4918
rect 9126 4884 9160 4918
rect 9194 4884 9228 4918
rect 9262 4884 9296 4918
rect 9330 4884 9364 4918
rect 9398 4884 9432 4918
rect 9466 4884 9500 4918
rect 9534 4884 9568 4918
rect 9602 4884 9636 4918
rect 9670 4884 9704 4918
rect 9738 4884 9772 4918
rect 9806 4884 9840 4918
rect 9874 4884 9908 4918
rect 9942 4884 9976 4918
rect 10010 4884 10044 4918
rect 10078 4884 10112 4918
rect 10146 4884 10180 4918
rect 10214 4884 10248 4918
rect 10282 4884 10316 4918
rect 10350 4884 10384 4918
rect 10418 4884 10452 4918
rect 10486 4884 10520 4918
rect 10554 4884 10588 4918
rect 10622 4884 10656 4918
rect 10690 4884 10724 4918
rect 10758 4884 10792 4918
rect 10826 4884 10860 4918
rect 10894 4884 10928 4918
rect 10962 4884 10996 4918
rect 11030 4884 11064 4918
rect 11098 4884 11132 4918
rect 11166 4884 11200 4918
rect 11234 4884 11268 4918
rect 11302 4884 11336 4918
rect 11370 4884 11404 4918
rect 11438 4884 11472 4918
rect 11506 4884 11540 4918
rect 11574 4884 11608 4918
rect 11642 4884 11676 4918
rect 11710 4884 11744 4918
rect 11778 4884 11812 4918
rect 11846 4884 11880 4918
rect 11914 4884 11948 4918
rect 11982 4884 12016 4918
rect 12050 4884 12084 4918
rect 12118 4884 12152 4918
rect 12186 4884 12220 4918
rect 12254 4884 12288 4918
rect 12322 4884 12356 4918
rect 12390 4884 12424 4918
rect 12458 4884 12492 4918
rect 12526 4884 12560 4918
rect 12594 4884 12628 4918
rect 12662 4884 12696 4918
rect 12730 4884 12764 4918
rect 12798 4884 12832 4918
rect 12866 4884 12900 4918
rect 12934 4884 12968 4918
rect 13002 4884 13036 4918
rect 13070 4884 13104 4918
rect 13138 4884 13172 4918
rect 13206 4884 13240 4918
rect 13274 4884 13308 4918
rect 13342 4884 13376 4918
rect 13410 4884 13444 4918
rect 13478 4884 13512 4918
rect 13546 4884 13580 4918
rect 13614 4884 13648 4918
rect 13682 4884 13716 4918
rect 13750 4884 13784 4918
rect 13818 4884 13852 4918
rect 13886 4884 13920 4918
rect 13954 4884 13988 4918
rect 14022 4884 14056 4918
rect 14090 4884 14124 4918
rect 14158 4884 14192 4918
rect 14226 4884 14260 4918
rect 14294 4884 14328 4918
rect 14362 4884 14396 4918
rect 14430 4884 14464 4918
rect 14498 4884 14532 4918
rect 14566 4884 14600 4918
rect 14634 4884 14668 4918
rect 14702 4884 14736 4918
rect 14770 4884 14804 4918
rect 231 4883 14835 4884
rect 231 4849 269 4883
rect 303 4849 329 4883
rect 295 4810 329 4849
rect 303 4776 329 4810
rect 295 4737 329 4776
rect 303 4703 329 4737
rect 295 4664 329 4703
rect 303 4630 329 4664
rect 14806 4849 14835 4883
rect 14806 4781 14835 4815
rect 14806 4713 14835 4747
rect 295 4591 329 4630
rect 303 4557 329 4591
rect 295 4518 329 4557
rect 303 4484 329 4518
rect 295 4445 329 4484
rect 303 4411 329 4445
rect 295 4372 329 4411
rect 303 4338 329 4372
rect 295 4299 329 4338
rect 303 4265 329 4299
rect 295 4226 329 4265
rect 303 4192 329 4226
rect 295 4153 329 4192
rect 303 4119 329 4153
rect 295 4080 329 4119
rect 303 4046 329 4080
rect 295 4007 329 4046
rect 303 3973 329 4007
rect 295 3934 329 3973
rect 303 3900 329 3934
rect 295 3861 329 3900
rect 303 3827 329 3861
rect 295 3788 329 3827
rect 303 3754 329 3788
rect 295 3715 329 3754
rect 303 3681 329 3715
rect 295 3642 329 3681
rect 303 3608 329 3642
rect 295 3569 329 3608
rect 303 3535 329 3569
rect 295 3496 329 3535
rect 303 3462 329 3496
rect 295 3423 329 3462
rect 303 3389 329 3423
rect 295 3350 329 3389
rect 303 3316 329 3350
rect 295 3277 329 3316
rect 303 3243 329 3277
rect 295 3204 329 3243
rect 303 3170 329 3204
rect 295 3131 329 3170
rect 303 3097 329 3131
rect 295 3058 329 3097
rect 303 3024 329 3058
rect 295 2985 329 3024
rect 303 2951 329 2985
rect 295 2912 329 2951
rect 303 2878 329 2912
rect 295 2839 329 2878
rect 303 2805 329 2839
rect 295 2766 329 2805
rect 303 2732 329 2766
rect 295 2693 329 2732
rect 303 2659 329 2693
rect 295 2620 329 2659
rect 303 2586 329 2620
rect 295 2547 329 2586
rect 303 2513 329 2547
rect 295 2474 329 2513
rect 303 2440 329 2474
rect 295 2401 329 2440
rect 303 2367 329 2401
rect 295 2328 329 2367
rect 303 2294 329 2328
rect 295 2255 329 2294
rect 303 2221 329 2255
rect 295 2182 329 2221
rect 303 2148 329 2182
rect 295 2109 329 2148
rect 303 2075 329 2109
rect 295 2036 329 2075
rect 303 2002 329 2036
rect 295 1963 329 2002
rect 303 1929 329 1963
rect 295 1890 329 1929
rect 303 1856 329 1890
rect 295 1817 329 1856
rect 303 1783 329 1817
rect 295 1744 329 1783
rect 303 1710 329 1744
rect 295 1671 329 1710
rect 303 1637 329 1671
rect 295 1598 329 1637
rect 303 1564 329 1598
rect 295 1525 329 1564
rect 303 1491 329 1525
rect 295 1452 329 1491
rect 303 1418 329 1452
rect 295 1379 329 1418
rect 303 1345 329 1379
rect 295 1306 329 1345
rect 303 1272 329 1306
rect 295 1233 329 1272
rect 303 1199 329 1233
rect 295 1159 329 1199
rect 303 1125 329 1159
rect 295 1085 329 1125
rect 303 1051 329 1085
rect 295 1011 329 1051
rect 303 977 329 1011
rect 295 937 329 977
rect 303 903 329 937
rect 295 863 329 903
rect 303 829 329 863
rect 295 789 329 829
rect 303 755 329 789
rect 295 715 329 755
rect 303 681 329 715
rect 295 641 329 681
rect 482 4638 14653 4653
rect 482 4619 584 4638
rect 482 4585 497 4619
rect 531 4585 584 4619
rect 10410 4606 10445 4638
rect 10479 4606 10514 4638
rect 10548 4606 10583 4638
rect 10617 4606 10652 4638
rect 10686 4606 10721 4638
rect 10755 4606 10790 4638
rect 10824 4606 10859 4638
rect 10893 4606 10928 4638
rect 10962 4606 10997 4638
rect 11031 4606 11066 4638
rect 11100 4606 11135 4638
rect 11169 4606 11204 4638
rect 11238 4606 11273 4638
rect 11307 4606 11342 4638
rect 11376 4606 11411 4638
rect 11445 4606 11480 4638
rect 11514 4606 11549 4638
rect 11583 4606 11618 4638
rect 11652 4606 11687 4638
rect 11721 4606 11756 4638
rect 11790 4606 11825 4638
rect 11859 4606 11894 4638
rect 11928 4606 11963 4638
rect 11997 4606 12032 4638
rect 12066 4606 12101 4638
rect 12135 4606 12170 4638
rect 12204 4606 12239 4638
rect 12273 4606 12308 4638
rect 12342 4606 12377 4638
rect 12411 4606 12446 4638
rect 12480 4606 12515 4638
rect 12549 4606 12584 4638
rect 12618 4606 12653 4638
rect 12687 4606 12722 4638
rect 12756 4606 12791 4638
rect 12825 4606 12860 4638
rect 12894 4606 12929 4638
rect 12963 4606 12998 4638
rect 13032 4606 13067 4638
rect 13101 4606 13136 4638
rect 13170 4606 13205 4638
rect 13239 4606 13274 4638
rect 13308 4606 13343 4638
rect 13377 4606 13412 4638
rect 13446 4606 13481 4638
rect 13515 4606 13550 4638
rect 13584 4606 13619 4638
rect 13653 4606 13688 4638
rect 13722 4606 13757 4638
rect 13791 4606 13826 4638
rect 13860 4606 13895 4638
rect 13929 4606 13964 4638
rect 13998 4606 14033 4638
rect 14067 4606 14102 4638
rect 14136 4606 14171 4638
rect 14205 4606 14240 4638
rect 14274 4606 14309 4638
rect 14343 4606 14378 4638
rect 14412 4606 14447 4638
rect 482 4570 584 4585
rect 14207 4604 14240 4606
rect 14280 4604 14309 4606
rect 14353 4604 14378 4606
rect 14426 4604 14447 4606
rect 14481 4604 14516 4638
rect 14550 4604 14585 4638
rect 14619 4604 14653 4638
rect 14207 4572 14246 4604
rect 14280 4572 14319 4604
rect 14353 4572 14392 4604
rect 14426 4572 14653 4604
rect 14207 4570 14653 4572
rect 482 4549 565 4570
rect 482 4515 497 4549
rect 531 4536 565 4549
rect 531 4515 633 4536
rect 482 4498 633 4515
rect 14225 4536 14260 4570
rect 14294 4536 14329 4570
rect 14363 4536 14398 4570
rect 14432 4536 14467 4570
rect 14501 4536 14536 4570
rect 14570 4551 14653 4570
rect 14207 4534 14536 4536
rect 14207 4502 14246 4534
rect 14280 4502 14319 4534
rect 14353 4502 14392 4534
rect 14426 4502 14536 4534
rect 14226 4500 14246 4502
rect 14295 4500 14319 4502
rect 14364 4500 14392 4502
rect 482 4479 565 4498
rect 482 4445 497 4479
rect 531 4464 565 4479
rect 599 4468 633 4498
rect 12363 4468 12398 4500
rect 12432 4468 12467 4500
rect 12501 4468 12536 4500
rect 12570 4468 12605 4500
rect 12639 4468 12674 4500
rect 12708 4468 12743 4500
rect 12777 4468 12812 4500
rect 12846 4468 12881 4500
rect 12915 4468 12950 4500
rect 12984 4468 13019 4500
rect 13053 4468 13088 4500
rect 13122 4468 13157 4500
rect 13191 4468 13226 4500
rect 13260 4468 13295 4500
rect 13329 4468 13364 4500
rect 13398 4468 13433 4500
rect 13467 4468 13502 4500
rect 13536 4468 13571 4500
rect 13605 4468 13640 4500
rect 13674 4468 13709 4500
rect 13743 4468 13778 4500
rect 13812 4468 13847 4500
rect 13881 4468 13916 4500
rect 13950 4468 13985 4500
rect 14019 4468 14054 4500
rect 14088 4468 14123 4500
rect 14157 4468 14192 4500
rect 14226 4468 14261 4500
rect 14295 4468 14330 4500
rect 14364 4468 14399 4500
rect 14433 4468 14468 4502
rect 599 4464 14468 4468
rect 531 4456 14468 4464
rect 531 4445 674 4456
rect 708 4453 14428 4456
rect 708 4445 780 4453
rect 482 4429 674 4445
rect 482 4426 633 4429
rect 482 4409 529 4426
rect 482 4375 497 4409
rect 563 4392 565 4426
rect 599 4392 601 4426
rect 667 4395 674 4429
rect 635 4392 674 4395
rect 531 4375 674 4392
rect 482 4356 674 4375
rect 482 4354 633 4356
rect 482 4351 565 4354
rect 482 4339 529 4351
rect 482 4305 497 4339
rect 563 4320 565 4351
rect 599 4351 633 4354
rect 599 4320 601 4351
rect 667 4322 674 4356
rect 563 4317 601 4320
rect 635 4317 674 4322
rect 531 4305 674 4317
rect 482 4283 674 4305
rect 482 4282 633 4283
rect 482 4276 565 4282
rect 482 4269 529 4276
rect 482 4235 497 4269
rect 563 4248 565 4276
rect 599 4276 633 4282
rect 599 4248 601 4276
rect 667 4249 674 4283
rect 563 4242 601 4248
rect 635 4242 674 4249
rect 531 4235 674 4242
rect 482 4211 674 4235
rect 482 4210 633 4211
rect 482 4201 565 4210
rect 482 4199 529 4201
rect 482 4165 497 4199
rect 563 4176 565 4201
rect 599 4201 633 4210
rect 599 4176 601 4201
rect 667 4177 674 4211
rect 563 4167 601 4176
rect 635 4167 674 4177
rect 531 4165 674 4167
rect 482 4139 674 4165
rect 482 4138 633 4139
rect 482 4129 565 4138
rect 482 4095 497 4129
rect 531 4126 565 4129
rect 563 4104 565 4126
rect 599 4126 633 4138
rect 599 4104 601 4126
rect 667 4105 674 4139
rect 482 4092 529 4095
rect 563 4092 601 4104
rect 635 4092 674 4105
rect 482 4067 674 4092
rect 14356 4432 14428 4453
rect 14390 4398 14428 4432
rect 14462 4426 14468 4456
rect 14356 4359 14428 4398
rect 14390 4325 14428 4359
rect 482 4066 633 4067
rect 482 4059 565 4066
rect 482 4025 497 4059
rect 531 4052 565 4059
rect 563 4032 565 4052
rect 599 4052 633 4066
rect 599 4032 601 4052
rect 667 4033 674 4067
rect 482 4018 529 4025
rect 563 4018 601 4032
rect 635 4018 674 4033
rect 482 3995 674 4018
rect 482 3994 633 3995
rect 482 3989 565 3994
rect 482 3955 497 3989
rect 531 3978 565 3989
rect 563 3960 565 3978
rect 599 3978 633 3994
rect 599 3960 601 3978
rect 667 3961 674 3995
rect 482 3944 529 3955
rect 563 3944 601 3960
rect 635 3944 674 3961
rect 482 3923 674 3944
rect 482 3922 633 3923
rect 482 3920 565 3922
rect 482 3886 497 3920
rect 531 3904 565 3920
rect 563 3888 565 3904
rect 599 3904 633 3922
rect 599 3888 601 3904
rect 667 3889 674 3923
rect 482 3870 529 3886
rect 563 3870 601 3888
rect 635 3870 674 3889
rect 482 3851 674 3870
rect 482 3817 497 3851
rect 531 3817 565 3851
rect 599 3817 633 3851
rect 667 3817 674 3851
rect 482 3794 674 3817
rect 482 3760 529 3794
rect 563 3760 601 3794
rect 635 3760 674 3794
rect 482 3749 674 3760
rect 482 3715 497 3749
rect 531 3720 565 3749
rect 563 3715 565 3720
rect 599 3720 633 3749
rect 599 3715 601 3720
rect 667 3715 674 3749
rect 482 3686 529 3715
rect 563 3686 601 3715
rect 635 3686 674 3715
rect 482 3680 674 3686
rect 482 3646 497 3680
rect 531 3646 565 3680
rect 599 3646 633 3680
rect 667 3646 674 3680
rect 482 3612 529 3646
rect 563 3612 601 3646
rect 635 3612 674 3646
rect 482 3611 674 3612
rect 482 3577 497 3611
rect 531 3577 565 3611
rect 599 3577 633 3611
rect 667 3577 674 3611
rect 482 3572 674 3577
rect 482 3542 529 3572
rect 563 3542 601 3572
rect 635 3542 674 3572
rect 482 3508 497 3542
rect 563 3538 565 3542
rect 531 3508 565 3538
rect 599 3538 601 3542
rect 599 3508 633 3538
rect 667 3508 674 3542
rect 482 3498 674 3508
rect 482 3473 529 3498
rect 563 3473 601 3498
rect 635 3473 674 3498
rect 482 3439 497 3473
rect 563 3464 565 3473
rect 531 3439 565 3464
rect 599 3464 601 3473
rect 599 3439 633 3464
rect 667 3439 674 3473
rect 482 3424 674 3439
rect 482 3404 529 3424
rect 563 3404 601 3424
rect 635 3404 674 3424
rect 482 3370 497 3404
rect 563 3390 565 3404
rect 531 3370 565 3390
rect 599 3390 601 3404
rect 599 3370 633 3390
rect 667 3370 674 3404
rect 482 3350 674 3370
rect 482 3335 529 3350
rect 563 3335 601 3350
rect 635 3335 674 3350
rect 482 3301 497 3335
rect 563 3316 565 3335
rect 531 3301 565 3316
rect 599 3316 601 3335
rect 599 3301 633 3316
rect 667 3301 674 3335
rect 482 3276 674 3301
rect 482 3266 529 3276
rect 563 3266 601 3276
rect 635 3266 674 3276
rect 482 3232 497 3266
rect 563 3242 565 3266
rect 531 3232 565 3242
rect 599 3242 601 3266
rect 599 3232 633 3242
rect 667 3232 674 3266
rect 482 3202 674 3232
rect 482 3197 529 3202
rect 563 3197 601 3202
rect 635 3197 674 3202
rect 482 3163 497 3197
rect 563 3168 565 3197
rect 531 3163 565 3168
rect 599 3168 601 3197
rect 599 3163 633 3168
rect 667 3163 674 3197
rect 482 3128 674 3163
rect 482 3094 497 3128
rect 563 3094 565 3128
rect 599 3094 601 3128
rect 667 3094 674 3128
rect 482 3059 674 3094
rect 482 3025 497 3059
rect 531 3054 565 3059
rect 563 3025 565 3054
rect 599 3054 633 3059
rect 599 3025 601 3054
rect 667 3025 674 3059
rect 482 3020 529 3025
rect 563 3020 601 3025
rect 635 3020 674 3025
rect 482 2990 674 3020
rect 482 2956 497 2990
rect 531 2980 565 2990
rect 563 2956 565 2980
rect 599 2980 633 2990
rect 599 2956 601 2980
rect 667 2956 674 2990
rect 482 2946 529 2956
rect 563 2946 601 2956
rect 635 2946 674 2956
rect 482 2921 674 2946
rect 482 2887 497 2921
rect 531 2906 565 2921
rect 563 2887 565 2906
rect 599 2906 633 2921
rect 599 2887 601 2906
rect 667 2887 674 2921
rect 482 2872 529 2887
rect 563 2872 601 2887
rect 635 2872 674 2887
rect 482 2852 674 2872
rect 482 2818 497 2852
rect 531 2832 565 2852
rect 563 2818 565 2832
rect 599 2832 633 2852
rect 599 2818 601 2832
rect 667 2818 674 2852
rect 482 2798 529 2818
rect 563 2798 601 2818
rect 635 2798 674 2818
rect 482 2783 674 2798
rect 482 2749 497 2783
rect 531 2758 565 2783
rect 563 2749 565 2758
rect 599 2758 633 2783
rect 599 2749 601 2758
rect 667 2749 674 2783
rect 482 2724 529 2749
rect 563 2724 601 2749
rect 635 2724 674 2749
rect 482 2714 674 2724
rect 482 2680 497 2714
rect 531 2684 565 2714
rect 563 2680 565 2684
rect 599 2684 633 2714
rect 599 2680 601 2684
rect 667 2680 674 2714
rect 482 2650 529 2680
rect 563 2650 601 2680
rect 635 2650 674 2680
rect 482 2645 674 2650
rect 482 2611 497 2645
rect 531 2611 565 2645
rect 599 2611 633 2645
rect 667 2611 674 2645
rect 482 2610 674 2611
rect 482 2576 529 2610
rect 563 2576 601 2610
rect 635 2576 674 2610
rect 482 2542 497 2576
rect 531 2542 565 2576
rect 599 2542 633 2576
rect 667 2542 674 2576
rect 482 2536 674 2542
rect 482 2507 529 2536
rect 563 2507 601 2536
rect 635 2507 674 2536
rect 482 2473 497 2507
rect 563 2502 565 2507
rect 531 2473 565 2502
rect 599 2502 601 2507
rect 599 2473 633 2502
rect 667 2473 674 2507
rect 482 2462 674 2473
rect 482 2438 529 2462
rect 563 2438 601 2462
rect 635 2438 674 2462
rect 482 2404 497 2438
rect 563 2428 565 2438
rect 531 2404 565 2428
rect 599 2428 601 2438
rect 599 2404 633 2428
rect 667 2404 674 2438
rect 482 2389 674 2404
rect 482 2369 529 2389
rect 563 2369 601 2389
rect 635 2369 674 2389
rect 482 2335 497 2369
rect 563 2355 565 2369
rect 531 2335 565 2355
rect 599 2355 601 2369
rect 599 2335 633 2355
rect 667 2335 674 2369
rect 482 2316 674 2335
rect 482 2300 529 2316
rect 563 2300 601 2316
rect 635 2300 674 2316
rect 482 2266 497 2300
rect 563 2282 565 2300
rect 531 2266 565 2282
rect 599 2282 601 2300
rect 599 2266 633 2282
rect 667 2266 674 2300
rect 482 2243 674 2266
rect 482 2231 529 2243
rect 563 2231 601 2243
rect 635 2231 674 2243
rect 482 2197 497 2231
rect 563 2209 565 2231
rect 531 2197 565 2209
rect 599 2209 601 2231
rect 599 2197 633 2209
rect 667 2197 674 2231
rect 482 2170 674 2197
rect 482 2163 529 2170
rect 482 2129 497 2163
rect 563 2162 601 2170
rect 635 2162 674 2170
rect 563 2136 565 2162
rect 531 2129 565 2136
rect 482 2128 565 2129
rect 599 2136 601 2162
rect 599 2128 633 2136
rect 667 2128 674 2162
rect 482 2097 674 2128
rect 482 2095 529 2097
rect 482 2061 497 2095
rect 563 2093 601 2097
rect 635 2093 674 2097
rect 563 2063 565 2093
rect 531 2061 565 2063
rect 482 2059 565 2061
rect 599 2063 601 2093
rect 599 2059 633 2063
rect 667 2059 674 2093
rect 482 2027 674 2059
rect 482 1993 497 2027
rect 531 2024 674 2027
rect 482 1990 529 1993
rect 563 1990 565 2024
rect 599 1990 601 2024
rect 667 1990 674 2024
rect 482 1959 674 1990
rect 482 1925 497 1959
rect 531 1955 674 1959
rect 531 1951 565 1955
rect 482 1917 529 1925
rect 563 1921 565 1951
rect 599 1951 633 1955
rect 599 1921 601 1951
rect 667 1921 674 1955
rect 563 1917 601 1921
rect 635 1917 674 1921
rect 482 1891 674 1917
rect 482 1857 497 1891
rect 531 1886 674 1891
rect 531 1878 565 1886
rect 482 1844 529 1857
rect 563 1852 565 1878
rect 599 1878 633 1886
rect 599 1852 601 1878
rect 667 1852 674 1886
rect 563 1844 601 1852
rect 635 1844 674 1852
rect 482 1823 674 1844
rect 482 1789 497 1823
rect 531 1817 674 1823
rect 531 1805 565 1817
rect 482 1771 529 1789
rect 563 1783 565 1805
rect 599 1805 633 1817
rect 599 1783 601 1805
rect 667 1783 674 1817
rect 563 1771 601 1783
rect 635 1771 674 1783
rect 482 1755 674 1771
rect 482 1721 497 1755
rect 531 1748 674 1755
rect 531 1732 565 1748
rect 482 1698 529 1721
rect 563 1714 565 1732
rect 599 1732 633 1748
rect 599 1714 601 1732
rect 667 1714 674 1748
rect 563 1698 601 1714
rect 635 1698 674 1714
rect 482 1687 674 1698
rect 482 1653 497 1687
rect 531 1679 674 1687
rect 531 1659 565 1679
rect 482 1625 529 1653
rect 563 1645 565 1659
rect 599 1659 633 1679
rect 599 1645 601 1659
rect 667 1645 674 1679
rect 563 1625 601 1645
rect 635 1625 674 1645
rect 482 1619 674 1625
rect 482 1585 497 1619
rect 531 1610 674 1619
rect 531 1586 565 1610
rect 482 1552 529 1585
rect 563 1576 565 1586
rect 599 1586 633 1610
rect 599 1576 601 1586
rect 667 1576 674 1610
rect 563 1552 601 1576
rect 635 1552 674 1576
rect 482 1551 674 1552
rect 482 1517 497 1551
rect 531 1541 674 1551
rect 531 1517 565 1541
rect 482 1513 565 1517
rect 482 1483 529 1513
rect 563 1507 565 1513
rect 599 1513 633 1541
rect 599 1507 601 1513
rect 667 1507 674 1541
rect 482 1449 497 1483
rect 563 1479 601 1507
rect 635 1479 674 1507
rect 531 1472 674 1479
rect 531 1449 565 1472
rect 482 1440 565 1449
rect 482 1415 529 1440
rect 563 1438 565 1440
rect 599 1440 633 1472
rect 599 1438 601 1440
rect 667 1438 674 1472
rect 482 1381 497 1415
rect 563 1406 601 1438
rect 635 1406 674 1438
rect 531 1403 674 1406
rect 531 1381 565 1403
rect 482 1369 565 1381
rect 599 1369 633 1403
rect 667 1369 674 1403
rect 482 1367 674 1369
rect 482 1347 529 1367
rect 482 1313 497 1347
rect 563 1334 601 1367
rect 635 1334 674 1367
rect 563 1333 565 1334
rect 531 1313 565 1333
rect 482 1300 565 1313
rect 599 1333 601 1334
rect 599 1300 633 1333
rect 667 1300 674 1334
rect 482 1294 674 1300
rect 482 1279 529 1294
rect 482 1245 497 1279
rect 563 1265 601 1294
rect 635 1265 674 1294
rect 563 1260 565 1265
rect 531 1245 565 1260
rect 482 1231 565 1245
rect 599 1260 601 1265
rect 599 1231 633 1260
rect 667 1231 674 1265
rect 482 1221 674 1231
rect 482 1211 529 1221
rect 482 1177 497 1211
rect 563 1196 601 1221
rect 635 1196 674 1221
rect 563 1187 565 1196
rect 531 1177 565 1187
rect 482 1162 565 1177
rect 599 1187 601 1196
rect 599 1162 633 1187
rect 667 1162 674 1196
rect 482 1148 674 1162
rect 482 1143 529 1148
rect 482 1109 497 1143
rect 563 1127 601 1148
rect 635 1127 674 1148
rect 563 1114 565 1127
rect 531 1109 565 1114
rect 482 1093 565 1109
rect 599 1114 601 1127
rect 599 1093 633 1114
rect 667 1093 674 1127
rect 482 1075 674 1093
rect 482 1041 497 1075
rect 563 1058 601 1075
rect 635 1058 674 1075
rect 563 1041 565 1058
rect 482 1024 565 1041
rect 599 1041 601 1058
rect 599 1024 633 1041
rect 667 1024 674 1058
rect 482 1007 674 1024
rect 482 973 497 1007
rect 531 1002 674 1007
rect 563 989 601 1002
rect 635 989 674 1002
rect 482 968 529 973
rect 563 968 565 989
rect 482 955 565 968
rect 599 968 601 989
rect 599 955 633 968
rect 667 955 674 989
rect 482 939 674 955
rect 482 769 497 939
rect 531 929 674 939
rect 563 920 601 929
rect 635 920 674 929
rect 667 894 674 920
rect 881 4308 1001 4324
rect 881 4274 924 4308
rect 958 4274 1001 4308
rect 881 4234 1001 4274
rect 881 4200 924 4234
rect 958 4200 1001 4234
rect 881 3104 1001 4200
rect 1311 4308 1431 4324
rect 1311 4274 1354 4308
rect 1388 4274 1431 4308
rect 1311 4234 1431 4274
rect 1311 4200 1354 4234
rect 1388 4200 1431 4234
rect 881 3070 924 3104
rect 958 3070 1001 3104
rect 881 3026 1001 3070
rect 881 2992 924 3026
rect 958 2992 1001 3026
rect 881 2948 1001 2992
rect 881 2914 924 2948
rect 958 2914 1001 2948
rect 881 2870 1001 2914
rect 881 2836 924 2870
rect 958 2836 1001 2870
rect 881 2792 1001 2836
rect 881 2758 924 2792
rect 958 2758 1001 2792
rect 881 2713 1001 2758
rect 881 2679 924 2713
rect 958 2679 1001 2713
rect 881 2634 1001 2679
rect 881 2600 924 2634
rect 958 2600 1001 2634
rect 881 1504 1001 2600
rect 1066 4064 1067 4098
rect 1101 4082 1139 4098
rect 1101 4064 1103 4082
rect 1066 4048 1103 4064
rect 1137 4064 1139 4082
rect 1173 4082 1211 4098
rect 1173 4064 1175 4082
rect 1137 4048 1175 4064
rect 1209 4064 1211 4082
rect 1245 4064 1246 4098
rect 1209 4048 1246 4064
rect 1066 4025 1246 4048
rect 1066 3991 1067 4025
rect 1101 4014 1139 4025
rect 1101 3991 1103 4014
rect 1066 3980 1103 3991
rect 1137 3991 1139 4014
rect 1173 4014 1211 4025
rect 1173 3991 1175 4014
rect 1137 3980 1175 3991
rect 1209 3991 1211 4014
rect 1245 3991 1246 4025
rect 1209 3980 1246 3991
rect 1066 3952 1246 3980
rect 1066 3918 1067 3952
rect 1101 3946 1139 3952
rect 1101 3918 1103 3946
rect 1066 3912 1103 3918
rect 1137 3918 1139 3946
rect 1173 3946 1211 3952
rect 1173 3918 1175 3946
rect 1137 3912 1175 3918
rect 1209 3918 1211 3946
rect 1245 3918 1246 3952
rect 1209 3912 1246 3918
rect 1066 3879 1246 3912
rect 1066 3845 1067 3879
rect 1101 3878 1139 3879
rect 1101 3845 1103 3878
rect 1066 3844 1103 3845
rect 1137 3845 1139 3878
rect 1173 3878 1211 3879
rect 1173 3845 1175 3878
rect 1137 3844 1175 3845
rect 1209 3845 1211 3878
rect 1245 3845 1246 3879
rect 1209 3844 1246 3845
rect 1066 3810 1246 3844
rect 1066 3806 1103 3810
rect 1066 3772 1067 3806
rect 1101 3776 1103 3806
rect 1137 3806 1175 3810
rect 1137 3776 1139 3806
rect 1101 3772 1139 3776
rect 1173 3776 1175 3806
rect 1209 3806 1246 3810
rect 1209 3776 1211 3806
rect 1173 3772 1211 3776
rect 1245 3772 1246 3806
rect 1066 3742 1246 3772
rect 1066 3733 1103 3742
rect 1066 3699 1067 3733
rect 1101 3708 1103 3733
rect 1137 3733 1175 3742
rect 1137 3708 1139 3733
rect 1101 3699 1139 3708
rect 1173 3708 1175 3733
rect 1209 3733 1246 3742
rect 1209 3708 1211 3733
rect 1173 3699 1211 3708
rect 1245 3699 1246 3733
rect 1066 3674 1246 3699
rect 1066 3660 1103 3674
rect 1066 3626 1067 3660
rect 1101 3640 1103 3660
rect 1137 3660 1175 3674
rect 1137 3640 1139 3660
rect 1101 3626 1139 3640
rect 1173 3640 1175 3660
rect 1209 3660 1246 3674
rect 1209 3640 1211 3660
rect 1173 3626 1211 3640
rect 1245 3626 1246 3660
rect 1066 3606 1246 3626
rect 1066 3587 1103 3606
rect 1066 3553 1067 3587
rect 1101 3572 1103 3587
rect 1137 3587 1175 3606
rect 1137 3572 1139 3587
rect 1101 3553 1139 3572
rect 1173 3572 1175 3587
rect 1209 3587 1246 3606
rect 1209 3572 1211 3587
rect 1173 3553 1211 3572
rect 1245 3553 1246 3587
rect 1066 3538 1246 3553
rect 1066 3514 1103 3538
rect 1066 3480 1067 3514
rect 1101 3504 1103 3514
rect 1137 3514 1175 3538
rect 1137 3504 1139 3514
rect 1101 3480 1139 3504
rect 1173 3504 1175 3514
rect 1209 3514 1246 3538
rect 1209 3504 1211 3514
rect 1173 3480 1211 3504
rect 1245 3480 1246 3514
rect 1066 3470 1246 3480
rect 1066 3441 1103 3470
rect 1066 3407 1067 3441
rect 1101 3436 1103 3441
rect 1137 3441 1175 3470
rect 1137 3436 1139 3441
rect 1101 3407 1139 3436
rect 1173 3436 1175 3441
rect 1209 3441 1246 3470
rect 1209 3436 1211 3441
rect 1173 3407 1211 3436
rect 1245 3407 1246 3441
rect 1066 3402 1246 3407
rect 1066 3368 1103 3402
rect 1137 3368 1175 3402
rect 1209 3368 1246 3402
rect 1066 3334 1067 3368
rect 1101 3334 1139 3368
rect 1173 3334 1211 3368
rect 1245 3334 1246 3368
rect 1066 3300 1103 3334
rect 1137 3300 1175 3334
rect 1209 3300 1246 3334
rect 1066 3295 1246 3300
rect 1066 3261 1067 3295
rect 1101 3266 1139 3295
rect 1101 3261 1103 3266
rect 1066 3232 1103 3261
rect 1137 3261 1139 3266
rect 1173 3266 1211 3295
rect 1173 3261 1175 3266
rect 1137 3232 1175 3261
rect 1209 3261 1211 3266
rect 1245 3261 1246 3295
rect 1209 3232 1246 3261
rect 1066 3222 1246 3232
rect 1066 3188 1067 3222
rect 1101 3198 1139 3222
rect 1101 3188 1103 3198
rect 1066 3164 1103 3188
rect 1137 3188 1139 3198
rect 1173 3198 1211 3222
rect 1173 3188 1175 3198
rect 1137 3164 1175 3188
rect 1209 3188 1211 3198
rect 1245 3188 1246 3222
rect 1209 3164 1246 3188
rect 1066 3149 1246 3164
rect 1066 3115 1067 3149
rect 1101 3115 1139 3149
rect 1173 3115 1211 3149
rect 1245 3115 1246 3149
rect 1066 3076 1246 3115
rect 1066 3042 1067 3076
rect 1101 3042 1139 3076
rect 1173 3042 1211 3076
rect 1245 3042 1246 3076
rect 1066 3003 1246 3042
rect 1066 2969 1067 3003
rect 1101 2969 1139 3003
rect 1173 2969 1211 3003
rect 1245 2969 1246 3003
rect 1066 2930 1246 2969
rect 1066 2896 1067 2930
rect 1101 2896 1139 2930
rect 1173 2896 1211 2930
rect 1245 2896 1246 2930
rect 1066 2857 1246 2896
rect 1066 2823 1067 2857
rect 1101 2823 1139 2857
rect 1173 2823 1211 2857
rect 1245 2823 1246 2857
rect 1066 2784 1246 2823
rect 1066 2750 1067 2784
rect 1101 2750 1139 2784
rect 1173 2750 1211 2784
rect 1245 2750 1246 2784
rect 1066 2711 1246 2750
rect 1066 2677 1067 2711
rect 1101 2677 1139 2711
rect 1173 2677 1211 2711
rect 1245 2677 1246 2711
rect 1066 2638 1246 2677
rect 1066 2604 1067 2638
rect 1101 2604 1139 2638
rect 1173 2604 1211 2638
rect 1245 2604 1246 2638
rect 1066 2565 1246 2604
rect 1066 2531 1067 2565
rect 1101 2531 1139 2565
rect 1173 2531 1211 2565
rect 1245 2531 1246 2565
rect 1066 2492 1246 2531
rect 1066 2458 1067 2492
rect 1101 2482 1139 2492
rect 1101 2458 1103 2482
rect 1066 2448 1103 2458
rect 1137 2458 1139 2482
rect 1173 2482 1211 2492
rect 1173 2458 1175 2482
rect 1137 2448 1175 2458
rect 1209 2458 1211 2482
rect 1245 2458 1246 2492
rect 1209 2448 1246 2458
rect 1066 2419 1246 2448
rect 1066 2385 1067 2419
rect 1101 2414 1139 2419
rect 1101 2385 1103 2414
rect 1066 2380 1103 2385
rect 1137 2385 1139 2414
rect 1173 2414 1211 2419
rect 1173 2385 1175 2414
rect 1137 2380 1175 2385
rect 1209 2385 1211 2414
rect 1245 2385 1246 2419
rect 1209 2380 1246 2385
rect 1066 2346 1246 2380
rect 1066 2312 1067 2346
rect 1101 2312 1103 2346
rect 1137 2312 1139 2346
rect 1173 2312 1175 2346
rect 1209 2312 1211 2346
rect 1245 2312 1246 2346
rect 1066 2278 1246 2312
rect 1066 2273 1103 2278
rect 1066 2239 1067 2273
rect 1101 2244 1103 2273
rect 1137 2273 1175 2278
rect 1137 2244 1139 2273
rect 1101 2239 1139 2244
rect 1173 2244 1175 2273
rect 1209 2273 1246 2278
rect 1209 2244 1211 2273
rect 1173 2239 1211 2244
rect 1245 2239 1246 2273
rect 1066 2210 1246 2239
rect 1066 2200 1103 2210
rect 1066 2166 1067 2200
rect 1101 2176 1103 2200
rect 1137 2200 1175 2210
rect 1137 2176 1139 2200
rect 1101 2166 1139 2176
rect 1173 2176 1175 2200
rect 1209 2200 1246 2210
rect 1209 2176 1211 2200
rect 1173 2166 1211 2176
rect 1245 2166 1246 2200
rect 1066 2142 1246 2166
rect 1066 2126 1103 2142
rect 1066 2092 1067 2126
rect 1101 2108 1103 2126
rect 1137 2126 1175 2142
rect 1137 2108 1139 2126
rect 1101 2092 1139 2108
rect 1173 2108 1175 2126
rect 1209 2126 1246 2142
rect 1209 2108 1211 2126
rect 1173 2092 1211 2108
rect 1245 2092 1246 2126
rect 1066 2074 1246 2092
rect 1066 2052 1103 2074
rect 1066 2018 1067 2052
rect 1101 2040 1103 2052
rect 1137 2052 1175 2074
rect 1137 2040 1139 2052
rect 1101 2018 1139 2040
rect 1173 2040 1175 2052
rect 1209 2052 1246 2074
rect 1209 2040 1211 2052
rect 1173 2018 1211 2040
rect 1245 2018 1246 2052
rect 1066 2006 1246 2018
rect 1066 1978 1103 2006
rect 1066 1944 1067 1978
rect 1101 1972 1103 1978
rect 1137 1978 1175 2006
rect 1137 1972 1139 1978
rect 1101 1944 1139 1972
rect 1173 1972 1175 1978
rect 1209 1978 1246 2006
rect 1209 1972 1211 1978
rect 1173 1944 1211 1972
rect 1245 1944 1246 1978
rect 1066 1938 1246 1944
rect 1066 1904 1103 1938
rect 1137 1904 1175 1938
rect 1209 1904 1246 1938
rect 1066 1870 1067 1904
rect 1101 1870 1139 1904
rect 1173 1870 1211 1904
rect 1245 1870 1246 1904
rect 1066 1836 1103 1870
rect 1137 1836 1175 1870
rect 1209 1836 1246 1870
rect 1066 1830 1246 1836
rect 1066 1796 1067 1830
rect 1101 1802 1139 1830
rect 1101 1796 1103 1802
rect 1066 1768 1103 1796
rect 1137 1796 1139 1802
rect 1173 1802 1211 1830
rect 1173 1796 1175 1802
rect 1137 1768 1175 1796
rect 1209 1796 1211 1802
rect 1245 1796 1246 1830
rect 1209 1768 1246 1796
rect 1066 1756 1246 1768
rect 1066 1722 1067 1756
rect 1101 1734 1139 1756
rect 1101 1722 1103 1734
rect 1066 1700 1103 1722
rect 1137 1722 1139 1734
rect 1173 1734 1211 1756
rect 1173 1722 1175 1734
rect 1137 1700 1175 1722
rect 1209 1722 1211 1734
rect 1245 1722 1246 1756
rect 1209 1700 1246 1722
rect 1066 1682 1246 1700
rect 1066 1648 1067 1682
rect 1101 1666 1139 1682
rect 1101 1648 1103 1666
rect 1066 1632 1103 1648
rect 1137 1648 1139 1666
rect 1173 1666 1211 1682
rect 1173 1648 1175 1666
rect 1137 1632 1175 1648
rect 1209 1648 1211 1666
rect 1245 1648 1246 1682
rect 1209 1632 1246 1648
rect 1066 1608 1246 1632
rect 1066 1574 1067 1608
rect 1101 1598 1139 1608
rect 1101 1574 1103 1598
rect 1066 1564 1103 1574
rect 1137 1574 1139 1598
rect 1173 1598 1211 1608
rect 1173 1574 1175 1598
rect 1137 1564 1175 1574
rect 1209 1574 1211 1598
rect 1245 1574 1246 1608
rect 1209 1564 1246 1574
rect 1066 1548 1246 1564
rect 1311 3104 1431 4200
rect 1873 4308 1993 4324
rect 1873 4274 1916 4308
rect 1950 4274 1993 4308
rect 1873 4234 1993 4274
rect 1873 4200 1916 4234
rect 1950 4200 1993 4234
rect 1311 3070 1354 3104
rect 1388 3070 1431 3104
rect 1311 3026 1431 3070
rect 1311 2992 1354 3026
rect 1388 2992 1431 3026
rect 1311 2948 1431 2992
rect 1311 2914 1354 2948
rect 1388 2914 1431 2948
rect 1311 2870 1431 2914
rect 1311 2836 1354 2870
rect 1388 2836 1431 2870
rect 1311 2792 1431 2836
rect 1311 2758 1354 2792
rect 1388 2758 1431 2792
rect 1311 2713 1431 2758
rect 1311 2679 1354 2713
rect 1388 2679 1431 2713
rect 1311 2634 1431 2679
rect 1311 2600 1354 2634
rect 1388 2600 1431 2634
rect 881 1470 924 1504
rect 958 1470 1001 1504
rect 881 1430 1001 1470
rect 881 1396 924 1430
rect 958 1396 1001 1430
rect 881 1250 1001 1396
rect 881 1216 924 1250
rect 958 1216 1001 1250
rect 881 1178 1001 1216
rect 881 1144 924 1178
rect 958 1144 1001 1178
rect 1311 1504 1431 2600
rect 1533 4092 1635 4118
rect 1669 4092 1771 4118
rect 1533 4082 1563 4092
rect 1741 4082 1771 4092
rect 1533 4014 1563 4048
rect 1741 4014 1771 4048
rect 1533 3946 1563 3980
rect 1741 3946 1771 3980
rect 1533 3878 1563 3912
rect 1741 3878 1771 3912
rect 1533 3810 1563 3844
rect 1741 3810 1771 3844
rect 1533 3742 1563 3776
rect 1741 3742 1771 3776
rect 1533 3674 1563 3708
rect 1741 3674 1771 3708
rect 1533 3606 1563 3640
rect 1741 3606 1771 3640
rect 1533 3538 1563 3572
rect 1741 3538 1771 3572
rect 1533 3470 1563 3504
rect 1741 3470 1771 3504
rect 1533 3402 1563 3436
rect 1741 3402 1771 3436
rect 1533 3334 1563 3368
rect 1741 3334 1771 3368
rect 1533 3266 1563 3300
rect 1741 3266 1771 3300
rect 1533 3198 1563 3232
rect 1741 3198 1771 3232
rect 1567 3164 1635 3194
rect 1669 3164 1737 3194
rect 1533 3148 1635 3164
rect 1669 3148 1771 3164
rect 1533 3108 1771 3148
rect 1533 3074 1563 3108
rect 1597 3074 1635 3108
rect 1669 3074 1707 3108
rect 1741 3074 1771 3108
rect 1533 3044 1771 3074
rect 1533 3028 1601 3044
rect 1533 2994 1563 3028
rect 1597 3010 1601 3028
rect 1635 3028 1669 3044
rect 1597 2994 1635 3010
rect 1703 3028 1771 3044
rect 1703 3010 1707 3028
rect 1669 2994 1707 3010
rect 1741 2994 1771 3028
rect 1533 2974 1771 2994
rect 1533 2948 1601 2974
rect 1533 2914 1563 2948
rect 1597 2940 1601 2948
rect 1635 2948 1669 2974
rect 1597 2914 1635 2940
rect 1703 2948 1771 2974
rect 1703 2940 1707 2948
rect 1669 2914 1707 2940
rect 1741 2914 1771 2948
rect 1533 2904 1771 2914
rect 1533 2870 1601 2904
rect 1635 2870 1669 2904
rect 1703 2870 1771 2904
rect 1533 2868 1771 2870
rect 1533 2834 1563 2868
rect 1597 2834 1635 2868
rect 1669 2834 1707 2868
rect 1741 2834 1771 2868
rect 1533 2800 1601 2834
rect 1635 2800 1669 2834
rect 1703 2800 1771 2834
rect 1533 2788 1771 2800
rect 1533 2754 1563 2788
rect 1597 2764 1635 2788
rect 1597 2754 1601 2764
rect 1533 2730 1601 2754
rect 1669 2764 1707 2788
rect 1635 2730 1669 2754
rect 1703 2754 1707 2764
rect 1741 2754 1771 2788
rect 1703 2730 1771 2754
rect 1533 2708 1771 2730
rect 1533 2674 1563 2708
rect 1597 2694 1635 2708
rect 1597 2674 1601 2694
rect 1533 2660 1601 2674
rect 1669 2694 1707 2708
rect 1635 2660 1669 2674
rect 1703 2674 1707 2694
rect 1741 2674 1771 2708
rect 1703 2660 1771 2674
rect 1533 2628 1771 2660
rect 1533 2594 1563 2628
rect 1597 2594 1635 2628
rect 1669 2594 1707 2628
rect 1741 2594 1771 2628
rect 1533 2556 1771 2594
rect 1533 2540 1635 2556
rect 1669 2540 1771 2556
rect 1567 2518 1635 2540
rect 1669 2518 1737 2540
rect 1533 2472 1563 2506
rect 1741 2472 1771 2506
rect 1533 2404 1563 2438
rect 1741 2404 1771 2438
rect 1533 2336 1563 2370
rect 1741 2336 1771 2370
rect 1533 2268 1563 2302
rect 1741 2268 1771 2302
rect 1533 2200 1563 2234
rect 1741 2200 1771 2234
rect 1533 2132 1563 2166
rect 1741 2132 1771 2166
rect 1533 2064 1563 2098
rect 1741 2064 1771 2098
rect 1533 1996 1563 2030
rect 1741 1996 1771 2030
rect 1533 1928 1563 1962
rect 1741 1928 1771 1962
rect 1533 1860 1563 1894
rect 1741 1860 1771 1894
rect 1533 1792 1563 1826
rect 1741 1792 1771 1826
rect 1533 1724 1563 1758
rect 1741 1724 1771 1758
rect 1533 1656 1563 1690
rect 1741 1656 1771 1690
rect 1533 1620 1563 1622
rect 1741 1620 1771 1622
rect 1533 1586 1635 1620
rect 1669 1586 1771 1620
rect 1533 1536 1771 1586
rect 1873 3104 1993 4200
rect 2303 4308 2423 4324
rect 2303 4274 2346 4308
rect 2380 4274 2423 4308
rect 2303 4234 2423 4274
rect 2303 4200 2346 4234
rect 2380 4200 2423 4234
rect 1873 3070 1916 3104
rect 1950 3070 1993 3104
rect 1873 3026 1993 3070
rect 1873 2992 1916 3026
rect 1950 2992 1993 3026
rect 1873 2948 1993 2992
rect 1873 2914 1916 2948
rect 1950 2914 1993 2948
rect 1873 2870 1993 2914
rect 1873 2836 1916 2870
rect 1950 2836 1993 2870
rect 1873 2792 1993 2836
rect 1873 2758 1916 2792
rect 1950 2758 1993 2792
rect 1873 2713 1993 2758
rect 1873 2679 1916 2713
rect 1950 2679 1993 2713
rect 1873 2634 1993 2679
rect 1873 2600 1916 2634
rect 1950 2600 1993 2634
rect 1311 1470 1354 1504
rect 1388 1470 1431 1504
rect 1311 1430 1431 1470
rect 1311 1396 1354 1430
rect 1388 1396 1431 1430
rect 1311 1250 1431 1396
rect 1311 1144 1318 1250
rect 1424 1144 1431 1250
rect 1873 1504 1993 2600
rect 2058 4064 2059 4098
rect 2093 4082 2131 4098
rect 2093 4064 2095 4082
rect 2058 4048 2095 4064
rect 2129 4064 2131 4082
rect 2165 4082 2203 4098
rect 2165 4064 2167 4082
rect 2129 4048 2167 4064
rect 2201 4064 2203 4082
rect 2237 4064 2238 4098
rect 2201 4048 2238 4064
rect 2058 4025 2238 4048
rect 2058 3991 2059 4025
rect 2093 4014 2131 4025
rect 2093 3991 2095 4014
rect 2058 3980 2095 3991
rect 2129 3991 2131 4014
rect 2165 4014 2203 4025
rect 2165 3991 2167 4014
rect 2129 3980 2167 3991
rect 2201 3991 2203 4014
rect 2237 3991 2238 4025
rect 2201 3980 2238 3991
rect 2058 3952 2238 3980
rect 2058 3918 2059 3952
rect 2093 3946 2131 3952
rect 2093 3918 2095 3946
rect 2058 3912 2095 3918
rect 2129 3918 2131 3946
rect 2165 3946 2203 3952
rect 2165 3918 2167 3946
rect 2129 3912 2167 3918
rect 2201 3918 2203 3946
rect 2237 3918 2238 3952
rect 2201 3912 2238 3918
rect 2058 3879 2238 3912
rect 2058 3845 2059 3879
rect 2093 3878 2131 3879
rect 2093 3845 2095 3878
rect 2058 3844 2095 3845
rect 2129 3845 2131 3878
rect 2165 3878 2203 3879
rect 2165 3845 2167 3878
rect 2129 3844 2167 3845
rect 2201 3845 2203 3878
rect 2237 3845 2238 3879
rect 2201 3844 2238 3845
rect 2058 3810 2238 3844
rect 2058 3806 2095 3810
rect 2058 3772 2059 3806
rect 2093 3776 2095 3806
rect 2129 3806 2167 3810
rect 2129 3776 2131 3806
rect 2093 3772 2131 3776
rect 2165 3776 2167 3806
rect 2201 3806 2238 3810
rect 2201 3776 2203 3806
rect 2165 3772 2203 3776
rect 2237 3772 2238 3806
rect 2058 3742 2238 3772
rect 2058 3733 2095 3742
rect 2058 3699 2059 3733
rect 2093 3708 2095 3733
rect 2129 3733 2167 3742
rect 2129 3708 2131 3733
rect 2093 3699 2131 3708
rect 2165 3708 2167 3733
rect 2201 3733 2238 3742
rect 2201 3708 2203 3733
rect 2165 3699 2203 3708
rect 2237 3699 2238 3733
rect 2058 3674 2238 3699
rect 2058 3660 2095 3674
rect 2058 3626 2059 3660
rect 2093 3640 2095 3660
rect 2129 3660 2167 3674
rect 2129 3640 2131 3660
rect 2093 3626 2131 3640
rect 2165 3640 2167 3660
rect 2201 3660 2238 3674
rect 2201 3640 2203 3660
rect 2165 3626 2203 3640
rect 2237 3626 2238 3660
rect 2058 3606 2238 3626
rect 2058 3587 2095 3606
rect 2058 3553 2059 3587
rect 2093 3572 2095 3587
rect 2129 3587 2167 3606
rect 2129 3572 2131 3587
rect 2093 3553 2131 3572
rect 2165 3572 2167 3587
rect 2201 3587 2238 3606
rect 2201 3572 2203 3587
rect 2165 3553 2203 3572
rect 2237 3553 2238 3587
rect 2058 3538 2238 3553
rect 2058 3514 2095 3538
rect 2058 3480 2059 3514
rect 2093 3504 2095 3514
rect 2129 3514 2167 3538
rect 2129 3504 2131 3514
rect 2093 3480 2131 3504
rect 2165 3504 2167 3514
rect 2201 3514 2238 3538
rect 2201 3504 2203 3514
rect 2165 3480 2203 3504
rect 2237 3480 2238 3514
rect 2058 3470 2238 3480
rect 2058 3441 2095 3470
rect 2058 3407 2059 3441
rect 2093 3436 2095 3441
rect 2129 3441 2167 3470
rect 2129 3436 2131 3441
rect 2093 3407 2131 3436
rect 2165 3436 2167 3441
rect 2201 3441 2238 3470
rect 2201 3436 2203 3441
rect 2165 3407 2203 3436
rect 2237 3407 2238 3441
rect 2058 3402 2238 3407
rect 2058 3368 2095 3402
rect 2129 3368 2167 3402
rect 2201 3368 2238 3402
rect 2058 3334 2059 3368
rect 2093 3334 2131 3368
rect 2165 3334 2203 3368
rect 2237 3334 2238 3368
rect 2058 3300 2095 3334
rect 2129 3300 2167 3334
rect 2201 3300 2238 3334
rect 2058 3295 2238 3300
rect 2058 3261 2059 3295
rect 2093 3266 2131 3295
rect 2093 3261 2095 3266
rect 2058 3232 2095 3261
rect 2129 3261 2131 3266
rect 2165 3266 2203 3295
rect 2165 3261 2167 3266
rect 2129 3232 2167 3261
rect 2201 3261 2203 3266
rect 2237 3261 2238 3295
rect 2201 3232 2238 3261
rect 2058 3222 2238 3232
rect 2058 3188 2059 3222
rect 2093 3198 2131 3222
rect 2093 3188 2095 3198
rect 2058 3164 2095 3188
rect 2129 3188 2131 3198
rect 2165 3198 2203 3222
rect 2165 3188 2167 3198
rect 2129 3164 2167 3188
rect 2201 3188 2203 3198
rect 2237 3188 2238 3222
rect 2201 3164 2238 3188
rect 2058 3149 2238 3164
rect 2058 3115 2059 3149
rect 2093 3115 2131 3149
rect 2165 3115 2203 3149
rect 2237 3115 2238 3149
rect 2058 3076 2238 3115
rect 2058 3042 2059 3076
rect 2093 3042 2131 3076
rect 2165 3042 2203 3076
rect 2237 3042 2238 3076
rect 2058 3003 2238 3042
rect 2058 2969 2059 3003
rect 2093 2969 2131 3003
rect 2165 2969 2203 3003
rect 2237 2969 2238 3003
rect 2058 2930 2238 2969
rect 2058 2896 2059 2930
rect 2093 2896 2131 2930
rect 2165 2896 2203 2930
rect 2237 2896 2238 2930
rect 2058 2857 2238 2896
rect 2058 2823 2059 2857
rect 2093 2823 2131 2857
rect 2165 2823 2203 2857
rect 2237 2823 2238 2857
rect 2058 2784 2238 2823
rect 2058 2750 2059 2784
rect 2093 2750 2131 2784
rect 2165 2750 2203 2784
rect 2237 2750 2238 2784
rect 2058 2711 2238 2750
rect 2058 2677 2059 2711
rect 2093 2677 2131 2711
rect 2165 2677 2203 2711
rect 2237 2677 2238 2711
rect 2058 2638 2238 2677
rect 2058 2604 2059 2638
rect 2093 2604 2131 2638
rect 2165 2604 2203 2638
rect 2237 2604 2238 2638
rect 2058 2565 2238 2604
rect 2058 2531 2059 2565
rect 2093 2531 2131 2565
rect 2165 2531 2203 2565
rect 2237 2531 2238 2565
rect 2058 2492 2238 2531
rect 2058 2458 2059 2492
rect 2093 2482 2131 2492
rect 2093 2458 2095 2482
rect 2058 2448 2095 2458
rect 2129 2458 2131 2482
rect 2165 2482 2203 2492
rect 2165 2458 2167 2482
rect 2129 2448 2167 2458
rect 2201 2458 2203 2482
rect 2237 2458 2238 2492
rect 2201 2448 2238 2458
rect 2058 2419 2238 2448
rect 2058 2385 2059 2419
rect 2093 2414 2131 2419
rect 2093 2385 2095 2414
rect 2058 2380 2095 2385
rect 2129 2385 2131 2414
rect 2165 2414 2203 2419
rect 2165 2385 2167 2414
rect 2129 2380 2167 2385
rect 2201 2385 2203 2414
rect 2237 2385 2238 2419
rect 2201 2380 2238 2385
rect 2058 2346 2238 2380
rect 2058 2312 2059 2346
rect 2093 2312 2095 2346
rect 2129 2312 2131 2346
rect 2165 2312 2167 2346
rect 2201 2312 2203 2346
rect 2237 2312 2238 2346
rect 2058 2278 2238 2312
rect 2058 2273 2095 2278
rect 2058 2239 2059 2273
rect 2093 2244 2095 2273
rect 2129 2273 2167 2278
rect 2129 2244 2131 2273
rect 2093 2239 2131 2244
rect 2165 2244 2167 2273
rect 2201 2273 2238 2278
rect 2201 2244 2203 2273
rect 2165 2239 2203 2244
rect 2237 2239 2238 2273
rect 2058 2210 2238 2239
rect 2058 2200 2095 2210
rect 2058 2166 2059 2200
rect 2093 2176 2095 2200
rect 2129 2200 2167 2210
rect 2129 2176 2131 2200
rect 2093 2166 2131 2176
rect 2165 2176 2167 2200
rect 2201 2200 2238 2210
rect 2201 2176 2203 2200
rect 2165 2166 2203 2176
rect 2237 2166 2238 2200
rect 2058 2142 2238 2166
rect 2058 2126 2095 2142
rect 2058 2092 2059 2126
rect 2093 2108 2095 2126
rect 2129 2126 2167 2142
rect 2129 2108 2131 2126
rect 2093 2092 2131 2108
rect 2165 2108 2167 2126
rect 2201 2126 2238 2142
rect 2201 2108 2203 2126
rect 2165 2092 2203 2108
rect 2237 2092 2238 2126
rect 2058 2074 2238 2092
rect 2058 2052 2095 2074
rect 2058 2018 2059 2052
rect 2093 2040 2095 2052
rect 2129 2052 2167 2074
rect 2129 2040 2131 2052
rect 2093 2018 2131 2040
rect 2165 2040 2167 2052
rect 2201 2052 2238 2074
rect 2201 2040 2203 2052
rect 2165 2018 2203 2040
rect 2237 2018 2238 2052
rect 2058 2006 2238 2018
rect 2058 1978 2095 2006
rect 2058 1944 2059 1978
rect 2093 1972 2095 1978
rect 2129 1978 2167 2006
rect 2129 1972 2131 1978
rect 2093 1944 2131 1972
rect 2165 1972 2167 1978
rect 2201 1978 2238 2006
rect 2201 1972 2203 1978
rect 2165 1944 2203 1972
rect 2237 1944 2238 1978
rect 2058 1938 2238 1944
rect 2058 1904 2095 1938
rect 2129 1904 2167 1938
rect 2201 1904 2238 1938
rect 2058 1870 2059 1904
rect 2093 1870 2131 1904
rect 2165 1870 2203 1904
rect 2237 1870 2238 1904
rect 2058 1836 2095 1870
rect 2129 1836 2167 1870
rect 2201 1836 2238 1870
rect 2058 1830 2238 1836
rect 2058 1796 2059 1830
rect 2093 1802 2131 1830
rect 2093 1796 2095 1802
rect 2058 1768 2095 1796
rect 2129 1796 2131 1802
rect 2165 1802 2203 1830
rect 2165 1796 2167 1802
rect 2129 1768 2167 1796
rect 2201 1796 2203 1802
rect 2237 1796 2238 1830
rect 2201 1768 2238 1796
rect 2058 1756 2238 1768
rect 2058 1722 2059 1756
rect 2093 1734 2131 1756
rect 2093 1722 2095 1734
rect 2058 1700 2095 1722
rect 2129 1722 2131 1734
rect 2165 1734 2203 1756
rect 2165 1722 2167 1734
rect 2129 1700 2167 1722
rect 2201 1722 2203 1734
rect 2237 1722 2238 1756
rect 2201 1700 2238 1722
rect 2058 1682 2238 1700
rect 2058 1648 2059 1682
rect 2093 1666 2131 1682
rect 2093 1648 2095 1666
rect 2058 1632 2095 1648
rect 2129 1648 2131 1666
rect 2165 1666 2203 1682
rect 2165 1648 2167 1666
rect 2129 1632 2167 1648
rect 2201 1648 2203 1666
rect 2237 1648 2238 1682
rect 2201 1632 2238 1648
rect 2058 1608 2238 1632
rect 2058 1574 2059 1608
rect 2093 1598 2131 1608
rect 2093 1574 2095 1598
rect 2058 1564 2095 1574
rect 2129 1574 2131 1598
rect 2165 1598 2203 1608
rect 2165 1574 2167 1598
rect 2129 1564 2167 1574
rect 2201 1574 2203 1598
rect 2237 1574 2238 1608
rect 2201 1564 2238 1574
rect 2058 1548 2238 1564
rect 2303 3104 2423 4200
rect 2865 4308 2985 4324
rect 2865 4274 2908 4308
rect 2942 4274 2985 4308
rect 2865 4234 2985 4274
rect 2865 4200 2908 4234
rect 2942 4200 2985 4234
rect 2303 3070 2346 3104
rect 2380 3070 2423 3104
rect 2303 3026 2423 3070
rect 2303 2992 2346 3026
rect 2380 2992 2423 3026
rect 2303 2948 2423 2992
rect 2303 2914 2346 2948
rect 2380 2914 2423 2948
rect 2303 2870 2423 2914
rect 2303 2836 2346 2870
rect 2380 2836 2423 2870
rect 2303 2792 2423 2836
rect 2303 2758 2346 2792
rect 2380 2758 2423 2792
rect 2303 2713 2423 2758
rect 2303 2679 2346 2713
rect 2380 2679 2423 2713
rect 2303 2634 2423 2679
rect 2303 2600 2346 2634
rect 2380 2600 2423 2634
rect 1873 1470 1916 1504
rect 1950 1470 1993 1504
rect 1873 1430 1993 1470
rect 1873 1396 1916 1430
rect 1950 1396 1993 1430
rect 1873 1250 1993 1396
rect 1873 1144 1880 1250
rect 1986 1144 1993 1250
rect 2303 1504 2423 2600
rect 2525 4092 2627 4118
rect 2661 4092 2763 4118
rect 2525 4082 2555 4092
rect 2733 4082 2763 4092
rect 2525 4014 2555 4048
rect 2733 4014 2763 4048
rect 2525 3946 2555 3980
rect 2733 3946 2763 3980
rect 2525 3878 2555 3912
rect 2733 3878 2763 3912
rect 2525 3810 2555 3844
rect 2733 3810 2763 3844
rect 2525 3742 2555 3776
rect 2733 3742 2763 3776
rect 2525 3674 2555 3708
rect 2733 3674 2763 3708
rect 2525 3606 2555 3640
rect 2733 3606 2763 3640
rect 2525 3538 2555 3572
rect 2733 3538 2763 3572
rect 2525 3470 2555 3504
rect 2733 3470 2763 3504
rect 2525 3402 2555 3436
rect 2733 3402 2763 3436
rect 2525 3334 2555 3368
rect 2733 3334 2763 3368
rect 2525 3266 2555 3300
rect 2733 3266 2763 3300
rect 2525 3198 2555 3232
rect 2733 3198 2763 3232
rect 2559 3164 2627 3194
rect 2661 3164 2729 3194
rect 2525 3148 2627 3164
rect 2661 3148 2763 3164
rect 2525 3108 2763 3148
rect 2525 3074 2555 3108
rect 2589 3074 2627 3108
rect 2661 3074 2699 3108
rect 2733 3074 2763 3108
rect 2525 3044 2763 3074
rect 2525 3028 2593 3044
rect 2525 2994 2555 3028
rect 2589 3010 2593 3028
rect 2627 3028 2661 3044
rect 2589 2994 2627 3010
rect 2695 3028 2763 3044
rect 2695 3010 2699 3028
rect 2661 2994 2699 3010
rect 2733 2994 2763 3028
rect 2525 2974 2763 2994
rect 2525 2948 2593 2974
rect 2525 2914 2555 2948
rect 2589 2940 2593 2948
rect 2627 2948 2661 2974
rect 2589 2914 2627 2940
rect 2695 2948 2763 2974
rect 2695 2940 2699 2948
rect 2661 2914 2699 2940
rect 2733 2914 2763 2948
rect 2525 2904 2763 2914
rect 2525 2870 2593 2904
rect 2627 2870 2661 2904
rect 2695 2870 2763 2904
rect 2525 2868 2763 2870
rect 2525 2834 2555 2868
rect 2589 2834 2627 2868
rect 2661 2834 2699 2868
rect 2733 2834 2763 2868
rect 2525 2800 2593 2834
rect 2627 2800 2661 2834
rect 2695 2800 2763 2834
rect 2525 2788 2763 2800
rect 2525 2754 2555 2788
rect 2589 2764 2627 2788
rect 2589 2754 2593 2764
rect 2525 2730 2593 2754
rect 2661 2764 2699 2788
rect 2627 2730 2661 2754
rect 2695 2754 2699 2764
rect 2733 2754 2763 2788
rect 2695 2730 2763 2754
rect 2525 2708 2763 2730
rect 2525 2674 2555 2708
rect 2589 2694 2627 2708
rect 2589 2674 2593 2694
rect 2525 2660 2593 2674
rect 2661 2694 2699 2708
rect 2627 2660 2661 2674
rect 2695 2674 2699 2694
rect 2733 2674 2763 2708
rect 2695 2660 2763 2674
rect 2525 2628 2763 2660
rect 2525 2594 2555 2628
rect 2589 2594 2627 2628
rect 2661 2594 2699 2628
rect 2733 2594 2763 2628
rect 2525 2556 2763 2594
rect 2525 2540 2627 2556
rect 2661 2540 2763 2556
rect 2559 2518 2627 2540
rect 2661 2518 2729 2540
rect 2525 2472 2555 2506
rect 2733 2472 2763 2506
rect 2525 2404 2555 2438
rect 2733 2404 2763 2438
rect 2525 2336 2555 2370
rect 2733 2336 2763 2370
rect 2525 2268 2555 2302
rect 2733 2268 2763 2302
rect 2525 2200 2555 2234
rect 2733 2200 2763 2234
rect 2525 2132 2555 2166
rect 2733 2132 2763 2166
rect 2525 2064 2555 2098
rect 2733 2064 2763 2098
rect 2525 1996 2555 2030
rect 2733 1996 2763 2030
rect 2525 1928 2555 1962
rect 2733 1928 2763 1962
rect 2525 1860 2555 1894
rect 2733 1860 2763 1894
rect 2525 1792 2555 1826
rect 2733 1792 2763 1826
rect 2525 1724 2555 1758
rect 2733 1724 2763 1758
rect 2525 1656 2555 1690
rect 2733 1656 2763 1690
rect 2525 1620 2555 1622
rect 2733 1620 2763 1622
rect 2525 1586 2627 1620
rect 2661 1586 2763 1620
rect 2525 1536 2763 1586
rect 2865 3104 2985 4200
rect 3295 4308 3415 4324
rect 3295 4274 3338 4308
rect 3372 4274 3415 4308
rect 3295 4234 3415 4274
rect 3295 4200 3338 4234
rect 3372 4200 3415 4234
rect 2865 3070 2908 3104
rect 2942 3070 2985 3104
rect 2865 3026 2985 3070
rect 2865 2992 2908 3026
rect 2942 2992 2985 3026
rect 2865 2948 2985 2992
rect 2865 2914 2908 2948
rect 2942 2914 2985 2948
rect 2865 2870 2985 2914
rect 2865 2836 2908 2870
rect 2942 2836 2985 2870
rect 2865 2792 2985 2836
rect 2865 2758 2908 2792
rect 2942 2758 2985 2792
rect 2865 2713 2985 2758
rect 2865 2679 2908 2713
rect 2942 2679 2985 2713
rect 2865 2634 2985 2679
rect 2865 2600 2908 2634
rect 2942 2600 2985 2634
rect 2303 1470 2346 1504
rect 2380 1470 2423 1504
rect 2303 1430 2423 1470
rect 2303 1396 2346 1430
rect 2380 1396 2423 1430
rect 2303 1250 2423 1396
rect 2303 1144 2310 1250
rect 2416 1144 2423 1250
rect 2865 1504 2985 2600
rect 3050 4064 3051 4098
rect 3085 4082 3123 4098
rect 3085 4064 3087 4082
rect 3050 4048 3087 4064
rect 3121 4064 3123 4082
rect 3157 4082 3195 4098
rect 3157 4064 3159 4082
rect 3121 4048 3159 4064
rect 3193 4064 3195 4082
rect 3229 4064 3230 4098
rect 3193 4048 3230 4064
rect 3050 4025 3230 4048
rect 3050 3991 3051 4025
rect 3085 4014 3123 4025
rect 3085 3991 3087 4014
rect 3050 3980 3087 3991
rect 3121 3991 3123 4014
rect 3157 4014 3195 4025
rect 3157 3991 3159 4014
rect 3121 3980 3159 3991
rect 3193 3991 3195 4014
rect 3229 3991 3230 4025
rect 3193 3980 3230 3991
rect 3050 3952 3230 3980
rect 3050 3918 3051 3952
rect 3085 3946 3123 3952
rect 3085 3918 3087 3946
rect 3050 3912 3087 3918
rect 3121 3918 3123 3946
rect 3157 3946 3195 3952
rect 3157 3918 3159 3946
rect 3121 3912 3159 3918
rect 3193 3918 3195 3946
rect 3229 3918 3230 3952
rect 3193 3912 3230 3918
rect 3050 3879 3230 3912
rect 3050 3845 3051 3879
rect 3085 3878 3123 3879
rect 3085 3845 3087 3878
rect 3050 3844 3087 3845
rect 3121 3845 3123 3878
rect 3157 3878 3195 3879
rect 3157 3845 3159 3878
rect 3121 3844 3159 3845
rect 3193 3845 3195 3878
rect 3229 3845 3230 3879
rect 3193 3844 3230 3845
rect 3050 3810 3230 3844
rect 3050 3806 3087 3810
rect 3050 3772 3051 3806
rect 3085 3776 3087 3806
rect 3121 3806 3159 3810
rect 3121 3776 3123 3806
rect 3085 3772 3123 3776
rect 3157 3776 3159 3806
rect 3193 3806 3230 3810
rect 3193 3776 3195 3806
rect 3157 3772 3195 3776
rect 3229 3772 3230 3806
rect 3050 3742 3230 3772
rect 3050 3733 3087 3742
rect 3050 3699 3051 3733
rect 3085 3708 3087 3733
rect 3121 3733 3159 3742
rect 3121 3708 3123 3733
rect 3085 3699 3123 3708
rect 3157 3708 3159 3733
rect 3193 3733 3230 3742
rect 3193 3708 3195 3733
rect 3157 3699 3195 3708
rect 3229 3699 3230 3733
rect 3050 3674 3230 3699
rect 3050 3660 3087 3674
rect 3050 3626 3051 3660
rect 3085 3640 3087 3660
rect 3121 3660 3159 3674
rect 3121 3640 3123 3660
rect 3085 3626 3123 3640
rect 3157 3640 3159 3660
rect 3193 3660 3230 3674
rect 3193 3640 3195 3660
rect 3157 3626 3195 3640
rect 3229 3626 3230 3660
rect 3050 3606 3230 3626
rect 3050 3587 3087 3606
rect 3050 3553 3051 3587
rect 3085 3572 3087 3587
rect 3121 3587 3159 3606
rect 3121 3572 3123 3587
rect 3085 3553 3123 3572
rect 3157 3572 3159 3587
rect 3193 3587 3230 3606
rect 3193 3572 3195 3587
rect 3157 3553 3195 3572
rect 3229 3553 3230 3587
rect 3050 3538 3230 3553
rect 3050 3514 3087 3538
rect 3050 3480 3051 3514
rect 3085 3504 3087 3514
rect 3121 3514 3159 3538
rect 3121 3504 3123 3514
rect 3085 3480 3123 3504
rect 3157 3504 3159 3514
rect 3193 3514 3230 3538
rect 3193 3504 3195 3514
rect 3157 3480 3195 3504
rect 3229 3480 3230 3514
rect 3050 3470 3230 3480
rect 3050 3441 3087 3470
rect 3050 3407 3051 3441
rect 3085 3436 3087 3441
rect 3121 3441 3159 3470
rect 3121 3436 3123 3441
rect 3085 3407 3123 3436
rect 3157 3436 3159 3441
rect 3193 3441 3230 3470
rect 3193 3436 3195 3441
rect 3157 3407 3195 3436
rect 3229 3407 3230 3441
rect 3050 3402 3230 3407
rect 3050 3368 3087 3402
rect 3121 3368 3159 3402
rect 3193 3368 3230 3402
rect 3050 3334 3051 3368
rect 3085 3334 3123 3368
rect 3157 3334 3195 3368
rect 3229 3334 3230 3368
rect 3050 3300 3087 3334
rect 3121 3300 3159 3334
rect 3193 3300 3230 3334
rect 3050 3295 3230 3300
rect 3050 3261 3051 3295
rect 3085 3266 3123 3295
rect 3085 3261 3087 3266
rect 3050 3232 3087 3261
rect 3121 3261 3123 3266
rect 3157 3266 3195 3295
rect 3157 3261 3159 3266
rect 3121 3232 3159 3261
rect 3193 3261 3195 3266
rect 3229 3261 3230 3295
rect 3193 3232 3230 3261
rect 3050 3222 3230 3232
rect 3050 3188 3051 3222
rect 3085 3198 3123 3222
rect 3085 3188 3087 3198
rect 3050 3164 3087 3188
rect 3121 3188 3123 3198
rect 3157 3198 3195 3222
rect 3157 3188 3159 3198
rect 3121 3164 3159 3188
rect 3193 3188 3195 3198
rect 3229 3188 3230 3222
rect 3193 3164 3230 3188
rect 3050 3149 3230 3164
rect 3050 3115 3051 3149
rect 3085 3115 3123 3149
rect 3157 3115 3195 3149
rect 3229 3115 3230 3149
rect 3050 3076 3230 3115
rect 3050 3042 3051 3076
rect 3085 3042 3123 3076
rect 3157 3042 3195 3076
rect 3229 3042 3230 3076
rect 3050 3003 3230 3042
rect 3050 2969 3051 3003
rect 3085 2969 3123 3003
rect 3157 2969 3195 3003
rect 3229 2969 3230 3003
rect 3050 2930 3230 2969
rect 3050 2896 3051 2930
rect 3085 2896 3123 2930
rect 3157 2896 3195 2930
rect 3229 2896 3230 2930
rect 3050 2857 3230 2896
rect 3050 2823 3051 2857
rect 3085 2823 3123 2857
rect 3157 2823 3195 2857
rect 3229 2823 3230 2857
rect 3050 2784 3230 2823
rect 3050 2750 3051 2784
rect 3085 2750 3123 2784
rect 3157 2750 3195 2784
rect 3229 2750 3230 2784
rect 3050 2711 3230 2750
rect 3050 2677 3051 2711
rect 3085 2677 3123 2711
rect 3157 2677 3195 2711
rect 3229 2677 3230 2711
rect 3050 2638 3230 2677
rect 3050 2604 3051 2638
rect 3085 2604 3123 2638
rect 3157 2604 3195 2638
rect 3229 2604 3230 2638
rect 3050 2565 3230 2604
rect 3050 2531 3051 2565
rect 3085 2531 3123 2565
rect 3157 2531 3195 2565
rect 3229 2531 3230 2565
rect 3050 2492 3230 2531
rect 3050 2458 3051 2492
rect 3085 2482 3123 2492
rect 3085 2458 3087 2482
rect 3050 2448 3087 2458
rect 3121 2458 3123 2482
rect 3157 2482 3195 2492
rect 3157 2458 3159 2482
rect 3121 2448 3159 2458
rect 3193 2458 3195 2482
rect 3229 2458 3230 2492
rect 3193 2448 3230 2458
rect 3050 2419 3230 2448
rect 3050 2385 3051 2419
rect 3085 2414 3123 2419
rect 3085 2385 3087 2414
rect 3050 2380 3087 2385
rect 3121 2385 3123 2414
rect 3157 2414 3195 2419
rect 3157 2385 3159 2414
rect 3121 2380 3159 2385
rect 3193 2385 3195 2414
rect 3229 2385 3230 2419
rect 3193 2380 3230 2385
rect 3050 2346 3230 2380
rect 3050 2312 3051 2346
rect 3085 2312 3087 2346
rect 3121 2312 3123 2346
rect 3157 2312 3159 2346
rect 3193 2312 3195 2346
rect 3229 2312 3230 2346
rect 3050 2278 3230 2312
rect 3050 2273 3087 2278
rect 3050 2239 3051 2273
rect 3085 2244 3087 2273
rect 3121 2273 3159 2278
rect 3121 2244 3123 2273
rect 3085 2239 3123 2244
rect 3157 2244 3159 2273
rect 3193 2273 3230 2278
rect 3193 2244 3195 2273
rect 3157 2239 3195 2244
rect 3229 2239 3230 2273
rect 3050 2210 3230 2239
rect 3050 2200 3087 2210
rect 3050 2166 3051 2200
rect 3085 2176 3087 2200
rect 3121 2200 3159 2210
rect 3121 2176 3123 2200
rect 3085 2166 3123 2176
rect 3157 2176 3159 2200
rect 3193 2200 3230 2210
rect 3193 2176 3195 2200
rect 3157 2166 3195 2176
rect 3229 2166 3230 2200
rect 3050 2142 3230 2166
rect 3050 2126 3087 2142
rect 3050 2092 3051 2126
rect 3085 2108 3087 2126
rect 3121 2126 3159 2142
rect 3121 2108 3123 2126
rect 3085 2092 3123 2108
rect 3157 2108 3159 2126
rect 3193 2126 3230 2142
rect 3193 2108 3195 2126
rect 3157 2092 3195 2108
rect 3229 2092 3230 2126
rect 3050 2074 3230 2092
rect 3050 2052 3087 2074
rect 3050 2018 3051 2052
rect 3085 2040 3087 2052
rect 3121 2052 3159 2074
rect 3121 2040 3123 2052
rect 3085 2018 3123 2040
rect 3157 2040 3159 2052
rect 3193 2052 3230 2074
rect 3193 2040 3195 2052
rect 3157 2018 3195 2040
rect 3229 2018 3230 2052
rect 3050 2006 3230 2018
rect 3050 1978 3087 2006
rect 3050 1944 3051 1978
rect 3085 1972 3087 1978
rect 3121 1978 3159 2006
rect 3121 1972 3123 1978
rect 3085 1944 3123 1972
rect 3157 1972 3159 1978
rect 3193 1978 3230 2006
rect 3193 1972 3195 1978
rect 3157 1944 3195 1972
rect 3229 1944 3230 1978
rect 3050 1938 3230 1944
rect 3050 1904 3087 1938
rect 3121 1904 3159 1938
rect 3193 1904 3230 1938
rect 3050 1870 3051 1904
rect 3085 1870 3123 1904
rect 3157 1870 3195 1904
rect 3229 1870 3230 1904
rect 3050 1836 3087 1870
rect 3121 1836 3159 1870
rect 3193 1836 3230 1870
rect 3050 1830 3230 1836
rect 3050 1796 3051 1830
rect 3085 1802 3123 1830
rect 3085 1796 3087 1802
rect 3050 1768 3087 1796
rect 3121 1796 3123 1802
rect 3157 1802 3195 1830
rect 3157 1796 3159 1802
rect 3121 1768 3159 1796
rect 3193 1796 3195 1802
rect 3229 1796 3230 1830
rect 3193 1768 3230 1796
rect 3050 1756 3230 1768
rect 3050 1722 3051 1756
rect 3085 1734 3123 1756
rect 3085 1722 3087 1734
rect 3050 1700 3087 1722
rect 3121 1722 3123 1734
rect 3157 1734 3195 1756
rect 3157 1722 3159 1734
rect 3121 1700 3159 1722
rect 3193 1722 3195 1734
rect 3229 1722 3230 1756
rect 3193 1700 3230 1722
rect 3050 1682 3230 1700
rect 3050 1648 3051 1682
rect 3085 1666 3123 1682
rect 3085 1648 3087 1666
rect 3050 1632 3087 1648
rect 3121 1648 3123 1666
rect 3157 1666 3195 1682
rect 3157 1648 3159 1666
rect 3121 1632 3159 1648
rect 3193 1648 3195 1666
rect 3229 1648 3230 1682
rect 3193 1632 3230 1648
rect 3050 1608 3230 1632
rect 3050 1574 3051 1608
rect 3085 1598 3123 1608
rect 3085 1574 3087 1598
rect 3050 1564 3087 1574
rect 3121 1574 3123 1598
rect 3157 1598 3195 1608
rect 3157 1574 3159 1598
rect 3121 1564 3159 1574
rect 3193 1574 3195 1598
rect 3229 1574 3230 1608
rect 3193 1564 3230 1574
rect 3050 1548 3230 1564
rect 3295 3104 3415 4200
rect 3857 4308 3977 4324
rect 3857 4274 3900 4308
rect 3934 4274 3977 4308
rect 3857 4234 3977 4274
rect 3857 4200 3900 4234
rect 3934 4200 3977 4234
rect 3295 3070 3338 3104
rect 3372 3070 3415 3104
rect 3295 3026 3415 3070
rect 3295 2992 3338 3026
rect 3372 2992 3415 3026
rect 3295 2948 3415 2992
rect 3295 2914 3338 2948
rect 3372 2914 3415 2948
rect 3295 2870 3415 2914
rect 3295 2836 3338 2870
rect 3372 2836 3415 2870
rect 3295 2792 3415 2836
rect 3295 2758 3338 2792
rect 3372 2758 3415 2792
rect 3295 2713 3415 2758
rect 3295 2679 3338 2713
rect 3372 2679 3415 2713
rect 3295 2634 3415 2679
rect 3295 2600 3338 2634
rect 3372 2600 3415 2634
rect 2865 1470 2908 1504
rect 2942 1470 2985 1504
rect 2865 1430 2985 1470
rect 2865 1396 2908 1430
rect 2942 1396 2985 1430
rect 2865 1250 2985 1396
rect 2865 1144 2872 1250
rect 2978 1144 2985 1250
rect 3295 1504 3415 2600
rect 3517 4092 3619 4118
rect 3653 4092 3755 4118
rect 3517 4082 3547 4092
rect 3725 4082 3755 4092
rect 3517 4014 3547 4048
rect 3725 4014 3755 4048
rect 3517 3946 3547 3980
rect 3725 3946 3755 3980
rect 3517 3878 3547 3912
rect 3725 3878 3755 3912
rect 3517 3810 3547 3844
rect 3725 3810 3755 3844
rect 3517 3742 3547 3776
rect 3725 3742 3755 3776
rect 3517 3674 3547 3708
rect 3725 3674 3755 3708
rect 3517 3606 3547 3640
rect 3725 3606 3755 3640
rect 3517 3538 3547 3572
rect 3725 3538 3755 3572
rect 3517 3470 3547 3504
rect 3725 3470 3755 3504
rect 3517 3402 3547 3436
rect 3725 3402 3755 3436
rect 3517 3334 3547 3368
rect 3725 3334 3755 3368
rect 3517 3266 3547 3300
rect 3725 3266 3755 3300
rect 3517 3198 3547 3232
rect 3725 3198 3755 3232
rect 3551 3164 3619 3194
rect 3653 3164 3721 3194
rect 3517 3148 3619 3164
rect 3653 3148 3755 3164
rect 3517 3108 3755 3148
rect 3517 3074 3547 3108
rect 3581 3074 3619 3108
rect 3653 3074 3691 3108
rect 3725 3074 3755 3108
rect 3517 3044 3755 3074
rect 3517 3028 3585 3044
rect 3517 2994 3547 3028
rect 3581 3010 3585 3028
rect 3619 3028 3653 3044
rect 3581 2994 3619 3010
rect 3687 3028 3755 3044
rect 3687 3010 3691 3028
rect 3653 2994 3691 3010
rect 3725 2994 3755 3028
rect 3517 2974 3755 2994
rect 3517 2948 3585 2974
rect 3517 2914 3547 2948
rect 3581 2940 3585 2948
rect 3619 2948 3653 2974
rect 3581 2914 3619 2940
rect 3687 2948 3755 2974
rect 3687 2940 3691 2948
rect 3653 2914 3691 2940
rect 3725 2914 3755 2948
rect 3517 2904 3755 2914
rect 3517 2870 3585 2904
rect 3619 2870 3653 2904
rect 3687 2870 3755 2904
rect 3517 2868 3755 2870
rect 3517 2834 3547 2868
rect 3581 2834 3619 2868
rect 3653 2834 3691 2868
rect 3725 2834 3755 2868
rect 3517 2800 3585 2834
rect 3619 2800 3653 2834
rect 3687 2800 3755 2834
rect 3517 2788 3755 2800
rect 3517 2754 3547 2788
rect 3581 2764 3619 2788
rect 3581 2754 3585 2764
rect 3517 2730 3585 2754
rect 3653 2764 3691 2788
rect 3619 2730 3653 2754
rect 3687 2754 3691 2764
rect 3725 2754 3755 2788
rect 3687 2730 3755 2754
rect 3517 2708 3755 2730
rect 3517 2674 3547 2708
rect 3581 2694 3619 2708
rect 3581 2674 3585 2694
rect 3517 2660 3585 2674
rect 3653 2694 3691 2708
rect 3619 2660 3653 2674
rect 3687 2674 3691 2694
rect 3725 2674 3755 2708
rect 3687 2660 3755 2674
rect 3517 2628 3755 2660
rect 3517 2594 3547 2628
rect 3581 2594 3619 2628
rect 3653 2594 3691 2628
rect 3725 2594 3755 2628
rect 3517 2556 3755 2594
rect 3517 2540 3619 2556
rect 3653 2540 3755 2556
rect 3551 2518 3619 2540
rect 3653 2518 3721 2540
rect 3517 2472 3547 2506
rect 3725 2472 3755 2506
rect 3517 2404 3547 2438
rect 3725 2404 3755 2438
rect 3517 2336 3547 2370
rect 3725 2336 3755 2370
rect 3517 2268 3547 2302
rect 3725 2268 3755 2302
rect 3517 2200 3547 2234
rect 3725 2200 3755 2234
rect 3517 2132 3547 2166
rect 3725 2132 3755 2166
rect 3517 2064 3547 2098
rect 3725 2064 3755 2098
rect 3517 1996 3547 2030
rect 3725 1996 3755 2030
rect 3517 1928 3547 1962
rect 3725 1928 3755 1962
rect 3517 1860 3547 1894
rect 3725 1860 3755 1894
rect 3517 1792 3547 1826
rect 3725 1792 3755 1826
rect 3517 1724 3547 1758
rect 3725 1724 3755 1758
rect 3517 1656 3547 1690
rect 3725 1656 3755 1690
rect 3517 1620 3547 1622
rect 3725 1620 3755 1622
rect 3517 1586 3619 1620
rect 3653 1586 3755 1620
rect 3517 1536 3755 1586
rect 3857 3104 3977 4200
rect 4287 4308 4407 4324
rect 4287 4274 4330 4308
rect 4364 4274 4407 4308
rect 4287 4234 4407 4274
rect 4287 4200 4330 4234
rect 4364 4200 4407 4234
rect 3857 3070 3900 3104
rect 3934 3070 3977 3104
rect 3857 3026 3977 3070
rect 3857 2992 3900 3026
rect 3934 2992 3977 3026
rect 3857 2948 3977 2992
rect 3857 2914 3900 2948
rect 3934 2914 3977 2948
rect 3857 2870 3977 2914
rect 3857 2836 3900 2870
rect 3934 2836 3977 2870
rect 3857 2792 3977 2836
rect 3857 2758 3900 2792
rect 3934 2758 3977 2792
rect 3857 2713 3977 2758
rect 3857 2679 3900 2713
rect 3934 2679 3977 2713
rect 3857 2634 3977 2679
rect 3857 2600 3900 2634
rect 3934 2600 3977 2634
rect 3295 1470 3338 1504
rect 3372 1470 3415 1504
rect 3295 1430 3415 1470
rect 3295 1396 3338 1430
rect 3372 1396 3415 1430
rect 3295 1250 3415 1396
rect 3295 1144 3302 1250
rect 3408 1144 3415 1250
rect 3857 1504 3977 2600
rect 4042 4064 4043 4098
rect 4077 4082 4115 4098
rect 4077 4064 4079 4082
rect 4042 4048 4079 4064
rect 4113 4064 4115 4082
rect 4149 4082 4187 4098
rect 4149 4064 4151 4082
rect 4113 4048 4151 4064
rect 4185 4064 4187 4082
rect 4221 4064 4222 4098
rect 4185 4048 4222 4064
rect 4042 4025 4222 4048
rect 4042 3991 4043 4025
rect 4077 4014 4115 4025
rect 4077 3991 4079 4014
rect 4042 3980 4079 3991
rect 4113 3991 4115 4014
rect 4149 4014 4187 4025
rect 4149 3991 4151 4014
rect 4113 3980 4151 3991
rect 4185 3991 4187 4014
rect 4221 3991 4222 4025
rect 4185 3980 4222 3991
rect 4042 3952 4222 3980
rect 4042 3918 4043 3952
rect 4077 3946 4115 3952
rect 4077 3918 4079 3946
rect 4042 3912 4079 3918
rect 4113 3918 4115 3946
rect 4149 3946 4187 3952
rect 4149 3918 4151 3946
rect 4113 3912 4151 3918
rect 4185 3918 4187 3946
rect 4221 3918 4222 3952
rect 4185 3912 4222 3918
rect 4042 3879 4222 3912
rect 4042 3845 4043 3879
rect 4077 3878 4115 3879
rect 4077 3845 4079 3878
rect 4042 3844 4079 3845
rect 4113 3845 4115 3878
rect 4149 3878 4187 3879
rect 4149 3845 4151 3878
rect 4113 3844 4151 3845
rect 4185 3845 4187 3878
rect 4221 3845 4222 3879
rect 4185 3844 4222 3845
rect 4042 3810 4222 3844
rect 4042 3806 4079 3810
rect 4042 3772 4043 3806
rect 4077 3776 4079 3806
rect 4113 3806 4151 3810
rect 4113 3776 4115 3806
rect 4077 3772 4115 3776
rect 4149 3776 4151 3806
rect 4185 3806 4222 3810
rect 4185 3776 4187 3806
rect 4149 3772 4187 3776
rect 4221 3772 4222 3806
rect 4042 3742 4222 3772
rect 4042 3733 4079 3742
rect 4042 3699 4043 3733
rect 4077 3708 4079 3733
rect 4113 3733 4151 3742
rect 4113 3708 4115 3733
rect 4077 3699 4115 3708
rect 4149 3708 4151 3733
rect 4185 3733 4222 3742
rect 4185 3708 4187 3733
rect 4149 3699 4187 3708
rect 4221 3699 4222 3733
rect 4042 3674 4222 3699
rect 4042 3660 4079 3674
rect 4042 3626 4043 3660
rect 4077 3640 4079 3660
rect 4113 3660 4151 3674
rect 4113 3640 4115 3660
rect 4077 3626 4115 3640
rect 4149 3640 4151 3660
rect 4185 3660 4222 3674
rect 4185 3640 4187 3660
rect 4149 3626 4187 3640
rect 4221 3626 4222 3660
rect 4042 3606 4222 3626
rect 4042 3587 4079 3606
rect 4042 3553 4043 3587
rect 4077 3572 4079 3587
rect 4113 3587 4151 3606
rect 4113 3572 4115 3587
rect 4077 3553 4115 3572
rect 4149 3572 4151 3587
rect 4185 3587 4222 3606
rect 4185 3572 4187 3587
rect 4149 3553 4187 3572
rect 4221 3553 4222 3587
rect 4042 3538 4222 3553
rect 4042 3514 4079 3538
rect 4042 3480 4043 3514
rect 4077 3504 4079 3514
rect 4113 3514 4151 3538
rect 4113 3504 4115 3514
rect 4077 3480 4115 3504
rect 4149 3504 4151 3514
rect 4185 3514 4222 3538
rect 4185 3504 4187 3514
rect 4149 3480 4187 3504
rect 4221 3480 4222 3514
rect 4042 3470 4222 3480
rect 4042 3441 4079 3470
rect 4042 3407 4043 3441
rect 4077 3436 4079 3441
rect 4113 3441 4151 3470
rect 4113 3436 4115 3441
rect 4077 3407 4115 3436
rect 4149 3436 4151 3441
rect 4185 3441 4222 3470
rect 4185 3436 4187 3441
rect 4149 3407 4187 3436
rect 4221 3407 4222 3441
rect 4042 3402 4222 3407
rect 4042 3368 4079 3402
rect 4113 3368 4151 3402
rect 4185 3368 4222 3402
rect 4042 3334 4043 3368
rect 4077 3334 4115 3368
rect 4149 3334 4187 3368
rect 4221 3334 4222 3368
rect 4042 3300 4079 3334
rect 4113 3300 4151 3334
rect 4185 3300 4222 3334
rect 4042 3295 4222 3300
rect 4042 3261 4043 3295
rect 4077 3266 4115 3295
rect 4077 3261 4079 3266
rect 4042 3232 4079 3261
rect 4113 3261 4115 3266
rect 4149 3266 4187 3295
rect 4149 3261 4151 3266
rect 4113 3232 4151 3261
rect 4185 3261 4187 3266
rect 4221 3261 4222 3295
rect 4185 3232 4222 3261
rect 4042 3222 4222 3232
rect 4042 3188 4043 3222
rect 4077 3198 4115 3222
rect 4077 3188 4079 3198
rect 4042 3164 4079 3188
rect 4113 3188 4115 3198
rect 4149 3198 4187 3222
rect 4149 3188 4151 3198
rect 4113 3164 4151 3188
rect 4185 3188 4187 3198
rect 4221 3188 4222 3222
rect 4185 3164 4222 3188
rect 4042 3149 4222 3164
rect 4042 3115 4043 3149
rect 4077 3115 4115 3149
rect 4149 3115 4187 3149
rect 4221 3115 4222 3149
rect 4042 3076 4222 3115
rect 4042 3042 4043 3076
rect 4077 3042 4115 3076
rect 4149 3042 4187 3076
rect 4221 3042 4222 3076
rect 4042 3003 4222 3042
rect 4042 2969 4043 3003
rect 4077 2969 4115 3003
rect 4149 2969 4187 3003
rect 4221 2969 4222 3003
rect 4042 2930 4222 2969
rect 4042 2896 4043 2930
rect 4077 2896 4115 2930
rect 4149 2896 4187 2930
rect 4221 2896 4222 2930
rect 4042 2857 4222 2896
rect 4042 2823 4043 2857
rect 4077 2823 4115 2857
rect 4149 2823 4187 2857
rect 4221 2823 4222 2857
rect 4042 2784 4222 2823
rect 4042 2750 4043 2784
rect 4077 2750 4115 2784
rect 4149 2750 4187 2784
rect 4221 2750 4222 2784
rect 4042 2711 4222 2750
rect 4042 2677 4043 2711
rect 4077 2677 4115 2711
rect 4149 2677 4187 2711
rect 4221 2677 4222 2711
rect 4042 2638 4222 2677
rect 4042 2604 4043 2638
rect 4077 2604 4115 2638
rect 4149 2604 4187 2638
rect 4221 2604 4222 2638
rect 4042 2565 4222 2604
rect 4042 2531 4043 2565
rect 4077 2531 4115 2565
rect 4149 2531 4187 2565
rect 4221 2531 4222 2565
rect 4042 2492 4222 2531
rect 4042 2458 4043 2492
rect 4077 2482 4115 2492
rect 4077 2458 4079 2482
rect 4042 2448 4079 2458
rect 4113 2458 4115 2482
rect 4149 2482 4187 2492
rect 4149 2458 4151 2482
rect 4113 2448 4151 2458
rect 4185 2458 4187 2482
rect 4221 2458 4222 2492
rect 4185 2448 4222 2458
rect 4042 2419 4222 2448
rect 4042 2385 4043 2419
rect 4077 2414 4115 2419
rect 4077 2385 4079 2414
rect 4042 2380 4079 2385
rect 4113 2385 4115 2414
rect 4149 2414 4187 2419
rect 4149 2385 4151 2414
rect 4113 2380 4151 2385
rect 4185 2385 4187 2414
rect 4221 2385 4222 2419
rect 4185 2380 4222 2385
rect 4042 2346 4222 2380
rect 4042 2312 4043 2346
rect 4077 2312 4079 2346
rect 4113 2312 4115 2346
rect 4149 2312 4151 2346
rect 4185 2312 4187 2346
rect 4221 2312 4222 2346
rect 4042 2278 4222 2312
rect 4042 2273 4079 2278
rect 4042 2239 4043 2273
rect 4077 2244 4079 2273
rect 4113 2273 4151 2278
rect 4113 2244 4115 2273
rect 4077 2239 4115 2244
rect 4149 2244 4151 2273
rect 4185 2273 4222 2278
rect 4185 2244 4187 2273
rect 4149 2239 4187 2244
rect 4221 2239 4222 2273
rect 4042 2210 4222 2239
rect 4042 2200 4079 2210
rect 4042 2166 4043 2200
rect 4077 2176 4079 2200
rect 4113 2200 4151 2210
rect 4113 2176 4115 2200
rect 4077 2166 4115 2176
rect 4149 2176 4151 2200
rect 4185 2200 4222 2210
rect 4185 2176 4187 2200
rect 4149 2166 4187 2176
rect 4221 2166 4222 2200
rect 4042 2142 4222 2166
rect 4042 2126 4079 2142
rect 4042 2092 4043 2126
rect 4077 2108 4079 2126
rect 4113 2126 4151 2142
rect 4113 2108 4115 2126
rect 4077 2092 4115 2108
rect 4149 2108 4151 2126
rect 4185 2126 4222 2142
rect 4185 2108 4187 2126
rect 4149 2092 4187 2108
rect 4221 2092 4222 2126
rect 4042 2074 4222 2092
rect 4042 2052 4079 2074
rect 4042 2018 4043 2052
rect 4077 2040 4079 2052
rect 4113 2052 4151 2074
rect 4113 2040 4115 2052
rect 4077 2018 4115 2040
rect 4149 2040 4151 2052
rect 4185 2052 4222 2074
rect 4185 2040 4187 2052
rect 4149 2018 4187 2040
rect 4221 2018 4222 2052
rect 4042 2006 4222 2018
rect 4042 1978 4079 2006
rect 4042 1944 4043 1978
rect 4077 1972 4079 1978
rect 4113 1978 4151 2006
rect 4113 1972 4115 1978
rect 4077 1944 4115 1972
rect 4149 1972 4151 1978
rect 4185 1978 4222 2006
rect 4185 1972 4187 1978
rect 4149 1944 4187 1972
rect 4221 1944 4222 1978
rect 4042 1938 4222 1944
rect 4042 1904 4079 1938
rect 4113 1904 4151 1938
rect 4185 1904 4222 1938
rect 4042 1870 4043 1904
rect 4077 1870 4115 1904
rect 4149 1870 4187 1904
rect 4221 1870 4222 1904
rect 4042 1836 4079 1870
rect 4113 1836 4151 1870
rect 4185 1836 4222 1870
rect 4042 1830 4222 1836
rect 4042 1796 4043 1830
rect 4077 1802 4115 1830
rect 4077 1796 4079 1802
rect 4042 1768 4079 1796
rect 4113 1796 4115 1802
rect 4149 1802 4187 1830
rect 4149 1796 4151 1802
rect 4113 1768 4151 1796
rect 4185 1796 4187 1802
rect 4221 1796 4222 1830
rect 4185 1768 4222 1796
rect 4042 1756 4222 1768
rect 4042 1722 4043 1756
rect 4077 1734 4115 1756
rect 4077 1722 4079 1734
rect 4042 1700 4079 1722
rect 4113 1722 4115 1734
rect 4149 1734 4187 1756
rect 4149 1722 4151 1734
rect 4113 1700 4151 1722
rect 4185 1722 4187 1734
rect 4221 1722 4222 1756
rect 4185 1700 4222 1722
rect 4042 1682 4222 1700
rect 4042 1648 4043 1682
rect 4077 1666 4115 1682
rect 4077 1648 4079 1666
rect 4042 1632 4079 1648
rect 4113 1648 4115 1666
rect 4149 1666 4187 1682
rect 4149 1648 4151 1666
rect 4113 1632 4151 1648
rect 4185 1648 4187 1666
rect 4221 1648 4222 1682
rect 4185 1632 4222 1648
rect 4042 1608 4222 1632
rect 4042 1574 4043 1608
rect 4077 1598 4115 1608
rect 4077 1574 4079 1598
rect 4042 1564 4079 1574
rect 4113 1574 4115 1598
rect 4149 1598 4187 1608
rect 4149 1574 4151 1598
rect 4113 1564 4151 1574
rect 4185 1574 4187 1598
rect 4221 1574 4222 1608
rect 4185 1564 4222 1574
rect 4042 1548 4222 1564
rect 4287 3104 4407 4200
rect 4849 4308 4969 4324
rect 4849 4274 4892 4308
rect 4926 4274 4969 4308
rect 4849 4234 4969 4274
rect 4849 4200 4892 4234
rect 4926 4200 4969 4234
rect 4287 3070 4330 3104
rect 4364 3070 4407 3104
rect 4287 3026 4407 3070
rect 4287 2992 4330 3026
rect 4364 2992 4407 3026
rect 4287 2948 4407 2992
rect 4287 2914 4330 2948
rect 4364 2914 4407 2948
rect 4287 2870 4407 2914
rect 4287 2836 4330 2870
rect 4364 2836 4407 2870
rect 4287 2792 4407 2836
rect 4287 2758 4330 2792
rect 4364 2758 4407 2792
rect 4287 2713 4407 2758
rect 4287 2679 4330 2713
rect 4364 2679 4407 2713
rect 4287 2634 4407 2679
rect 4287 2600 4330 2634
rect 4364 2600 4407 2634
rect 3857 1470 3900 1504
rect 3934 1470 3977 1504
rect 3857 1430 3977 1470
rect 3857 1396 3900 1430
rect 3934 1396 3977 1430
rect 3857 1250 3977 1396
rect 3857 1144 3864 1250
rect 3970 1144 3977 1250
rect 4287 1504 4407 2600
rect 4509 4092 4611 4118
rect 4645 4092 4747 4118
rect 4509 4082 4539 4092
rect 4717 4082 4747 4092
rect 4509 4014 4539 4048
rect 4717 4014 4747 4048
rect 4509 3946 4539 3980
rect 4717 3946 4747 3980
rect 4509 3878 4539 3912
rect 4717 3878 4747 3912
rect 4509 3810 4539 3844
rect 4717 3810 4747 3844
rect 4509 3742 4539 3776
rect 4717 3742 4747 3776
rect 4509 3674 4539 3708
rect 4717 3674 4747 3708
rect 4509 3606 4539 3640
rect 4717 3606 4747 3640
rect 4509 3538 4539 3572
rect 4717 3538 4747 3572
rect 4509 3470 4539 3504
rect 4717 3470 4747 3504
rect 4509 3402 4539 3436
rect 4717 3402 4747 3436
rect 4509 3334 4539 3368
rect 4717 3334 4747 3368
rect 4509 3266 4539 3300
rect 4717 3266 4747 3300
rect 4509 3198 4539 3232
rect 4717 3198 4747 3232
rect 4543 3164 4611 3194
rect 4645 3164 4713 3194
rect 4509 3148 4611 3164
rect 4645 3148 4747 3164
rect 4509 3108 4747 3148
rect 4509 3074 4539 3108
rect 4573 3074 4611 3108
rect 4645 3074 4683 3108
rect 4717 3074 4747 3108
rect 4509 3044 4747 3074
rect 4509 3028 4577 3044
rect 4509 2994 4539 3028
rect 4573 3010 4577 3028
rect 4611 3028 4645 3044
rect 4573 2994 4611 3010
rect 4679 3028 4747 3044
rect 4679 3010 4683 3028
rect 4645 2994 4683 3010
rect 4717 2994 4747 3028
rect 4509 2974 4747 2994
rect 4509 2948 4577 2974
rect 4509 2914 4539 2948
rect 4573 2940 4577 2948
rect 4611 2948 4645 2974
rect 4573 2914 4611 2940
rect 4679 2948 4747 2974
rect 4679 2940 4683 2948
rect 4645 2914 4683 2940
rect 4717 2914 4747 2948
rect 4509 2904 4747 2914
rect 4509 2870 4577 2904
rect 4611 2870 4645 2904
rect 4679 2870 4747 2904
rect 4509 2868 4747 2870
rect 4509 2834 4539 2868
rect 4573 2834 4611 2868
rect 4645 2834 4683 2868
rect 4717 2834 4747 2868
rect 4509 2800 4577 2834
rect 4611 2800 4645 2834
rect 4679 2800 4747 2834
rect 4509 2788 4747 2800
rect 4509 2754 4539 2788
rect 4573 2764 4611 2788
rect 4573 2754 4577 2764
rect 4509 2730 4577 2754
rect 4645 2764 4683 2788
rect 4611 2730 4645 2754
rect 4679 2754 4683 2764
rect 4717 2754 4747 2788
rect 4679 2730 4747 2754
rect 4509 2708 4747 2730
rect 4509 2674 4539 2708
rect 4573 2694 4611 2708
rect 4573 2674 4577 2694
rect 4509 2660 4577 2674
rect 4645 2694 4683 2708
rect 4611 2660 4645 2674
rect 4679 2674 4683 2694
rect 4717 2674 4747 2708
rect 4679 2660 4747 2674
rect 4509 2628 4747 2660
rect 4509 2594 4539 2628
rect 4573 2594 4611 2628
rect 4645 2594 4683 2628
rect 4717 2594 4747 2628
rect 4509 2556 4747 2594
rect 4509 2540 4611 2556
rect 4645 2540 4747 2556
rect 4543 2518 4611 2540
rect 4645 2518 4713 2540
rect 4509 2472 4539 2506
rect 4717 2472 4747 2506
rect 4509 2404 4539 2438
rect 4717 2404 4747 2438
rect 4509 2336 4539 2370
rect 4717 2336 4747 2370
rect 4509 2268 4539 2302
rect 4717 2268 4747 2302
rect 4509 2200 4539 2234
rect 4717 2200 4747 2234
rect 4509 2132 4539 2166
rect 4717 2132 4747 2166
rect 4509 2064 4539 2098
rect 4717 2064 4747 2098
rect 4509 1996 4539 2030
rect 4717 1996 4747 2030
rect 4509 1928 4539 1962
rect 4717 1928 4747 1962
rect 4509 1860 4539 1894
rect 4717 1860 4747 1894
rect 4509 1792 4539 1826
rect 4717 1792 4747 1826
rect 4509 1724 4539 1758
rect 4717 1724 4747 1758
rect 4509 1656 4539 1690
rect 4717 1656 4747 1690
rect 4509 1620 4539 1622
rect 4717 1620 4747 1622
rect 4509 1586 4611 1620
rect 4645 1586 4747 1620
rect 4509 1536 4747 1586
rect 4849 3104 4969 4200
rect 5279 4308 5399 4324
rect 5279 4274 5322 4308
rect 5356 4274 5399 4308
rect 5279 4234 5399 4274
rect 5279 4200 5322 4234
rect 5356 4200 5399 4234
rect 4849 3070 4892 3104
rect 4926 3070 4969 3104
rect 4849 3026 4969 3070
rect 4849 2992 4892 3026
rect 4926 2992 4969 3026
rect 4849 2948 4969 2992
rect 4849 2914 4892 2948
rect 4926 2914 4969 2948
rect 4849 2870 4969 2914
rect 4849 2836 4892 2870
rect 4926 2836 4969 2870
rect 4849 2792 4969 2836
rect 4849 2758 4892 2792
rect 4926 2758 4969 2792
rect 4849 2713 4969 2758
rect 4849 2679 4892 2713
rect 4926 2679 4969 2713
rect 4849 2634 4969 2679
rect 4849 2600 4892 2634
rect 4926 2600 4969 2634
rect 4287 1470 4330 1504
rect 4364 1470 4407 1504
rect 4287 1430 4407 1470
rect 4287 1396 4330 1430
rect 4364 1396 4407 1430
rect 4287 1250 4407 1396
rect 4287 1144 4294 1250
rect 4400 1144 4407 1250
rect 4849 1504 4969 2600
rect 5034 4064 5035 4098
rect 5069 4082 5107 4098
rect 5069 4064 5071 4082
rect 5034 4048 5071 4064
rect 5105 4064 5107 4082
rect 5141 4082 5179 4098
rect 5141 4064 5143 4082
rect 5105 4048 5143 4064
rect 5177 4064 5179 4082
rect 5213 4064 5214 4098
rect 5177 4048 5214 4064
rect 5034 4025 5214 4048
rect 5034 3991 5035 4025
rect 5069 4014 5107 4025
rect 5069 3991 5071 4014
rect 5034 3980 5071 3991
rect 5105 3991 5107 4014
rect 5141 4014 5179 4025
rect 5141 3991 5143 4014
rect 5105 3980 5143 3991
rect 5177 3991 5179 4014
rect 5213 3991 5214 4025
rect 5177 3980 5214 3991
rect 5034 3952 5214 3980
rect 5034 3918 5035 3952
rect 5069 3946 5107 3952
rect 5069 3918 5071 3946
rect 5034 3912 5071 3918
rect 5105 3918 5107 3946
rect 5141 3946 5179 3952
rect 5141 3918 5143 3946
rect 5105 3912 5143 3918
rect 5177 3918 5179 3946
rect 5213 3918 5214 3952
rect 5177 3912 5214 3918
rect 5034 3879 5214 3912
rect 5034 3845 5035 3879
rect 5069 3878 5107 3879
rect 5069 3845 5071 3878
rect 5034 3844 5071 3845
rect 5105 3845 5107 3878
rect 5141 3878 5179 3879
rect 5141 3845 5143 3878
rect 5105 3844 5143 3845
rect 5177 3845 5179 3878
rect 5213 3845 5214 3879
rect 5177 3844 5214 3845
rect 5034 3810 5214 3844
rect 5034 3806 5071 3810
rect 5034 3772 5035 3806
rect 5069 3776 5071 3806
rect 5105 3806 5143 3810
rect 5105 3776 5107 3806
rect 5069 3772 5107 3776
rect 5141 3776 5143 3806
rect 5177 3806 5214 3810
rect 5177 3776 5179 3806
rect 5141 3772 5179 3776
rect 5213 3772 5214 3806
rect 5034 3742 5214 3772
rect 5034 3733 5071 3742
rect 5034 3699 5035 3733
rect 5069 3708 5071 3733
rect 5105 3733 5143 3742
rect 5105 3708 5107 3733
rect 5069 3699 5107 3708
rect 5141 3708 5143 3733
rect 5177 3733 5214 3742
rect 5177 3708 5179 3733
rect 5141 3699 5179 3708
rect 5213 3699 5214 3733
rect 5034 3674 5214 3699
rect 5034 3660 5071 3674
rect 5034 3626 5035 3660
rect 5069 3640 5071 3660
rect 5105 3660 5143 3674
rect 5105 3640 5107 3660
rect 5069 3626 5107 3640
rect 5141 3640 5143 3660
rect 5177 3660 5214 3674
rect 5177 3640 5179 3660
rect 5141 3626 5179 3640
rect 5213 3626 5214 3660
rect 5034 3606 5214 3626
rect 5034 3587 5071 3606
rect 5034 3553 5035 3587
rect 5069 3572 5071 3587
rect 5105 3587 5143 3606
rect 5105 3572 5107 3587
rect 5069 3553 5107 3572
rect 5141 3572 5143 3587
rect 5177 3587 5214 3606
rect 5177 3572 5179 3587
rect 5141 3553 5179 3572
rect 5213 3553 5214 3587
rect 5034 3538 5214 3553
rect 5034 3514 5071 3538
rect 5034 3480 5035 3514
rect 5069 3504 5071 3514
rect 5105 3514 5143 3538
rect 5105 3504 5107 3514
rect 5069 3480 5107 3504
rect 5141 3504 5143 3514
rect 5177 3514 5214 3538
rect 5177 3504 5179 3514
rect 5141 3480 5179 3504
rect 5213 3480 5214 3514
rect 5034 3470 5214 3480
rect 5034 3441 5071 3470
rect 5034 3407 5035 3441
rect 5069 3436 5071 3441
rect 5105 3441 5143 3470
rect 5105 3436 5107 3441
rect 5069 3407 5107 3436
rect 5141 3436 5143 3441
rect 5177 3441 5214 3470
rect 5177 3436 5179 3441
rect 5141 3407 5179 3436
rect 5213 3407 5214 3441
rect 5034 3402 5214 3407
rect 5034 3368 5071 3402
rect 5105 3368 5143 3402
rect 5177 3368 5214 3402
rect 5034 3334 5035 3368
rect 5069 3334 5107 3368
rect 5141 3334 5179 3368
rect 5213 3334 5214 3368
rect 5034 3300 5071 3334
rect 5105 3300 5143 3334
rect 5177 3300 5214 3334
rect 5034 3295 5214 3300
rect 5034 3261 5035 3295
rect 5069 3266 5107 3295
rect 5069 3261 5071 3266
rect 5034 3232 5071 3261
rect 5105 3261 5107 3266
rect 5141 3266 5179 3295
rect 5141 3261 5143 3266
rect 5105 3232 5143 3261
rect 5177 3261 5179 3266
rect 5213 3261 5214 3295
rect 5177 3232 5214 3261
rect 5034 3222 5214 3232
rect 5034 3188 5035 3222
rect 5069 3198 5107 3222
rect 5069 3188 5071 3198
rect 5034 3164 5071 3188
rect 5105 3188 5107 3198
rect 5141 3198 5179 3222
rect 5141 3188 5143 3198
rect 5105 3164 5143 3188
rect 5177 3188 5179 3198
rect 5213 3188 5214 3222
rect 5177 3164 5214 3188
rect 5034 3149 5214 3164
rect 5034 3115 5035 3149
rect 5069 3115 5107 3149
rect 5141 3115 5179 3149
rect 5213 3115 5214 3149
rect 5034 3076 5214 3115
rect 5034 3042 5035 3076
rect 5069 3042 5107 3076
rect 5141 3042 5179 3076
rect 5213 3042 5214 3076
rect 5034 3003 5214 3042
rect 5034 2969 5035 3003
rect 5069 2969 5107 3003
rect 5141 2969 5179 3003
rect 5213 2969 5214 3003
rect 5034 2930 5214 2969
rect 5034 2896 5035 2930
rect 5069 2896 5107 2930
rect 5141 2896 5179 2930
rect 5213 2896 5214 2930
rect 5034 2857 5214 2896
rect 5034 2823 5035 2857
rect 5069 2823 5107 2857
rect 5141 2823 5179 2857
rect 5213 2823 5214 2857
rect 5034 2784 5214 2823
rect 5034 2750 5035 2784
rect 5069 2750 5107 2784
rect 5141 2750 5179 2784
rect 5213 2750 5214 2784
rect 5034 2711 5214 2750
rect 5034 2677 5035 2711
rect 5069 2677 5107 2711
rect 5141 2677 5179 2711
rect 5213 2677 5214 2711
rect 5034 2638 5214 2677
rect 5034 2604 5035 2638
rect 5069 2604 5107 2638
rect 5141 2604 5179 2638
rect 5213 2604 5214 2638
rect 5034 2565 5214 2604
rect 5034 2531 5035 2565
rect 5069 2531 5107 2565
rect 5141 2531 5179 2565
rect 5213 2531 5214 2565
rect 5034 2492 5214 2531
rect 5034 2458 5035 2492
rect 5069 2482 5107 2492
rect 5069 2458 5071 2482
rect 5034 2448 5071 2458
rect 5105 2458 5107 2482
rect 5141 2482 5179 2492
rect 5141 2458 5143 2482
rect 5105 2448 5143 2458
rect 5177 2458 5179 2482
rect 5213 2458 5214 2492
rect 5177 2448 5214 2458
rect 5034 2419 5214 2448
rect 5034 2385 5035 2419
rect 5069 2414 5107 2419
rect 5069 2385 5071 2414
rect 5034 2380 5071 2385
rect 5105 2385 5107 2414
rect 5141 2414 5179 2419
rect 5141 2385 5143 2414
rect 5105 2380 5143 2385
rect 5177 2385 5179 2414
rect 5213 2385 5214 2419
rect 5177 2380 5214 2385
rect 5034 2346 5214 2380
rect 5034 2312 5035 2346
rect 5069 2312 5071 2346
rect 5105 2312 5107 2346
rect 5141 2312 5143 2346
rect 5177 2312 5179 2346
rect 5213 2312 5214 2346
rect 5034 2278 5214 2312
rect 5034 2273 5071 2278
rect 5034 2239 5035 2273
rect 5069 2244 5071 2273
rect 5105 2273 5143 2278
rect 5105 2244 5107 2273
rect 5069 2239 5107 2244
rect 5141 2244 5143 2273
rect 5177 2273 5214 2278
rect 5177 2244 5179 2273
rect 5141 2239 5179 2244
rect 5213 2239 5214 2273
rect 5034 2210 5214 2239
rect 5034 2200 5071 2210
rect 5034 2166 5035 2200
rect 5069 2176 5071 2200
rect 5105 2200 5143 2210
rect 5105 2176 5107 2200
rect 5069 2166 5107 2176
rect 5141 2176 5143 2200
rect 5177 2200 5214 2210
rect 5177 2176 5179 2200
rect 5141 2166 5179 2176
rect 5213 2166 5214 2200
rect 5034 2142 5214 2166
rect 5034 2126 5071 2142
rect 5034 2092 5035 2126
rect 5069 2108 5071 2126
rect 5105 2126 5143 2142
rect 5105 2108 5107 2126
rect 5069 2092 5107 2108
rect 5141 2108 5143 2126
rect 5177 2126 5214 2142
rect 5177 2108 5179 2126
rect 5141 2092 5179 2108
rect 5213 2092 5214 2126
rect 5034 2074 5214 2092
rect 5034 2052 5071 2074
rect 5034 2018 5035 2052
rect 5069 2040 5071 2052
rect 5105 2052 5143 2074
rect 5105 2040 5107 2052
rect 5069 2018 5107 2040
rect 5141 2040 5143 2052
rect 5177 2052 5214 2074
rect 5177 2040 5179 2052
rect 5141 2018 5179 2040
rect 5213 2018 5214 2052
rect 5034 2006 5214 2018
rect 5034 1978 5071 2006
rect 5034 1944 5035 1978
rect 5069 1972 5071 1978
rect 5105 1978 5143 2006
rect 5105 1972 5107 1978
rect 5069 1944 5107 1972
rect 5141 1972 5143 1978
rect 5177 1978 5214 2006
rect 5177 1972 5179 1978
rect 5141 1944 5179 1972
rect 5213 1944 5214 1978
rect 5034 1938 5214 1944
rect 5034 1904 5071 1938
rect 5105 1904 5143 1938
rect 5177 1904 5214 1938
rect 5034 1870 5035 1904
rect 5069 1870 5107 1904
rect 5141 1870 5179 1904
rect 5213 1870 5214 1904
rect 5034 1836 5071 1870
rect 5105 1836 5143 1870
rect 5177 1836 5214 1870
rect 5034 1830 5214 1836
rect 5034 1796 5035 1830
rect 5069 1802 5107 1830
rect 5069 1796 5071 1802
rect 5034 1768 5071 1796
rect 5105 1796 5107 1802
rect 5141 1802 5179 1830
rect 5141 1796 5143 1802
rect 5105 1768 5143 1796
rect 5177 1796 5179 1802
rect 5213 1796 5214 1830
rect 5177 1768 5214 1796
rect 5034 1756 5214 1768
rect 5034 1722 5035 1756
rect 5069 1734 5107 1756
rect 5069 1722 5071 1734
rect 5034 1700 5071 1722
rect 5105 1722 5107 1734
rect 5141 1734 5179 1756
rect 5141 1722 5143 1734
rect 5105 1700 5143 1722
rect 5177 1722 5179 1734
rect 5213 1722 5214 1756
rect 5177 1700 5214 1722
rect 5034 1682 5214 1700
rect 5034 1648 5035 1682
rect 5069 1666 5107 1682
rect 5069 1648 5071 1666
rect 5034 1632 5071 1648
rect 5105 1648 5107 1666
rect 5141 1666 5179 1682
rect 5141 1648 5143 1666
rect 5105 1632 5143 1648
rect 5177 1648 5179 1666
rect 5213 1648 5214 1682
rect 5177 1632 5214 1648
rect 5034 1608 5214 1632
rect 5034 1574 5035 1608
rect 5069 1598 5107 1608
rect 5069 1574 5071 1598
rect 5034 1564 5071 1574
rect 5105 1574 5107 1598
rect 5141 1598 5179 1608
rect 5141 1574 5143 1598
rect 5105 1564 5143 1574
rect 5177 1574 5179 1598
rect 5213 1574 5214 1608
rect 5177 1564 5214 1574
rect 5034 1548 5214 1564
rect 5279 3104 5399 4200
rect 5841 4308 5961 4324
rect 5841 4274 5884 4308
rect 5918 4274 5961 4308
rect 5841 4234 5961 4274
rect 5841 4200 5884 4234
rect 5918 4200 5961 4234
rect 5279 3070 5322 3104
rect 5356 3070 5399 3104
rect 5279 3026 5399 3070
rect 5279 2992 5322 3026
rect 5356 2992 5399 3026
rect 5279 2948 5399 2992
rect 5279 2914 5322 2948
rect 5356 2914 5399 2948
rect 5279 2870 5399 2914
rect 5279 2836 5322 2870
rect 5356 2836 5399 2870
rect 5279 2792 5399 2836
rect 5279 2758 5322 2792
rect 5356 2758 5399 2792
rect 5279 2713 5399 2758
rect 5279 2679 5322 2713
rect 5356 2679 5399 2713
rect 5279 2634 5399 2679
rect 5279 2600 5322 2634
rect 5356 2600 5399 2634
rect 4849 1470 4892 1504
rect 4926 1470 4969 1504
rect 4849 1430 4969 1470
rect 4849 1396 4892 1430
rect 4926 1396 4969 1430
rect 4849 1250 4969 1396
rect 4849 1144 4856 1250
rect 4962 1144 4969 1250
rect 5279 1504 5399 2600
rect 5501 4092 5603 4118
rect 5637 4092 5739 4118
rect 5501 4082 5531 4092
rect 5709 4082 5739 4092
rect 5501 4014 5531 4048
rect 5709 4014 5739 4048
rect 5501 3946 5531 3980
rect 5709 3946 5739 3980
rect 5501 3878 5531 3912
rect 5709 3878 5739 3912
rect 5501 3810 5531 3844
rect 5709 3810 5739 3844
rect 5501 3742 5531 3776
rect 5709 3742 5739 3776
rect 5501 3674 5531 3708
rect 5709 3674 5739 3708
rect 5501 3606 5531 3640
rect 5709 3606 5739 3640
rect 5501 3538 5531 3572
rect 5709 3538 5739 3572
rect 5501 3470 5531 3504
rect 5709 3470 5739 3504
rect 5501 3402 5531 3436
rect 5709 3402 5739 3436
rect 5501 3334 5531 3368
rect 5709 3334 5739 3368
rect 5501 3266 5531 3300
rect 5709 3266 5739 3300
rect 5501 3198 5531 3232
rect 5709 3198 5739 3232
rect 5535 3164 5603 3194
rect 5637 3164 5705 3194
rect 5501 3148 5603 3164
rect 5637 3148 5739 3164
rect 5501 3108 5739 3148
rect 5501 3074 5531 3108
rect 5565 3074 5603 3108
rect 5637 3074 5675 3108
rect 5709 3074 5739 3108
rect 5501 3044 5739 3074
rect 5501 3028 5569 3044
rect 5501 2994 5531 3028
rect 5565 3010 5569 3028
rect 5603 3028 5637 3044
rect 5565 2994 5603 3010
rect 5671 3028 5739 3044
rect 5671 3010 5675 3028
rect 5637 2994 5675 3010
rect 5709 2994 5739 3028
rect 5501 2974 5739 2994
rect 5501 2948 5569 2974
rect 5501 2914 5531 2948
rect 5565 2940 5569 2948
rect 5603 2948 5637 2974
rect 5565 2914 5603 2940
rect 5671 2948 5739 2974
rect 5671 2940 5675 2948
rect 5637 2914 5675 2940
rect 5709 2914 5739 2948
rect 5501 2904 5739 2914
rect 5501 2870 5569 2904
rect 5603 2870 5637 2904
rect 5671 2870 5739 2904
rect 5501 2868 5739 2870
rect 5501 2834 5531 2868
rect 5565 2834 5603 2868
rect 5637 2834 5675 2868
rect 5709 2834 5739 2868
rect 5501 2800 5569 2834
rect 5603 2800 5637 2834
rect 5671 2800 5739 2834
rect 5501 2788 5739 2800
rect 5501 2754 5531 2788
rect 5565 2764 5603 2788
rect 5565 2754 5569 2764
rect 5501 2730 5569 2754
rect 5637 2764 5675 2788
rect 5603 2730 5637 2754
rect 5671 2754 5675 2764
rect 5709 2754 5739 2788
rect 5671 2730 5739 2754
rect 5501 2708 5739 2730
rect 5501 2674 5531 2708
rect 5565 2694 5603 2708
rect 5565 2674 5569 2694
rect 5501 2660 5569 2674
rect 5637 2694 5675 2708
rect 5603 2660 5637 2674
rect 5671 2674 5675 2694
rect 5709 2674 5739 2708
rect 5671 2660 5739 2674
rect 5501 2628 5739 2660
rect 5501 2594 5531 2628
rect 5565 2594 5603 2628
rect 5637 2594 5675 2628
rect 5709 2594 5739 2628
rect 5501 2556 5739 2594
rect 5501 2540 5603 2556
rect 5637 2540 5739 2556
rect 5535 2518 5603 2540
rect 5637 2518 5705 2540
rect 5501 2472 5531 2506
rect 5709 2472 5739 2506
rect 5501 2404 5531 2438
rect 5709 2404 5739 2438
rect 5501 2336 5531 2370
rect 5709 2336 5739 2370
rect 5501 2268 5531 2302
rect 5709 2268 5739 2302
rect 5501 2200 5531 2234
rect 5709 2200 5739 2234
rect 5501 2132 5531 2166
rect 5709 2132 5739 2166
rect 5501 2064 5531 2098
rect 5709 2064 5739 2098
rect 5501 1996 5531 2030
rect 5709 1996 5739 2030
rect 5501 1928 5531 1962
rect 5709 1928 5739 1962
rect 5501 1860 5531 1894
rect 5709 1860 5739 1894
rect 5501 1792 5531 1826
rect 5709 1792 5739 1826
rect 5501 1724 5531 1758
rect 5709 1724 5739 1758
rect 5501 1656 5531 1690
rect 5709 1656 5739 1690
rect 5501 1620 5531 1622
rect 5709 1620 5739 1622
rect 5501 1586 5603 1620
rect 5637 1586 5739 1620
rect 5501 1536 5739 1586
rect 5841 3104 5961 4200
rect 6271 4308 6391 4324
rect 6271 4274 6314 4308
rect 6348 4274 6391 4308
rect 6271 4234 6391 4274
rect 6271 4200 6314 4234
rect 6348 4200 6391 4234
rect 5841 3070 5884 3104
rect 5918 3070 5961 3104
rect 5841 3026 5961 3070
rect 5841 2992 5884 3026
rect 5918 2992 5961 3026
rect 5841 2948 5961 2992
rect 5841 2914 5884 2948
rect 5918 2914 5961 2948
rect 5841 2870 5961 2914
rect 5841 2836 5884 2870
rect 5918 2836 5961 2870
rect 5841 2792 5961 2836
rect 5841 2758 5884 2792
rect 5918 2758 5961 2792
rect 5841 2713 5961 2758
rect 5841 2679 5884 2713
rect 5918 2679 5961 2713
rect 5841 2634 5961 2679
rect 5841 2600 5884 2634
rect 5918 2600 5961 2634
rect 5279 1470 5322 1504
rect 5356 1470 5399 1504
rect 5279 1430 5399 1470
rect 5279 1396 5322 1430
rect 5356 1396 5399 1430
rect 5279 1250 5399 1396
rect 5279 1144 5286 1250
rect 5392 1144 5399 1250
rect 5841 1504 5961 2600
rect 6026 4064 6027 4098
rect 6061 4082 6099 4098
rect 6061 4064 6063 4082
rect 6026 4048 6063 4064
rect 6097 4064 6099 4082
rect 6133 4082 6171 4098
rect 6133 4064 6135 4082
rect 6097 4048 6135 4064
rect 6169 4064 6171 4082
rect 6205 4064 6206 4098
rect 6169 4048 6206 4064
rect 6026 4025 6206 4048
rect 6026 3991 6027 4025
rect 6061 4014 6099 4025
rect 6061 3991 6063 4014
rect 6026 3980 6063 3991
rect 6097 3991 6099 4014
rect 6133 4014 6171 4025
rect 6133 3991 6135 4014
rect 6097 3980 6135 3991
rect 6169 3991 6171 4014
rect 6205 3991 6206 4025
rect 6169 3980 6206 3991
rect 6026 3952 6206 3980
rect 6026 3918 6027 3952
rect 6061 3946 6099 3952
rect 6061 3918 6063 3946
rect 6026 3912 6063 3918
rect 6097 3918 6099 3946
rect 6133 3946 6171 3952
rect 6133 3918 6135 3946
rect 6097 3912 6135 3918
rect 6169 3918 6171 3946
rect 6205 3918 6206 3952
rect 6169 3912 6206 3918
rect 6026 3879 6206 3912
rect 6026 3845 6027 3879
rect 6061 3878 6099 3879
rect 6061 3845 6063 3878
rect 6026 3844 6063 3845
rect 6097 3845 6099 3878
rect 6133 3878 6171 3879
rect 6133 3845 6135 3878
rect 6097 3844 6135 3845
rect 6169 3845 6171 3878
rect 6205 3845 6206 3879
rect 6169 3844 6206 3845
rect 6026 3810 6206 3844
rect 6026 3806 6063 3810
rect 6026 3772 6027 3806
rect 6061 3776 6063 3806
rect 6097 3806 6135 3810
rect 6097 3776 6099 3806
rect 6061 3772 6099 3776
rect 6133 3776 6135 3806
rect 6169 3806 6206 3810
rect 6169 3776 6171 3806
rect 6133 3772 6171 3776
rect 6205 3772 6206 3806
rect 6026 3742 6206 3772
rect 6026 3733 6063 3742
rect 6026 3699 6027 3733
rect 6061 3708 6063 3733
rect 6097 3733 6135 3742
rect 6097 3708 6099 3733
rect 6061 3699 6099 3708
rect 6133 3708 6135 3733
rect 6169 3733 6206 3742
rect 6169 3708 6171 3733
rect 6133 3699 6171 3708
rect 6205 3699 6206 3733
rect 6026 3674 6206 3699
rect 6026 3660 6063 3674
rect 6026 3626 6027 3660
rect 6061 3640 6063 3660
rect 6097 3660 6135 3674
rect 6097 3640 6099 3660
rect 6061 3626 6099 3640
rect 6133 3640 6135 3660
rect 6169 3660 6206 3674
rect 6169 3640 6171 3660
rect 6133 3626 6171 3640
rect 6205 3626 6206 3660
rect 6026 3606 6206 3626
rect 6026 3587 6063 3606
rect 6026 3553 6027 3587
rect 6061 3572 6063 3587
rect 6097 3587 6135 3606
rect 6097 3572 6099 3587
rect 6061 3553 6099 3572
rect 6133 3572 6135 3587
rect 6169 3587 6206 3606
rect 6169 3572 6171 3587
rect 6133 3553 6171 3572
rect 6205 3553 6206 3587
rect 6026 3538 6206 3553
rect 6026 3514 6063 3538
rect 6026 3480 6027 3514
rect 6061 3504 6063 3514
rect 6097 3514 6135 3538
rect 6097 3504 6099 3514
rect 6061 3480 6099 3504
rect 6133 3504 6135 3514
rect 6169 3514 6206 3538
rect 6169 3504 6171 3514
rect 6133 3480 6171 3504
rect 6205 3480 6206 3514
rect 6026 3470 6206 3480
rect 6026 3441 6063 3470
rect 6026 3407 6027 3441
rect 6061 3436 6063 3441
rect 6097 3441 6135 3470
rect 6097 3436 6099 3441
rect 6061 3407 6099 3436
rect 6133 3436 6135 3441
rect 6169 3441 6206 3470
rect 6169 3436 6171 3441
rect 6133 3407 6171 3436
rect 6205 3407 6206 3441
rect 6026 3402 6206 3407
rect 6026 3368 6063 3402
rect 6097 3368 6135 3402
rect 6169 3368 6206 3402
rect 6026 3334 6027 3368
rect 6061 3334 6099 3368
rect 6133 3334 6171 3368
rect 6205 3334 6206 3368
rect 6026 3300 6063 3334
rect 6097 3300 6135 3334
rect 6169 3300 6206 3334
rect 6026 3295 6206 3300
rect 6026 3261 6027 3295
rect 6061 3266 6099 3295
rect 6061 3261 6063 3266
rect 6026 3232 6063 3261
rect 6097 3261 6099 3266
rect 6133 3266 6171 3295
rect 6133 3261 6135 3266
rect 6097 3232 6135 3261
rect 6169 3261 6171 3266
rect 6205 3261 6206 3295
rect 6169 3232 6206 3261
rect 6026 3222 6206 3232
rect 6026 3188 6027 3222
rect 6061 3198 6099 3222
rect 6061 3188 6063 3198
rect 6026 3164 6063 3188
rect 6097 3188 6099 3198
rect 6133 3198 6171 3222
rect 6133 3188 6135 3198
rect 6097 3164 6135 3188
rect 6169 3188 6171 3198
rect 6205 3188 6206 3222
rect 6169 3164 6206 3188
rect 6026 3149 6206 3164
rect 6026 3115 6027 3149
rect 6061 3115 6099 3149
rect 6133 3115 6171 3149
rect 6205 3115 6206 3149
rect 6026 3076 6206 3115
rect 6026 3042 6027 3076
rect 6061 3042 6099 3076
rect 6133 3042 6171 3076
rect 6205 3042 6206 3076
rect 6026 3003 6206 3042
rect 6026 2969 6027 3003
rect 6061 2969 6099 3003
rect 6133 2969 6171 3003
rect 6205 2969 6206 3003
rect 6026 2930 6206 2969
rect 6026 2896 6027 2930
rect 6061 2896 6099 2930
rect 6133 2896 6171 2930
rect 6205 2896 6206 2930
rect 6026 2857 6206 2896
rect 6026 2823 6027 2857
rect 6061 2823 6099 2857
rect 6133 2823 6171 2857
rect 6205 2823 6206 2857
rect 6026 2784 6206 2823
rect 6026 2750 6027 2784
rect 6061 2750 6099 2784
rect 6133 2750 6171 2784
rect 6205 2750 6206 2784
rect 6026 2711 6206 2750
rect 6026 2677 6027 2711
rect 6061 2677 6099 2711
rect 6133 2677 6171 2711
rect 6205 2677 6206 2711
rect 6026 2638 6206 2677
rect 6026 2604 6027 2638
rect 6061 2604 6099 2638
rect 6133 2604 6171 2638
rect 6205 2604 6206 2638
rect 6026 2565 6206 2604
rect 6026 2531 6027 2565
rect 6061 2531 6099 2565
rect 6133 2531 6171 2565
rect 6205 2531 6206 2565
rect 6026 2492 6206 2531
rect 6026 2458 6027 2492
rect 6061 2482 6099 2492
rect 6061 2458 6063 2482
rect 6026 2448 6063 2458
rect 6097 2458 6099 2482
rect 6133 2482 6171 2492
rect 6133 2458 6135 2482
rect 6097 2448 6135 2458
rect 6169 2458 6171 2482
rect 6205 2458 6206 2492
rect 6169 2448 6206 2458
rect 6026 2419 6206 2448
rect 6026 2385 6027 2419
rect 6061 2414 6099 2419
rect 6061 2385 6063 2414
rect 6026 2380 6063 2385
rect 6097 2385 6099 2414
rect 6133 2414 6171 2419
rect 6133 2385 6135 2414
rect 6097 2380 6135 2385
rect 6169 2385 6171 2414
rect 6205 2385 6206 2419
rect 6169 2380 6206 2385
rect 6026 2346 6206 2380
rect 6026 2312 6027 2346
rect 6061 2312 6063 2346
rect 6097 2312 6099 2346
rect 6133 2312 6135 2346
rect 6169 2312 6171 2346
rect 6205 2312 6206 2346
rect 6026 2278 6206 2312
rect 6026 2273 6063 2278
rect 6026 2239 6027 2273
rect 6061 2244 6063 2273
rect 6097 2273 6135 2278
rect 6097 2244 6099 2273
rect 6061 2239 6099 2244
rect 6133 2244 6135 2273
rect 6169 2273 6206 2278
rect 6169 2244 6171 2273
rect 6133 2239 6171 2244
rect 6205 2239 6206 2273
rect 6026 2210 6206 2239
rect 6026 2200 6063 2210
rect 6026 2166 6027 2200
rect 6061 2176 6063 2200
rect 6097 2200 6135 2210
rect 6097 2176 6099 2200
rect 6061 2166 6099 2176
rect 6133 2176 6135 2200
rect 6169 2200 6206 2210
rect 6169 2176 6171 2200
rect 6133 2166 6171 2176
rect 6205 2166 6206 2200
rect 6026 2142 6206 2166
rect 6026 2126 6063 2142
rect 6026 2092 6027 2126
rect 6061 2108 6063 2126
rect 6097 2126 6135 2142
rect 6097 2108 6099 2126
rect 6061 2092 6099 2108
rect 6133 2108 6135 2126
rect 6169 2126 6206 2142
rect 6169 2108 6171 2126
rect 6133 2092 6171 2108
rect 6205 2092 6206 2126
rect 6026 2074 6206 2092
rect 6026 2052 6063 2074
rect 6026 2018 6027 2052
rect 6061 2040 6063 2052
rect 6097 2052 6135 2074
rect 6097 2040 6099 2052
rect 6061 2018 6099 2040
rect 6133 2040 6135 2052
rect 6169 2052 6206 2074
rect 6169 2040 6171 2052
rect 6133 2018 6171 2040
rect 6205 2018 6206 2052
rect 6026 2006 6206 2018
rect 6026 1978 6063 2006
rect 6026 1944 6027 1978
rect 6061 1972 6063 1978
rect 6097 1978 6135 2006
rect 6097 1972 6099 1978
rect 6061 1944 6099 1972
rect 6133 1972 6135 1978
rect 6169 1978 6206 2006
rect 6169 1972 6171 1978
rect 6133 1944 6171 1972
rect 6205 1944 6206 1978
rect 6026 1938 6206 1944
rect 6026 1904 6063 1938
rect 6097 1904 6135 1938
rect 6169 1904 6206 1938
rect 6026 1870 6027 1904
rect 6061 1870 6099 1904
rect 6133 1870 6171 1904
rect 6205 1870 6206 1904
rect 6026 1836 6063 1870
rect 6097 1836 6135 1870
rect 6169 1836 6206 1870
rect 6026 1830 6206 1836
rect 6026 1796 6027 1830
rect 6061 1802 6099 1830
rect 6061 1796 6063 1802
rect 6026 1768 6063 1796
rect 6097 1796 6099 1802
rect 6133 1802 6171 1830
rect 6133 1796 6135 1802
rect 6097 1768 6135 1796
rect 6169 1796 6171 1802
rect 6205 1796 6206 1830
rect 6169 1768 6206 1796
rect 6026 1756 6206 1768
rect 6026 1722 6027 1756
rect 6061 1734 6099 1756
rect 6061 1722 6063 1734
rect 6026 1700 6063 1722
rect 6097 1722 6099 1734
rect 6133 1734 6171 1756
rect 6133 1722 6135 1734
rect 6097 1700 6135 1722
rect 6169 1722 6171 1734
rect 6205 1722 6206 1756
rect 6169 1700 6206 1722
rect 6026 1682 6206 1700
rect 6026 1648 6027 1682
rect 6061 1666 6099 1682
rect 6061 1648 6063 1666
rect 6026 1632 6063 1648
rect 6097 1648 6099 1666
rect 6133 1666 6171 1682
rect 6133 1648 6135 1666
rect 6097 1632 6135 1648
rect 6169 1648 6171 1666
rect 6205 1648 6206 1682
rect 6169 1632 6206 1648
rect 6026 1608 6206 1632
rect 6026 1574 6027 1608
rect 6061 1598 6099 1608
rect 6061 1574 6063 1598
rect 6026 1564 6063 1574
rect 6097 1574 6099 1598
rect 6133 1598 6171 1608
rect 6133 1574 6135 1598
rect 6097 1564 6135 1574
rect 6169 1574 6171 1598
rect 6205 1574 6206 1608
rect 6169 1564 6206 1574
rect 6026 1548 6206 1564
rect 6271 3104 6391 4200
rect 6833 4308 6953 4324
rect 6833 4274 6876 4308
rect 6910 4274 6953 4308
rect 6833 4234 6953 4274
rect 6833 4200 6876 4234
rect 6910 4200 6953 4234
rect 6271 3070 6314 3104
rect 6348 3070 6391 3104
rect 6271 3026 6391 3070
rect 6271 2992 6314 3026
rect 6348 2992 6391 3026
rect 6271 2948 6391 2992
rect 6271 2914 6314 2948
rect 6348 2914 6391 2948
rect 6271 2870 6391 2914
rect 6271 2836 6314 2870
rect 6348 2836 6391 2870
rect 6271 2792 6391 2836
rect 6271 2758 6314 2792
rect 6348 2758 6391 2792
rect 6271 2713 6391 2758
rect 6271 2679 6314 2713
rect 6348 2679 6391 2713
rect 6271 2634 6391 2679
rect 6271 2600 6314 2634
rect 6348 2600 6391 2634
rect 5841 1470 5884 1504
rect 5918 1470 5961 1504
rect 5841 1430 5961 1470
rect 5841 1396 5884 1430
rect 5918 1396 5961 1430
rect 5841 1250 5961 1396
rect 5841 1144 5848 1250
rect 5954 1144 5961 1250
rect 6271 1504 6391 2600
rect 6493 4092 6595 4118
rect 6629 4092 6731 4118
rect 6493 4082 6523 4092
rect 6701 4082 6731 4092
rect 6493 4014 6523 4048
rect 6701 4014 6731 4048
rect 6493 3946 6523 3980
rect 6701 3946 6731 3980
rect 6493 3878 6523 3912
rect 6701 3878 6731 3912
rect 6493 3810 6523 3844
rect 6701 3810 6731 3844
rect 6493 3742 6523 3776
rect 6701 3742 6731 3776
rect 6493 3674 6523 3708
rect 6701 3674 6731 3708
rect 6493 3606 6523 3640
rect 6701 3606 6731 3640
rect 6493 3538 6523 3572
rect 6701 3538 6731 3572
rect 6493 3470 6523 3504
rect 6701 3470 6731 3504
rect 6493 3402 6523 3436
rect 6701 3402 6731 3436
rect 6493 3334 6523 3368
rect 6701 3334 6731 3368
rect 6493 3266 6523 3300
rect 6701 3266 6731 3300
rect 6493 3198 6523 3232
rect 6701 3198 6731 3232
rect 6527 3164 6595 3194
rect 6629 3164 6697 3194
rect 6493 3148 6595 3164
rect 6629 3148 6731 3164
rect 6493 3108 6731 3148
rect 6493 3074 6523 3108
rect 6557 3074 6595 3108
rect 6629 3074 6667 3108
rect 6701 3074 6731 3108
rect 6493 3044 6731 3074
rect 6493 3028 6561 3044
rect 6493 2994 6523 3028
rect 6557 3010 6561 3028
rect 6595 3028 6629 3044
rect 6557 2994 6595 3010
rect 6663 3028 6731 3044
rect 6663 3010 6667 3028
rect 6629 2994 6667 3010
rect 6701 2994 6731 3028
rect 6493 2974 6731 2994
rect 6493 2948 6561 2974
rect 6493 2914 6523 2948
rect 6557 2940 6561 2948
rect 6595 2948 6629 2974
rect 6557 2914 6595 2940
rect 6663 2948 6731 2974
rect 6663 2940 6667 2948
rect 6629 2914 6667 2940
rect 6701 2914 6731 2948
rect 6493 2904 6731 2914
rect 6493 2870 6561 2904
rect 6595 2870 6629 2904
rect 6663 2870 6731 2904
rect 6493 2868 6731 2870
rect 6493 2834 6523 2868
rect 6557 2834 6595 2868
rect 6629 2834 6667 2868
rect 6701 2834 6731 2868
rect 6493 2800 6561 2834
rect 6595 2800 6629 2834
rect 6663 2800 6731 2834
rect 6493 2788 6731 2800
rect 6493 2754 6523 2788
rect 6557 2764 6595 2788
rect 6557 2754 6561 2764
rect 6493 2730 6561 2754
rect 6629 2764 6667 2788
rect 6595 2730 6629 2754
rect 6663 2754 6667 2764
rect 6701 2754 6731 2788
rect 6663 2730 6731 2754
rect 6493 2708 6731 2730
rect 6493 2674 6523 2708
rect 6557 2694 6595 2708
rect 6557 2674 6561 2694
rect 6493 2660 6561 2674
rect 6629 2694 6667 2708
rect 6595 2660 6629 2674
rect 6663 2674 6667 2694
rect 6701 2674 6731 2708
rect 6663 2660 6731 2674
rect 6493 2628 6731 2660
rect 6493 2594 6523 2628
rect 6557 2594 6595 2628
rect 6629 2594 6667 2628
rect 6701 2594 6731 2628
rect 6493 2556 6731 2594
rect 6493 2540 6595 2556
rect 6629 2540 6731 2556
rect 6527 2518 6595 2540
rect 6629 2518 6697 2540
rect 6493 2472 6523 2506
rect 6701 2472 6731 2506
rect 6493 2404 6523 2438
rect 6701 2404 6731 2438
rect 6493 2336 6523 2370
rect 6701 2336 6731 2370
rect 6493 2268 6523 2302
rect 6701 2268 6731 2302
rect 6493 2200 6523 2234
rect 6701 2200 6731 2234
rect 6493 2132 6523 2166
rect 6701 2132 6731 2166
rect 6493 2064 6523 2098
rect 6701 2064 6731 2098
rect 6493 1996 6523 2030
rect 6701 1996 6731 2030
rect 6493 1928 6523 1962
rect 6701 1928 6731 1962
rect 6493 1860 6523 1894
rect 6701 1860 6731 1894
rect 6493 1792 6523 1826
rect 6701 1792 6731 1826
rect 6493 1724 6523 1758
rect 6701 1724 6731 1758
rect 6493 1656 6523 1690
rect 6701 1656 6731 1690
rect 6493 1620 6523 1622
rect 6701 1620 6731 1622
rect 6493 1586 6595 1620
rect 6629 1586 6731 1620
rect 6493 1536 6731 1586
rect 6833 3104 6953 4200
rect 7263 4308 7383 4324
rect 7263 4274 7306 4308
rect 7340 4274 7383 4308
rect 7263 4234 7383 4274
rect 7263 4200 7306 4234
rect 7340 4200 7383 4234
rect 6833 3070 6876 3104
rect 6910 3070 6953 3104
rect 6833 3026 6953 3070
rect 6833 2992 6876 3026
rect 6910 2992 6953 3026
rect 6833 2948 6953 2992
rect 6833 2914 6876 2948
rect 6910 2914 6953 2948
rect 6833 2870 6953 2914
rect 6833 2836 6876 2870
rect 6910 2836 6953 2870
rect 6833 2792 6953 2836
rect 6833 2758 6876 2792
rect 6910 2758 6953 2792
rect 6833 2713 6953 2758
rect 6833 2679 6876 2713
rect 6910 2679 6953 2713
rect 6833 2634 6953 2679
rect 6833 2600 6876 2634
rect 6910 2600 6953 2634
rect 6271 1470 6314 1504
rect 6348 1470 6391 1504
rect 6271 1430 6391 1470
rect 6271 1396 6314 1430
rect 6348 1396 6391 1430
rect 6271 1250 6391 1396
rect 6271 1144 6278 1250
rect 6384 1144 6391 1250
rect 6833 1504 6953 2600
rect 7018 4064 7019 4098
rect 7053 4082 7091 4098
rect 7053 4064 7055 4082
rect 7018 4048 7055 4064
rect 7089 4064 7091 4082
rect 7125 4082 7163 4098
rect 7125 4064 7127 4082
rect 7089 4048 7127 4064
rect 7161 4064 7163 4082
rect 7197 4064 7198 4098
rect 7161 4048 7198 4064
rect 7018 4025 7198 4048
rect 7018 3991 7019 4025
rect 7053 4014 7091 4025
rect 7053 3991 7055 4014
rect 7018 3980 7055 3991
rect 7089 3991 7091 4014
rect 7125 4014 7163 4025
rect 7125 3991 7127 4014
rect 7089 3980 7127 3991
rect 7161 3991 7163 4014
rect 7197 3991 7198 4025
rect 7161 3980 7198 3991
rect 7018 3952 7198 3980
rect 7018 3918 7019 3952
rect 7053 3946 7091 3952
rect 7053 3918 7055 3946
rect 7018 3912 7055 3918
rect 7089 3918 7091 3946
rect 7125 3946 7163 3952
rect 7125 3918 7127 3946
rect 7089 3912 7127 3918
rect 7161 3918 7163 3946
rect 7197 3918 7198 3952
rect 7161 3912 7198 3918
rect 7018 3879 7198 3912
rect 7018 3845 7019 3879
rect 7053 3878 7091 3879
rect 7053 3845 7055 3878
rect 7018 3844 7055 3845
rect 7089 3845 7091 3878
rect 7125 3878 7163 3879
rect 7125 3845 7127 3878
rect 7089 3844 7127 3845
rect 7161 3845 7163 3878
rect 7197 3845 7198 3879
rect 7161 3844 7198 3845
rect 7018 3810 7198 3844
rect 7018 3806 7055 3810
rect 7018 3772 7019 3806
rect 7053 3776 7055 3806
rect 7089 3806 7127 3810
rect 7089 3776 7091 3806
rect 7053 3772 7091 3776
rect 7125 3776 7127 3806
rect 7161 3806 7198 3810
rect 7161 3776 7163 3806
rect 7125 3772 7163 3776
rect 7197 3772 7198 3806
rect 7018 3742 7198 3772
rect 7018 3733 7055 3742
rect 7018 3699 7019 3733
rect 7053 3708 7055 3733
rect 7089 3733 7127 3742
rect 7089 3708 7091 3733
rect 7053 3699 7091 3708
rect 7125 3708 7127 3733
rect 7161 3733 7198 3742
rect 7161 3708 7163 3733
rect 7125 3699 7163 3708
rect 7197 3699 7198 3733
rect 7018 3674 7198 3699
rect 7018 3660 7055 3674
rect 7018 3626 7019 3660
rect 7053 3640 7055 3660
rect 7089 3660 7127 3674
rect 7089 3640 7091 3660
rect 7053 3626 7091 3640
rect 7125 3640 7127 3660
rect 7161 3660 7198 3674
rect 7161 3640 7163 3660
rect 7125 3626 7163 3640
rect 7197 3626 7198 3660
rect 7018 3606 7198 3626
rect 7018 3587 7055 3606
rect 7018 3553 7019 3587
rect 7053 3572 7055 3587
rect 7089 3587 7127 3606
rect 7089 3572 7091 3587
rect 7053 3553 7091 3572
rect 7125 3572 7127 3587
rect 7161 3587 7198 3606
rect 7161 3572 7163 3587
rect 7125 3553 7163 3572
rect 7197 3553 7198 3587
rect 7018 3538 7198 3553
rect 7018 3514 7055 3538
rect 7018 3480 7019 3514
rect 7053 3504 7055 3514
rect 7089 3514 7127 3538
rect 7089 3504 7091 3514
rect 7053 3480 7091 3504
rect 7125 3504 7127 3514
rect 7161 3514 7198 3538
rect 7161 3504 7163 3514
rect 7125 3480 7163 3504
rect 7197 3480 7198 3514
rect 7018 3470 7198 3480
rect 7018 3441 7055 3470
rect 7018 3407 7019 3441
rect 7053 3436 7055 3441
rect 7089 3441 7127 3470
rect 7089 3436 7091 3441
rect 7053 3407 7091 3436
rect 7125 3436 7127 3441
rect 7161 3441 7198 3470
rect 7161 3436 7163 3441
rect 7125 3407 7163 3436
rect 7197 3407 7198 3441
rect 7018 3402 7198 3407
rect 7018 3368 7055 3402
rect 7089 3368 7127 3402
rect 7161 3368 7198 3402
rect 7018 3334 7019 3368
rect 7053 3334 7091 3368
rect 7125 3334 7163 3368
rect 7197 3334 7198 3368
rect 7018 3300 7055 3334
rect 7089 3300 7127 3334
rect 7161 3300 7198 3334
rect 7018 3295 7198 3300
rect 7018 3261 7019 3295
rect 7053 3266 7091 3295
rect 7053 3261 7055 3266
rect 7018 3232 7055 3261
rect 7089 3261 7091 3266
rect 7125 3266 7163 3295
rect 7125 3261 7127 3266
rect 7089 3232 7127 3261
rect 7161 3261 7163 3266
rect 7197 3261 7198 3295
rect 7161 3232 7198 3261
rect 7018 3222 7198 3232
rect 7018 3188 7019 3222
rect 7053 3198 7091 3222
rect 7053 3188 7055 3198
rect 7018 3164 7055 3188
rect 7089 3188 7091 3198
rect 7125 3198 7163 3222
rect 7125 3188 7127 3198
rect 7089 3164 7127 3188
rect 7161 3188 7163 3198
rect 7197 3188 7198 3222
rect 7161 3164 7198 3188
rect 7018 3149 7198 3164
rect 7018 3115 7019 3149
rect 7053 3115 7091 3149
rect 7125 3115 7163 3149
rect 7197 3115 7198 3149
rect 7018 3076 7198 3115
rect 7018 3042 7019 3076
rect 7053 3042 7091 3076
rect 7125 3042 7163 3076
rect 7197 3042 7198 3076
rect 7018 3003 7198 3042
rect 7018 2969 7019 3003
rect 7053 2969 7091 3003
rect 7125 2969 7163 3003
rect 7197 2969 7198 3003
rect 7018 2930 7198 2969
rect 7018 2896 7019 2930
rect 7053 2896 7091 2930
rect 7125 2896 7163 2930
rect 7197 2896 7198 2930
rect 7018 2857 7198 2896
rect 7018 2823 7019 2857
rect 7053 2823 7091 2857
rect 7125 2823 7163 2857
rect 7197 2823 7198 2857
rect 7018 2784 7198 2823
rect 7018 2750 7019 2784
rect 7053 2750 7091 2784
rect 7125 2750 7163 2784
rect 7197 2750 7198 2784
rect 7018 2711 7198 2750
rect 7018 2677 7019 2711
rect 7053 2677 7091 2711
rect 7125 2677 7163 2711
rect 7197 2677 7198 2711
rect 7018 2638 7198 2677
rect 7018 2604 7019 2638
rect 7053 2604 7091 2638
rect 7125 2604 7163 2638
rect 7197 2604 7198 2638
rect 7018 2565 7198 2604
rect 7018 2531 7019 2565
rect 7053 2531 7091 2565
rect 7125 2531 7163 2565
rect 7197 2531 7198 2565
rect 7018 2492 7198 2531
rect 7018 2458 7019 2492
rect 7053 2482 7091 2492
rect 7053 2458 7055 2482
rect 7018 2448 7055 2458
rect 7089 2458 7091 2482
rect 7125 2482 7163 2492
rect 7125 2458 7127 2482
rect 7089 2448 7127 2458
rect 7161 2458 7163 2482
rect 7197 2458 7198 2492
rect 7161 2448 7198 2458
rect 7018 2419 7198 2448
rect 7018 2385 7019 2419
rect 7053 2414 7091 2419
rect 7053 2385 7055 2414
rect 7018 2380 7055 2385
rect 7089 2385 7091 2414
rect 7125 2414 7163 2419
rect 7125 2385 7127 2414
rect 7089 2380 7127 2385
rect 7161 2385 7163 2414
rect 7197 2385 7198 2419
rect 7161 2380 7198 2385
rect 7018 2346 7198 2380
rect 7018 2312 7019 2346
rect 7053 2312 7055 2346
rect 7089 2312 7091 2346
rect 7125 2312 7127 2346
rect 7161 2312 7163 2346
rect 7197 2312 7198 2346
rect 7018 2278 7198 2312
rect 7018 2273 7055 2278
rect 7018 2239 7019 2273
rect 7053 2244 7055 2273
rect 7089 2273 7127 2278
rect 7089 2244 7091 2273
rect 7053 2239 7091 2244
rect 7125 2244 7127 2273
rect 7161 2273 7198 2278
rect 7161 2244 7163 2273
rect 7125 2239 7163 2244
rect 7197 2239 7198 2273
rect 7018 2210 7198 2239
rect 7018 2200 7055 2210
rect 7018 2166 7019 2200
rect 7053 2176 7055 2200
rect 7089 2200 7127 2210
rect 7089 2176 7091 2200
rect 7053 2166 7091 2176
rect 7125 2176 7127 2200
rect 7161 2200 7198 2210
rect 7161 2176 7163 2200
rect 7125 2166 7163 2176
rect 7197 2166 7198 2200
rect 7018 2142 7198 2166
rect 7018 2126 7055 2142
rect 7018 2092 7019 2126
rect 7053 2108 7055 2126
rect 7089 2126 7127 2142
rect 7089 2108 7091 2126
rect 7053 2092 7091 2108
rect 7125 2108 7127 2126
rect 7161 2126 7198 2142
rect 7161 2108 7163 2126
rect 7125 2092 7163 2108
rect 7197 2092 7198 2126
rect 7018 2074 7198 2092
rect 7018 2052 7055 2074
rect 7018 2018 7019 2052
rect 7053 2040 7055 2052
rect 7089 2052 7127 2074
rect 7089 2040 7091 2052
rect 7053 2018 7091 2040
rect 7125 2040 7127 2052
rect 7161 2052 7198 2074
rect 7161 2040 7163 2052
rect 7125 2018 7163 2040
rect 7197 2018 7198 2052
rect 7018 2006 7198 2018
rect 7018 1978 7055 2006
rect 7018 1944 7019 1978
rect 7053 1972 7055 1978
rect 7089 1978 7127 2006
rect 7089 1972 7091 1978
rect 7053 1944 7091 1972
rect 7125 1972 7127 1978
rect 7161 1978 7198 2006
rect 7161 1972 7163 1978
rect 7125 1944 7163 1972
rect 7197 1944 7198 1978
rect 7018 1938 7198 1944
rect 7018 1904 7055 1938
rect 7089 1904 7127 1938
rect 7161 1904 7198 1938
rect 7018 1870 7019 1904
rect 7053 1870 7091 1904
rect 7125 1870 7163 1904
rect 7197 1870 7198 1904
rect 7018 1836 7055 1870
rect 7089 1836 7127 1870
rect 7161 1836 7198 1870
rect 7018 1830 7198 1836
rect 7018 1796 7019 1830
rect 7053 1802 7091 1830
rect 7053 1796 7055 1802
rect 7018 1768 7055 1796
rect 7089 1796 7091 1802
rect 7125 1802 7163 1830
rect 7125 1796 7127 1802
rect 7089 1768 7127 1796
rect 7161 1796 7163 1802
rect 7197 1796 7198 1830
rect 7161 1768 7198 1796
rect 7018 1756 7198 1768
rect 7018 1722 7019 1756
rect 7053 1734 7091 1756
rect 7053 1722 7055 1734
rect 7018 1700 7055 1722
rect 7089 1722 7091 1734
rect 7125 1734 7163 1756
rect 7125 1722 7127 1734
rect 7089 1700 7127 1722
rect 7161 1722 7163 1734
rect 7197 1722 7198 1756
rect 7161 1700 7198 1722
rect 7018 1682 7198 1700
rect 7018 1648 7019 1682
rect 7053 1666 7091 1682
rect 7053 1648 7055 1666
rect 7018 1632 7055 1648
rect 7089 1648 7091 1666
rect 7125 1666 7163 1682
rect 7125 1648 7127 1666
rect 7089 1632 7127 1648
rect 7161 1648 7163 1666
rect 7197 1648 7198 1682
rect 7161 1632 7198 1648
rect 7018 1608 7198 1632
rect 7018 1574 7019 1608
rect 7053 1598 7091 1608
rect 7053 1574 7055 1598
rect 7018 1564 7055 1574
rect 7089 1574 7091 1598
rect 7125 1598 7163 1608
rect 7125 1574 7127 1598
rect 7089 1564 7127 1574
rect 7161 1574 7163 1598
rect 7197 1574 7198 1608
rect 7161 1564 7198 1574
rect 7018 1548 7198 1564
rect 7263 3104 7383 4200
rect 7825 4308 7945 4324
rect 7825 4274 7868 4308
rect 7902 4274 7945 4308
rect 7825 4234 7945 4274
rect 7825 4200 7868 4234
rect 7902 4200 7945 4234
rect 7263 3070 7306 3104
rect 7340 3070 7383 3104
rect 7263 3026 7383 3070
rect 7263 2992 7306 3026
rect 7340 2992 7383 3026
rect 7263 2948 7383 2992
rect 7263 2914 7306 2948
rect 7340 2914 7383 2948
rect 7263 2870 7383 2914
rect 7263 2836 7306 2870
rect 7340 2836 7383 2870
rect 7263 2792 7383 2836
rect 7263 2758 7306 2792
rect 7340 2758 7383 2792
rect 7263 2713 7383 2758
rect 7263 2679 7306 2713
rect 7340 2679 7383 2713
rect 7263 2634 7383 2679
rect 7263 2600 7306 2634
rect 7340 2600 7383 2634
rect 6833 1470 6876 1504
rect 6910 1470 6953 1504
rect 6833 1430 6953 1470
rect 6833 1396 6876 1430
rect 6910 1396 6953 1430
rect 6833 1250 6953 1396
rect 6833 1144 6840 1250
rect 6946 1144 6953 1250
rect 7263 1504 7383 2600
rect 7485 4092 7587 4118
rect 7621 4092 7723 4118
rect 7485 4082 7515 4092
rect 7693 4082 7723 4092
rect 7485 4014 7515 4048
rect 7693 4014 7723 4048
rect 7485 3946 7515 3980
rect 7693 3946 7723 3980
rect 7485 3878 7515 3912
rect 7693 3878 7723 3912
rect 7485 3810 7515 3844
rect 7693 3810 7723 3844
rect 7485 3742 7515 3776
rect 7693 3742 7723 3776
rect 7485 3674 7515 3708
rect 7693 3674 7723 3708
rect 7485 3606 7515 3640
rect 7693 3606 7723 3640
rect 7485 3538 7515 3572
rect 7693 3538 7723 3572
rect 7485 3470 7515 3504
rect 7693 3470 7723 3504
rect 7485 3402 7515 3436
rect 7693 3402 7723 3436
rect 7485 3334 7515 3368
rect 7693 3334 7723 3368
rect 7485 3266 7515 3300
rect 7693 3266 7723 3300
rect 7485 3198 7515 3232
rect 7693 3198 7723 3232
rect 7519 3164 7587 3194
rect 7621 3164 7689 3194
rect 7485 3148 7587 3164
rect 7621 3148 7723 3164
rect 7485 3108 7723 3148
rect 7485 3074 7515 3108
rect 7549 3074 7587 3108
rect 7621 3074 7659 3108
rect 7693 3074 7723 3108
rect 7485 3044 7723 3074
rect 7485 3028 7553 3044
rect 7485 2994 7515 3028
rect 7549 3010 7553 3028
rect 7587 3028 7621 3044
rect 7549 2994 7587 3010
rect 7655 3028 7723 3044
rect 7655 3010 7659 3028
rect 7621 2994 7659 3010
rect 7693 2994 7723 3028
rect 7485 2974 7723 2994
rect 7485 2948 7553 2974
rect 7485 2914 7515 2948
rect 7549 2940 7553 2948
rect 7587 2948 7621 2974
rect 7549 2914 7587 2940
rect 7655 2948 7723 2974
rect 7655 2940 7659 2948
rect 7621 2914 7659 2940
rect 7693 2914 7723 2948
rect 7485 2904 7723 2914
rect 7485 2870 7553 2904
rect 7587 2870 7621 2904
rect 7655 2870 7723 2904
rect 7485 2868 7723 2870
rect 7485 2834 7515 2868
rect 7549 2834 7587 2868
rect 7621 2834 7659 2868
rect 7693 2834 7723 2868
rect 7485 2800 7553 2834
rect 7587 2800 7621 2834
rect 7655 2800 7723 2834
rect 7485 2788 7723 2800
rect 7485 2754 7515 2788
rect 7549 2764 7587 2788
rect 7549 2754 7553 2764
rect 7485 2730 7553 2754
rect 7621 2764 7659 2788
rect 7587 2730 7621 2754
rect 7655 2754 7659 2764
rect 7693 2754 7723 2788
rect 7655 2730 7723 2754
rect 7485 2708 7723 2730
rect 7485 2674 7515 2708
rect 7549 2694 7587 2708
rect 7549 2674 7553 2694
rect 7485 2660 7553 2674
rect 7621 2694 7659 2708
rect 7587 2660 7621 2674
rect 7655 2674 7659 2694
rect 7693 2674 7723 2708
rect 7655 2660 7723 2674
rect 7485 2628 7723 2660
rect 7485 2594 7515 2628
rect 7549 2594 7587 2628
rect 7621 2594 7659 2628
rect 7693 2594 7723 2628
rect 7485 2556 7723 2594
rect 7485 2540 7587 2556
rect 7621 2540 7723 2556
rect 7519 2518 7587 2540
rect 7621 2518 7689 2540
rect 7485 2472 7515 2506
rect 7693 2472 7723 2506
rect 7485 2404 7515 2438
rect 7693 2404 7723 2438
rect 7485 2336 7515 2370
rect 7693 2336 7723 2370
rect 7485 2268 7515 2302
rect 7693 2268 7723 2302
rect 7485 2200 7515 2234
rect 7693 2200 7723 2234
rect 7485 2132 7515 2166
rect 7693 2132 7723 2166
rect 7485 2064 7515 2098
rect 7693 2064 7723 2098
rect 7485 1996 7515 2030
rect 7693 1996 7723 2030
rect 7485 1928 7515 1962
rect 7693 1928 7723 1962
rect 7485 1860 7515 1894
rect 7693 1860 7723 1894
rect 7485 1792 7515 1826
rect 7693 1792 7723 1826
rect 7485 1724 7515 1758
rect 7693 1724 7723 1758
rect 7485 1656 7515 1690
rect 7693 1656 7723 1690
rect 7485 1620 7515 1622
rect 7693 1620 7723 1622
rect 7485 1586 7587 1620
rect 7621 1586 7723 1620
rect 7485 1536 7723 1586
rect 7825 3104 7945 4200
rect 8255 4308 8375 4324
rect 8255 4274 8298 4308
rect 8332 4274 8375 4308
rect 8255 4234 8375 4274
rect 8255 4200 8298 4234
rect 8332 4200 8375 4234
rect 7825 3070 7868 3104
rect 7902 3070 7945 3104
rect 7825 3026 7945 3070
rect 7825 2992 7868 3026
rect 7902 2992 7945 3026
rect 7825 2948 7945 2992
rect 7825 2914 7868 2948
rect 7902 2914 7945 2948
rect 7825 2870 7945 2914
rect 7825 2836 7868 2870
rect 7902 2836 7945 2870
rect 7825 2792 7945 2836
rect 7825 2758 7868 2792
rect 7902 2758 7945 2792
rect 7825 2713 7945 2758
rect 7825 2679 7868 2713
rect 7902 2679 7945 2713
rect 7825 2634 7945 2679
rect 7825 2600 7868 2634
rect 7902 2600 7945 2634
rect 7263 1470 7306 1504
rect 7340 1470 7383 1504
rect 7263 1430 7383 1470
rect 7263 1396 7306 1430
rect 7340 1396 7383 1430
rect 7263 1250 7383 1396
rect 7263 1144 7270 1250
rect 7376 1144 7383 1250
rect 7825 1504 7945 2600
rect 8010 4064 8011 4098
rect 8045 4082 8083 4098
rect 8045 4064 8047 4082
rect 8010 4048 8047 4064
rect 8081 4064 8083 4082
rect 8117 4082 8155 4098
rect 8117 4064 8119 4082
rect 8081 4048 8119 4064
rect 8153 4064 8155 4082
rect 8189 4064 8190 4098
rect 8153 4048 8190 4064
rect 8010 4025 8190 4048
rect 8010 3991 8011 4025
rect 8045 4014 8083 4025
rect 8045 3991 8047 4014
rect 8010 3980 8047 3991
rect 8081 3991 8083 4014
rect 8117 4014 8155 4025
rect 8117 3991 8119 4014
rect 8081 3980 8119 3991
rect 8153 3991 8155 4014
rect 8189 3991 8190 4025
rect 8153 3980 8190 3991
rect 8010 3952 8190 3980
rect 8010 3918 8011 3952
rect 8045 3946 8083 3952
rect 8045 3918 8047 3946
rect 8010 3912 8047 3918
rect 8081 3918 8083 3946
rect 8117 3946 8155 3952
rect 8117 3918 8119 3946
rect 8081 3912 8119 3918
rect 8153 3918 8155 3946
rect 8189 3918 8190 3952
rect 8153 3912 8190 3918
rect 8010 3879 8190 3912
rect 8010 3845 8011 3879
rect 8045 3878 8083 3879
rect 8045 3845 8047 3878
rect 8010 3844 8047 3845
rect 8081 3845 8083 3878
rect 8117 3878 8155 3879
rect 8117 3845 8119 3878
rect 8081 3844 8119 3845
rect 8153 3845 8155 3878
rect 8189 3845 8190 3879
rect 8153 3844 8190 3845
rect 8010 3810 8190 3844
rect 8010 3806 8047 3810
rect 8010 3772 8011 3806
rect 8045 3776 8047 3806
rect 8081 3806 8119 3810
rect 8081 3776 8083 3806
rect 8045 3772 8083 3776
rect 8117 3776 8119 3806
rect 8153 3806 8190 3810
rect 8153 3776 8155 3806
rect 8117 3772 8155 3776
rect 8189 3772 8190 3806
rect 8010 3742 8190 3772
rect 8010 3733 8047 3742
rect 8010 3699 8011 3733
rect 8045 3708 8047 3733
rect 8081 3733 8119 3742
rect 8081 3708 8083 3733
rect 8045 3699 8083 3708
rect 8117 3708 8119 3733
rect 8153 3733 8190 3742
rect 8153 3708 8155 3733
rect 8117 3699 8155 3708
rect 8189 3699 8190 3733
rect 8010 3674 8190 3699
rect 8010 3660 8047 3674
rect 8010 3626 8011 3660
rect 8045 3640 8047 3660
rect 8081 3660 8119 3674
rect 8081 3640 8083 3660
rect 8045 3626 8083 3640
rect 8117 3640 8119 3660
rect 8153 3660 8190 3674
rect 8153 3640 8155 3660
rect 8117 3626 8155 3640
rect 8189 3626 8190 3660
rect 8010 3606 8190 3626
rect 8010 3587 8047 3606
rect 8010 3553 8011 3587
rect 8045 3572 8047 3587
rect 8081 3587 8119 3606
rect 8081 3572 8083 3587
rect 8045 3553 8083 3572
rect 8117 3572 8119 3587
rect 8153 3587 8190 3606
rect 8153 3572 8155 3587
rect 8117 3553 8155 3572
rect 8189 3553 8190 3587
rect 8010 3538 8190 3553
rect 8010 3514 8047 3538
rect 8010 3480 8011 3514
rect 8045 3504 8047 3514
rect 8081 3514 8119 3538
rect 8081 3504 8083 3514
rect 8045 3480 8083 3504
rect 8117 3504 8119 3514
rect 8153 3514 8190 3538
rect 8153 3504 8155 3514
rect 8117 3480 8155 3504
rect 8189 3480 8190 3514
rect 8010 3470 8190 3480
rect 8010 3441 8047 3470
rect 8010 3407 8011 3441
rect 8045 3436 8047 3441
rect 8081 3441 8119 3470
rect 8081 3436 8083 3441
rect 8045 3407 8083 3436
rect 8117 3436 8119 3441
rect 8153 3441 8190 3470
rect 8153 3436 8155 3441
rect 8117 3407 8155 3436
rect 8189 3407 8190 3441
rect 8010 3402 8190 3407
rect 8010 3368 8047 3402
rect 8081 3368 8119 3402
rect 8153 3368 8190 3402
rect 8010 3334 8011 3368
rect 8045 3334 8083 3368
rect 8117 3334 8155 3368
rect 8189 3334 8190 3368
rect 8010 3300 8047 3334
rect 8081 3300 8119 3334
rect 8153 3300 8190 3334
rect 8010 3295 8190 3300
rect 8010 3261 8011 3295
rect 8045 3266 8083 3295
rect 8045 3261 8047 3266
rect 8010 3232 8047 3261
rect 8081 3261 8083 3266
rect 8117 3266 8155 3295
rect 8117 3261 8119 3266
rect 8081 3232 8119 3261
rect 8153 3261 8155 3266
rect 8189 3261 8190 3295
rect 8153 3232 8190 3261
rect 8010 3222 8190 3232
rect 8010 3188 8011 3222
rect 8045 3198 8083 3222
rect 8045 3188 8047 3198
rect 8010 3164 8047 3188
rect 8081 3188 8083 3198
rect 8117 3198 8155 3222
rect 8117 3188 8119 3198
rect 8081 3164 8119 3188
rect 8153 3188 8155 3198
rect 8189 3188 8190 3222
rect 8153 3164 8190 3188
rect 8010 3149 8190 3164
rect 8010 3115 8011 3149
rect 8045 3115 8083 3149
rect 8117 3115 8155 3149
rect 8189 3115 8190 3149
rect 8010 3076 8190 3115
rect 8010 3042 8011 3076
rect 8045 3042 8083 3076
rect 8117 3042 8155 3076
rect 8189 3042 8190 3076
rect 8010 3003 8190 3042
rect 8010 2969 8011 3003
rect 8045 2969 8083 3003
rect 8117 2969 8155 3003
rect 8189 2969 8190 3003
rect 8010 2930 8190 2969
rect 8010 2896 8011 2930
rect 8045 2896 8083 2930
rect 8117 2896 8155 2930
rect 8189 2896 8190 2930
rect 8010 2857 8190 2896
rect 8010 2823 8011 2857
rect 8045 2823 8083 2857
rect 8117 2823 8155 2857
rect 8189 2823 8190 2857
rect 8010 2784 8190 2823
rect 8010 2750 8011 2784
rect 8045 2750 8083 2784
rect 8117 2750 8155 2784
rect 8189 2750 8190 2784
rect 8010 2711 8190 2750
rect 8010 2677 8011 2711
rect 8045 2677 8083 2711
rect 8117 2677 8155 2711
rect 8189 2677 8190 2711
rect 8010 2638 8190 2677
rect 8010 2604 8011 2638
rect 8045 2604 8083 2638
rect 8117 2604 8155 2638
rect 8189 2604 8190 2638
rect 8010 2565 8190 2604
rect 8010 2531 8011 2565
rect 8045 2531 8083 2565
rect 8117 2531 8155 2565
rect 8189 2531 8190 2565
rect 8010 2492 8190 2531
rect 8010 2458 8011 2492
rect 8045 2482 8083 2492
rect 8045 2458 8047 2482
rect 8010 2448 8047 2458
rect 8081 2458 8083 2482
rect 8117 2482 8155 2492
rect 8117 2458 8119 2482
rect 8081 2448 8119 2458
rect 8153 2458 8155 2482
rect 8189 2458 8190 2492
rect 8153 2448 8190 2458
rect 8010 2419 8190 2448
rect 8010 2385 8011 2419
rect 8045 2414 8083 2419
rect 8045 2385 8047 2414
rect 8010 2380 8047 2385
rect 8081 2385 8083 2414
rect 8117 2414 8155 2419
rect 8117 2385 8119 2414
rect 8081 2380 8119 2385
rect 8153 2385 8155 2414
rect 8189 2385 8190 2419
rect 8153 2380 8190 2385
rect 8010 2346 8190 2380
rect 8010 2312 8011 2346
rect 8045 2312 8047 2346
rect 8081 2312 8083 2346
rect 8117 2312 8119 2346
rect 8153 2312 8155 2346
rect 8189 2312 8190 2346
rect 8010 2278 8190 2312
rect 8010 2273 8047 2278
rect 8010 2239 8011 2273
rect 8045 2244 8047 2273
rect 8081 2273 8119 2278
rect 8081 2244 8083 2273
rect 8045 2239 8083 2244
rect 8117 2244 8119 2273
rect 8153 2273 8190 2278
rect 8153 2244 8155 2273
rect 8117 2239 8155 2244
rect 8189 2239 8190 2273
rect 8010 2210 8190 2239
rect 8010 2200 8047 2210
rect 8010 2166 8011 2200
rect 8045 2176 8047 2200
rect 8081 2200 8119 2210
rect 8081 2176 8083 2200
rect 8045 2166 8083 2176
rect 8117 2176 8119 2200
rect 8153 2200 8190 2210
rect 8153 2176 8155 2200
rect 8117 2166 8155 2176
rect 8189 2166 8190 2200
rect 8010 2142 8190 2166
rect 8010 2126 8047 2142
rect 8010 2092 8011 2126
rect 8045 2108 8047 2126
rect 8081 2126 8119 2142
rect 8081 2108 8083 2126
rect 8045 2092 8083 2108
rect 8117 2108 8119 2126
rect 8153 2126 8190 2142
rect 8153 2108 8155 2126
rect 8117 2092 8155 2108
rect 8189 2092 8190 2126
rect 8010 2074 8190 2092
rect 8010 2052 8047 2074
rect 8010 2018 8011 2052
rect 8045 2040 8047 2052
rect 8081 2052 8119 2074
rect 8081 2040 8083 2052
rect 8045 2018 8083 2040
rect 8117 2040 8119 2052
rect 8153 2052 8190 2074
rect 8153 2040 8155 2052
rect 8117 2018 8155 2040
rect 8189 2018 8190 2052
rect 8010 2006 8190 2018
rect 8010 1978 8047 2006
rect 8010 1944 8011 1978
rect 8045 1972 8047 1978
rect 8081 1978 8119 2006
rect 8081 1972 8083 1978
rect 8045 1944 8083 1972
rect 8117 1972 8119 1978
rect 8153 1978 8190 2006
rect 8153 1972 8155 1978
rect 8117 1944 8155 1972
rect 8189 1944 8190 1978
rect 8010 1938 8190 1944
rect 8010 1904 8047 1938
rect 8081 1904 8119 1938
rect 8153 1904 8190 1938
rect 8010 1870 8011 1904
rect 8045 1870 8083 1904
rect 8117 1870 8155 1904
rect 8189 1870 8190 1904
rect 8010 1836 8047 1870
rect 8081 1836 8119 1870
rect 8153 1836 8190 1870
rect 8010 1830 8190 1836
rect 8010 1796 8011 1830
rect 8045 1802 8083 1830
rect 8045 1796 8047 1802
rect 8010 1768 8047 1796
rect 8081 1796 8083 1802
rect 8117 1802 8155 1830
rect 8117 1796 8119 1802
rect 8081 1768 8119 1796
rect 8153 1796 8155 1802
rect 8189 1796 8190 1830
rect 8153 1768 8190 1796
rect 8010 1756 8190 1768
rect 8010 1722 8011 1756
rect 8045 1734 8083 1756
rect 8045 1722 8047 1734
rect 8010 1700 8047 1722
rect 8081 1722 8083 1734
rect 8117 1734 8155 1756
rect 8117 1722 8119 1734
rect 8081 1700 8119 1722
rect 8153 1722 8155 1734
rect 8189 1722 8190 1756
rect 8153 1700 8190 1722
rect 8010 1682 8190 1700
rect 8010 1648 8011 1682
rect 8045 1666 8083 1682
rect 8045 1648 8047 1666
rect 8010 1632 8047 1648
rect 8081 1648 8083 1666
rect 8117 1666 8155 1682
rect 8117 1648 8119 1666
rect 8081 1632 8119 1648
rect 8153 1648 8155 1666
rect 8189 1648 8190 1682
rect 8153 1632 8190 1648
rect 8010 1608 8190 1632
rect 8010 1574 8011 1608
rect 8045 1598 8083 1608
rect 8045 1574 8047 1598
rect 8010 1564 8047 1574
rect 8081 1574 8083 1598
rect 8117 1598 8155 1608
rect 8117 1574 8119 1598
rect 8081 1564 8119 1574
rect 8153 1574 8155 1598
rect 8189 1574 8190 1608
rect 8153 1564 8190 1574
rect 8010 1548 8190 1564
rect 8255 3104 8375 4200
rect 8817 4308 8937 4324
rect 8817 4274 8860 4308
rect 8894 4274 8937 4308
rect 8817 4234 8937 4274
rect 8817 4200 8860 4234
rect 8894 4200 8937 4234
rect 8255 3070 8298 3104
rect 8332 3070 8375 3104
rect 8255 3026 8375 3070
rect 8255 2992 8298 3026
rect 8332 2992 8375 3026
rect 8255 2948 8375 2992
rect 8255 2914 8298 2948
rect 8332 2914 8375 2948
rect 8255 2870 8375 2914
rect 8255 2836 8298 2870
rect 8332 2836 8375 2870
rect 8255 2792 8375 2836
rect 8255 2758 8298 2792
rect 8332 2758 8375 2792
rect 8255 2713 8375 2758
rect 8255 2679 8298 2713
rect 8332 2679 8375 2713
rect 8255 2634 8375 2679
rect 8255 2600 8298 2634
rect 8332 2600 8375 2634
rect 7825 1470 7868 1504
rect 7902 1470 7945 1504
rect 7825 1430 7945 1470
rect 7825 1396 7868 1430
rect 7902 1396 7945 1430
rect 7825 1250 7945 1396
rect 7825 1144 7832 1250
rect 7938 1144 7945 1250
rect 8255 1504 8375 2600
rect 8477 4092 8579 4118
rect 8613 4092 8715 4118
rect 8477 4082 8507 4092
rect 8685 4082 8715 4092
rect 8477 4014 8507 4048
rect 8685 4014 8715 4048
rect 8477 3946 8507 3980
rect 8685 3946 8715 3980
rect 8477 3878 8507 3912
rect 8685 3878 8715 3912
rect 8477 3810 8507 3844
rect 8685 3810 8715 3844
rect 8477 3742 8507 3776
rect 8685 3742 8715 3776
rect 8477 3674 8507 3708
rect 8685 3674 8715 3708
rect 8477 3606 8507 3640
rect 8685 3606 8715 3640
rect 8477 3538 8507 3572
rect 8685 3538 8715 3572
rect 8477 3470 8507 3504
rect 8685 3470 8715 3504
rect 8477 3402 8507 3436
rect 8685 3402 8715 3436
rect 8477 3334 8507 3368
rect 8685 3334 8715 3368
rect 8477 3266 8507 3300
rect 8685 3266 8715 3300
rect 8477 3198 8507 3232
rect 8685 3198 8715 3232
rect 8511 3164 8579 3194
rect 8613 3164 8681 3194
rect 8477 3148 8579 3164
rect 8613 3148 8715 3164
rect 8477 3108 8715 3148
rect 8477 3074 8507 3108
rect 8541 3074 8579 3108
rect 8613 3074 8651 3108
rect 8685 3074 8715 3108
rect 8477 3044 8715 3074
rect 8477 3028 8545 3044
rect 8477 2994 8507 3028
rect 8541 3010 8545 3028
rect 8579 3028 8613 3044
rect 8541 2994 8579 3010
rect 8647 3028 8715 3044
rect 8647 3010 8651 3028
rect 8613 2994 8651 3010
rect 8685 2994 8715 3028
rect 8477 2974 8715 2994
rect 8477 2948 8545 2974
rect 8477 2914 8507 2948
rect 8541 2940 8545 2948
rect 8579 2948 8613 2974
rect 8541 2914 8579 2940
rect 8647 2948 8715 2974
rect 8647 2940 8651 2948
rect 8613 2914 8651 2940
rect 8685 2914 8715 2948
rect 8477 2904 8715 2914
rect 8477 2870 8545 2904
rect 8579 2870 8613 2904
rect 8647 2870 8715 2904
rect 8477 2868 8715 2870
rect 8477 2834 8507 2868
rect 8541 2834 8579 2868
rect 8613 2834 8651 2868
rect 8685 2834 8715 2868
rect 8477 2800 8545 2834
rect 8579 2800 8613 2834
rect 8647 2800 8715 2834
rect 8477 2788 8715 2800
rect 8477 2754 8507 2788
rect 8541 2764 8579 2788
rect 8541 2754 8545 2764
rect 8477 2730 8545 2754
rect 8613 2764 8651 2788
rect 8579 2730 8613 2754
rect 8647 2754 8651 2764
rect 8685 2754 8715 2788
rect 8647 2730 8715 2754
rect 8477 2708 8715 2730
rect 8477 2674 8507 2708
rect 8541 2694 8579 2708
rect 8541 2674 8545 2694
rect 8477 2660 8545 2674
rect 8613 2694 8651 2708
rect 8579 2660 8613 2674
rect 8647 2674 8651 2694
rect 8685 2674 8715 2708
rect 8647 2660 8715 2674
rect 8477 2628 8715 2660
rect 8477 2594 8507 2628
rect 8541 2594 8579 2628
rect 8613 2594 8651 2628
rect 8685 2594 8715 2628
rect 8477 2556 8715 2594
rect 8477 2540 8579 2556
rect 8613 2540 8715 2556
rect 8511 2518 8579 2540
rect 8613 2518 8681 2540
rect 8477 2472 8507 2506
rect 8685 2472 8715 2506
rect 8477 2404 8507 2438
rect 8685 2404 8715 2438
rect 8477 2336 8507 2370
rect 8685 2336 8715 2370
rect 8477 2268 8507 2302
rect 8685 2268 8715 2302
rect 8477 2200 8507 2234
rect 8685 2200 8715 2234
rect 8477 2132 8507 2166
rect 8685 2132 8715 2166
rect 8477 2064 8507 2098
rect 8685 2064 8715 2098
rect 8477 1996 8507 2030
rect 8685 1996 8715 2030
rect 8477 1928 8507 1962
rect 8685 1928 8715 1962
rect 8477 1860 8507 1894
rect 8685 1860 8715 1894
rect 8477 1792 8507 1826
rect 8685 1792 8715 1826
rect 8477 1724 8507 1758
rect 8685 1724 8715 1758
rect 8477 1656 8507 1690
rect 8685 1656 8715 1690
rect 8477 1620 8507 1622
rect 8685 1620 8715 1622
rect 8477 1586 8579 1620
rect 8613 1586 8715 1620
rect 8477 1536 8715 1586
rect 8817 3104 8937 4200
rect 9247 4308 9367 4324
rect 9247 4274 9290 4308
rect 9324 4274 9367 4308
rect 9247 4234 9367 4274
rect 9247 4200 9290 4234
rect 9324 4200 9367 4234
rect 8817 3070 8860 3104
rect 8894 3070 8937 3104
rect 8817 3026 8937 3070
rect 8817 2992 8860 3026
rect 8894 2992 8937 3026
rect 8817 2948 8937 2992
rect 8817 2914 8860 2948
rect 8894 2914 8937 2948
rect 8817 2870 8937 2914
rect 8817 2836 8860 2870
rect 8894 2836 8937 2870
rect 8817 2792 8937 2836
rect 8817 2758 8860 2792
rect 8894 2758 8937 2792
rect 8817 2713 8937 2758
rect 8817 2679 8860 2713
rect 8894 2679 8937 2713
rect 8817 2634 8937 2679
rect 8817 2600 8860 2634
rect 8894 2600 8937 2634
rect 8255 1470 8298 1504
rect 8332 1470 8375 1504
rect 8255 1430 8375 1470
rect 8255 1396 8298 1430
rect 8332 1396 8375 1430
rect 8255 1250 8375 1396
rect 8255 1144 8262 1250
rect 8368 1144 8375 1250
rect 8817 1504 8937 2600
rect 9002 4098 9182 4099
rect 9002 4064 9003 4098
rect 9037 4082 9075 4098
rect 9037 4064 9039 4082
rect 9002 4048 9039 4064
rect 9073 4064 9075 4082
rect 9109 4082 9147 4098
rect 9109 4064 9111 4082
rect 9073 4048 9111 4064
rect 9145 4064 9147 4082
rect 9181 4064 9182 4098
rect 9145 4048 9182 4064
rect 9002 4025 9182 4048
rect 9002 3991 9003 4025
rect 9037 4014 9075 4025
rect 9037 3991 9039 4014
rect 9002 3980 9039 3991
rect 9073 3991 9075 4014
rect 9109 4014 9147 4025
rect 9109 3991 9111 4014
rect 9073 3980 9111 3991
rect 9145 3991 9147 4014
rect 9181 3991 9182 4025
rect 9145 3980 9182 3991
rect 9002 3952 9182 3980
rect 9002 3918 9003 3952
rect 9037 3946 9075 3952
rect 9037 3918 9039 3946
rect 9002 3912 9039 3918
rect 9073 3918 9075 3946
rect 9109 3946 9147 3952
rect 9109 3918 9111 3946
rect 9073 3912 9111 3918
rect 9145 3918 9147 3946
rect 9181 3918 9182 3952
rect 9145 3912 9182 3918
rect 9002 3879 9182 3912
rect 9002 3845 9003 3879
rect 9037 3878 9075 3879
rect 9037 3845 9039 3878
rect 9002 3844 9039 3845
rect 9073 3845 9075 3878
rect 9109 3878 9147 3879
rect 9109 3845 9111 3878
rect 9073 3844 9111 3845
rect 9145 3845 9147 3878
rect 9181 3845 9182 3879
rect 9145 3844 9182 3845
rect 9002 3810 9182 3844
rect 9002 3806 9039 3810
rect 9002 3772 9003 3806
rect 9037 3776 9039 3806
rect 9073 3806 9111 3810
rect 9073 3776 9075 3806
rect 9037 3772 9075 3776
rect 9109 3776 9111 3806
rect 9145 3806 9182 3810
rect 9145 3776 9147 3806
rect 9109 3772 9147 3776
rect 9181 3772 9182 3806
rect 9002 3742 9182 3772
rect 9002 3733 9039 3742
rect 9002 3699 9003 3733
rect 9037 3708 9039 3733
rect 9073 3733 9111 3742
rect 9073 3708 9075 3733
rect 9037 3699 9075 3708
rect 9109 3708 9111 3733
rect 9145 3733 9182 3742
rect 9145 3708 9147 3733
rect 9109 3699 9147 3708
rect 9181 3699 9182 3733
rect 9002 3674 9182 3699
rect 9002 3660 9039 3674
rect 9002 3626 9003 3660
rect 9037 3640 9039 3660
rect 9073 3660 9111 3674
rect 9073 3640 9075 3660
rect 9037 3626 9075 3640
rect 9109 3640 9111 3660
rect 9145 3660 9182 3674
rect 9145 3640 9147 3660
rect 9109 3626 9147 3640
rect 9181 3626 9182 3660
rect 9002 3606 9182 3626
rect 9002 3587 9039 3606
rect 9002 3553 9003 3587
rect 9037 3572 9039 3587
rect 9073 3587 9111 3606
rect 9073 3572 9075 3587
rect 9037 3553 9075 3572
rect 9109 3572 9111 3587
rect 9145 3587 9182 3606
rect 9145 3572 9147 3587
rect 9109 3553 9147 3572
rect 9181 3553 9182 3587
rect 9002 3538 9182 3553
rect 9002 3514 9039 3538
rect 9002 3480 9003 3514
rect 9037 3504 9039 3514
rect 9073 3514 9111 3538
rect 9073 3504 9075 3514
rect 9037 3480 9075 3504
rect 9109 3504 9111 3514
rect 9145 3514 9182 3538
rect 9145 3504 9147 3514
rect 9109 3480 9147 3504
rect 9181 3480 9182 3514
rect 9002 3470 9182 3480
rect 9002 3441 9039 3470
rect 9002 3407 9003 3441
rect 9037 3436 9039 3441
rect 9073 3441 9111 3470
rect 9073 3436 9075 3441
rect 9037 3407 9075 3436
rect 9109 3436 9111 3441
rect 9145 3441 9182 3470
rect 9145 3436 9147 3441
rect 9109 3407 9147 3436
rect 9181 3407 9182 3441
rect 9002 3402 9182 3407
rect 9002 3368 9039 3402
rect 9073 3368 9111 3402
rect 9145 3368 9182 3402
rect 9002 3334 9003 3368
rect 9037 3334 9075 3368
rect 9109 3334 9147 3368
rect 9181 3334 9182 3368
rect 9002 3300 9039 3334
rect 9073 3300 9111 3334
rect 9145 3300 9182 3334
rect 9002 3295 9182 3300
rect 9002 3261 9003 3295
rect 9037 3266 9075 3295
rect 9037 3261 9039 3266
rect 9002 3232 9039 3261
rect 9073 3261 9075 3266
rect 9109 3266 9147 3295
rect 9109 3261 9111 3266
rect 9073 3232 9111 3261
rect 9145 3261 9147 3266
rect 9181 3261 9182 3295
rect 9145 3232 9182 3261
rect 9002 3222 9182 3232
rect 9002 3188 9003 3222
rect 9037 3198 9075 3222
rect 9037 3188 9039 3198
rect 9002 3164 9039 3188
rect 9073 3188 9075 3198
rect 9109 3198 9147 3222
rect 9109 3188 9111 3198
rect 9073 3164 9111 3188
rect 9145 3188 9147 3198
rect 9181 3188 9182 3222
rect 9145 3164 9182 3188
rect 9002 3149 9182 3164
rect 9002 3115 9003 3149
rect 9037 3115 9075 3149
rect 9109 3115 9147 3149
rect 9181 3115 9182 3149
rect 9002 3076 9182 3115
rect 9002 3042 9003 3076
rect 9037 3042 9075 3076
rect 9109 3042 9147 3076
rect 9181 3042 9182 3076
rect 9002 3003 9182 3042
rect 9002 2969 9003 3003
rect 9037 2969 9075 3003
rect 9109 2969 9147 3003
rect 9181 2969 9182 3003
rect 9002 2930 9182 2969
rect 9002 2896 9003 2930
rect 9037 2896 9075 2930
rect 9109 2896 9147 2930
rect 9181 2896 9182 2930
rect 9002 2857 9182 2896
rect 9002 2823 9003 2857
rect 9037 2823 9075 2857
rect 9109 2823 9147 2857
rect 9181 2823 9182 2857
rect 9002 2784 9182 2823
rect 9002 2750 9003 2784
rect 9037 2750 9075 2784
rect 9109 2750 9147 2784
rect 9181 2750 9182 2784
rect 9002 2711 9182 2750
rect 9002 2677 9003 2711
rect 9037 2677 9075 2711
rect 9109 2677 9147 2711
rect 9181 2677 9182 2711
rect 9002 2638 9182 2677
rect 9002 2604 9003 2638
rect 9037 2604 9075 2638
rect 9109 2604 9147 2638
rect 9181 2604 9182 2638
rect 9002 2565 9182 2604
rect 9002 2531 9003 2565
rect 9037 2531 9075 2565
rect 9109 2531 9147 2565
rect 9181 2531 9182 2565
rect 9002 2492 9182 2531
rect 9002 2458 9003 2492
rect 9037 2482 9075 2492
rect 9037 2458 9039 2482
rect 9002 2448 9039 2458
rect 9073 2458 9075 2482
rect 9109 2482 9147 2492
rect 9109 2458 9111 2482
rect 9073 2448 9111 2458
rect 9145 2458 9147 2482
rect 9181 2458 9182 2492
rect 9145 2448 9182 2458
rect 9002 2419 9182 2448
rect 9002 2385 9003 2419
rect 9037 2414 9075 2419
rect 9037 2385 9039 2414
rect 9002 2380 9039 2385
rect 9073 2385 9075 2414
rect 9109 2414 9147 2419
rect 9109 2385 9111 2414
rect 9073 2380 9111 2385
rect 9145 2385 9147 2414
rect 9181 2385 9182 2419
rect 9145 2380 9182 2385
rect 9002 2346 9182 2380
rect 9002 2312 9003 2346
rect 9037 2312 9039 2346
rect 9073 2312 9075 2346
rect 9109 2312 9111 2346
rect 9145 2312 9147 2346
rect 9181 2312 9182 2346
rect 9002 2278 9182 2312
rect 9002 2273 9039 2278
rect 9002 2239 9003 2273
rect 9037 2244 9039 2273
rect 9073 2273 9111 2278
rect 9073 2244 9075 2273
rect 9037 2239 9075 2244
rect 9109 2244 9111 2273
rect 9145 2273 9182 2278
rect 9145 2244 9147 2273
rect 9109 2239 9147 2244
rect 9181 2239 9182 2273
rect 9002 2210 9182 2239
rect 9002 2200 9039 2210
rect 9002 2166 9003 2200
rect 9037 2176 9039 2200
rect 9073 2200 9111 2210
rect 9073 2176 9075 2200
rect 9037 2166 9075 2176
rect 9109 2176 9111 2200
rect 9145 2200 9182 2210
rect 9145 2176 9147 2200
rect 9109 2166 9147 2176
rect 9181 2166 9182 2200
rect 9002 2142 9182 2166
rect 9002 2126 9039 2142
rect 9002 2092 9003 2126
rect 9037 2108 9039 2126
rect 9073 2126 9111 2142
rect 9073 2108 9075 2126
rect 9037 2092 9075 2108
rect 9109 2108 9111 2126
rect 9145 2126 9182 2142
rect 9145 2108 9147 2126
rect 9109 2092 9147 2108
rect 9181 2092 9182 2126
rect 9002 2074 9182 2092
rect 9002 2052 9039 2074
rect 9002 2018 9003 2052
rect 9037 2040 9039 2052
rect 9073 2052 9111 2074
rect 9073 2040 9075 2052
rect 9037 2018 9075 2040
rect 9109 2040 9111 2052
rect 9145 2052 9182 2074
rect 9145 2040 9147 2052
rect 9109 2018 9147 2040
rect 9181 2018 9182 2052
rect 9002 2006 9182 2018
rect 9002 1978 9039 2006
rect 9002 1944 9003 1978
rect 9037 1972 9039 1978
rect 9073 1978 9111 2006
rect 9073 1972 9075 1978
rect 9037 1944 9075 1972
rect 9109 1972 9111 1978
rect 9145 1978 9182 2006
rect 9145 1972 9147 1978
rect 9109 1944 9147 1972
rect 9181 1944 9182 1978
rect 9002 1938 9182 1944
rect 9002 1904 9039 1938
rect 9073 1904 9111 1938
rect 9145 1904 9182 1938
rect 9002 1870 9003 1904
rect 9037 1870 9075 1904
rect 9109 1870 9147 1904
rect 9181 1870 9182 1904
rect 9002 1836 9039 1870
rect 9073 1836 9111 1870
rect 9145 1836 9182 1870
rect 9002 1830 9182 1836
rect 9002 1796 9003 1830
rect 9037 1802 9075 1830
rect 9037 1796 9039 1802
rect 9002 1768 9039 1796
rect 9073 1796 9075 1802
rect 9109 1802 9147 1830
rect 9109 1796 9111 1802
rect 9073 1768 9111 1796
rect 9145 1796 9147 1802
rect 9181 1796 9182 1830
rect 9145 1768 9182 1796
rect 9002 1756 9182 1768
rect 9002 1722 9003 1756
rect 9037 1734 9075 1756
rect 9037 1722 9039 1734
rect 9002 1700 9039 1722
rect 9073 1722 9075 1734
rect 9109 1734 9147 1756
rect 9109 1722 9111 1734
rect 9073 1700 9111 1722
rect 9145 1722 9147 1734
rect 9181 1722 9182 1756
rect 9145 1700 9182 1722
rect 9002 1682 9182 1700
rect 9002 1648 9003 1682
rect 9037 1666 9075 1682
rect 9037 1648 9039 1666
rect 9002 1632 9039 1648
rect 9073 1648 9075 1666
rect 9109 1666 9147 1682
rect 9109 1648 9111 1666
rect 9073 1632 9111 1648
rect 9145 1648 9147 1666
rect 9181 1648 9182 1682
rect 9145 1632 9182 1648
rect 9002 1608 9182 1632
rect 9002 1574 9003 1608
rect 9037 1598 9075 1608
rect 9037 1574 9039 1598
rect 9002 1564 9039 1574
rect 9073 1574 9075 1598
rect 9109 1598 9147 1608
rect 9109 1574 9111 1598
rect 9073 1564 9111 1574
rect 9145 1574 9147 1598
rect 9181 1574 9182 1608
rect 9145 1564 9182 1574
rect 9002 1548 9182 1564
rect 9247 3104 9367 4200
rect 9809 4308 9929 4324
rect 9809 4274 9852 4308
rect 9886 4274 9929 4308
rect 9809 4234 9929 4274
rect 9809 4200 9852 4234
rect 9886 4200 9929 4234
rect 9247 3070 9290 3104
rect 9324 3070 9367 3104
rect 9247 3026 9367 3070
rect 9247 2992 9290 3026
rect 9324 2992 9367 3026
rect 9247 2948 9367 2992
rect 9247 2914 9290 2948
rect 9324 2914 9367 2948
rect 9247 2870 9367 2914
rect 9247 2836 9290 2870
rect 9324 2836 9367 2870
rect 9247 2792 9367 2836
rect 9247 2758 9290 2792
rect 9324 2758 9367 2792
rect 9247 2713 9367 2758
rect 9247 2679 9290 2713
rect 9324 2679 9367 2713
rect 9247 2634 9367 2679
rect 9247 2600 9290 2634
rect 9324 2600 9367 2634
rect 8817 1470 8860 1504
rect 8894 1470 8937 1504
rect 8817 1430 8937 1470
rect 8817 1396 8860 1430
rect 8894 1396 8937 1430
rect 8817 1250 8937 1396
rect 8817 1144 8824 1250
rect 8930 1144 8937 1250
rect 9247 1504 9367 2600
rect 9469 4092 9571 4118
rect 9605 4092 9707 4118
rect 9469 4082 9499 4092
rect 9677 4082 9707 4092
rect 9469 4014 9499 4048
rect 9677 4014 9707 4048
rect 9469 3946 9499 3980
rect 9677 3946 9707 3980
rect 9469 3878 9499 3912
rect 9677 3878 9707 3912
rect 9469 3810 9499 3844
rect 9677 3810 9707 3844
rect 9469 3742 9499 3776
rect 9677 3742 9707 3776
rect 9469 3674 9499 3708
rect 9677 3674 9707 3708
rect 9469 3606 9499 3640
rect 9677 3606 9707 3640
rect 9469 3538 9499 3572
rect 9677 3538 9707 3572
rect 9469 3470 9499 3504
rect 9677 3470 9707 3504
rect 9469 3402 9499 3436
rect 9677 3402 9707 3436
rect 9469 3334 9499 3368
rect 9677 3334 9707 3368
rect 9469 3266 9499 3300
rect 9677 3266 9707 3300
rect 9469 3198 9499 3232
rect 9677 3198 9707 3232
rect 9503 3164 9571 3194
rect 9605 3164 9673 3194
rect 9469 3148 9571 3164
rect 9605 3148 9707 3164
rect 9469 3108 9707 3148
rect 9469 3074 9499 3108
rect 9533 3074 9571 3108
rect 9605 3074 9643 3108
rect 9677 3074 9707 3108
rect 9469 3044 9707 3074
rect 9469 3028 9537 3044
rect 9469 2994 9499 3028
rect 9533 3010 9537 3028
rect 9571 3028 9605 3044
rect 9533 2994 9571 3010
rect 9639 3028 9707 3044
rect 9639 3010 9643 3028
rect 9605 2994 9643 3010
rect 9677 2994 9707 3028
rect 9469 2974 9707 2994
rect 9469 2948 9537 2974
rect 9469 2914 9499 2948
rect 9533 2940 9537 2948
rect 9571 2948 9605 2974
rect 9533 2914 9571 2940
rect 9639 2948 9707 2974
rect 9639 2940 9643 2948
rect 9605 2914 9643 2940
rect 9677 2914 9707 2948
rect 9469 2904 9707 2914
rect 9469 2870 9537 2904
rect 9571 2870 9605 2904
rect 9639 2870 9707 2904
rect 9469 2868 9707 2870
rect 9469 2834 9499 2868
rect 9533 2834 9571 2868
rect 9605 2834 9643 2868
rect 9677 2834 9707 2868
rect 9469 2800 9537 2834
rect 9571 2800 9605 2834
rect 9639 2800 9707 2834
rect 9469 2788 9707 2800
rect 9469 2754 9499 2788
rect 9533 2764 9571 2788
rect 9533 2754 9537 2764
rect 9469 2730 9537 2754
rect 9605 2764 9643 2788
rect 9571 2730 9605 2754
rect 9639 2754 9643 2764
rect 9677 2754 9707 2788
rect 9639 2730 9707 2754
rect 9469 2708 9707 2730
rect 9469 2674 9499 2708
rect 9533 2694 9571 2708
rect 9533 2674 9537 2694
rect 9469 2660 9537 2674
rect 9605 2694 9643 2708
rect 9571 2660 9605 2674
rect 9639 2674 9643 2694
rect 9677 2674 9707 2708
rect 9639 2660 9707 2674
rect 9469 2628 9707 2660
rect 9469 2594 9499 2628
rect 9533 2594 9571 2628
rect 9605 2594 9643 2628
rect 9677 2594 9707 2628
rect 9469 2556 9707 2594
rect 9469 2540 9571 2556
rect 9605 2540 9707 2556
rect 9503 2518 9571 2540
rect 9605 2518 9673 2540
rect 9469 2472 9499 2506
rect 9677 2472 9707 2506
rect 9469 2404 9499 2438
rect 9677 2404 9707 2438
rect 9469 2336 9499 2370
rect 9677 2336 9707 2370
rect 9469 2268 9499 2302
rect 9677 2268 9707 2302
rect 9469 2200 9499 2234
rect 9677 2200 9707 2234
rect 9469 2132 9499 2166
rect 9677 2132 9707 2166
rect 9469 2064 9499 2098
rect 9677 2064 9707 2098
rect 9469 1996 9499 2030
rect 9677 1996 9707 2030
rect 9469 1928 9499 1962
rect 9677 1928 9707 1962
rect 9469 1860 9499 1894
rect 9677 1860 9707 1894
rect 9469 1792 9499 1826
rect 9677 1792 9707 1826
rect 9469 1724 9499 1758
rect 9677 1724 9707 1758
rect 9469 1656 9499 1690
rect 9677 1656 9707 1690
rect 9469 1620 9499 1622
rect 9677 1620 9707 1622
rect 9469 1586 9571 1620
rect 9605 1586 9707 1620
rect 9469 1536 9707 1586
rect 9809 3104 9929 4200
rect 10239 4308 10359 4324
rect 10239 4274 10282 4308
rect 10316 4274 10359 4308
rect 10239 4234 10359 4274
rect 10239 4200 10282 4234
rect 10316 4200 10359 4234
rect 9809 3070 9852 3104
rect 9886 3070 9929 3104
rect 9809 3026 9929 3070
rect 9809 2992 9852 3026
rect 9886 2992 9929 3026
rect 9809 2948 9929 2992
rect 9809 2914 9852 2948
rect 9886 2914 9929 2948
rect 9809 2870 9929 2914
rect 9809 2836 9852 2870
rect 9886 2836 9929 2870
rect 9809 2792 9929 2836
rect 9809 2758 9852 2792
rect 9886 2758 9929 2792
rect 9809 2713 9929 2758
rect 9809 2679 9852 2713
rect 9886 2679 9929 2713
rect 9809 2634 9929 2679
rect 9809 2600 9852 2634
rect 9886 2600 9929 2634
rect 9247 1470 9290 1504
rect 9324 1470 9367 1504
rect 9247 1430 9367 1470
rect 9247 1396 9290 1430
rect 9324 1396 9367 1430
rect 9247 1250 9367 1396
rect 9247 1144 9254 1250
rect 9360 1144 9367 1250
rect 9809 1504 9929 2600
rect 9994 4098 10174 4118
rect 9994 4064 9995 4098
rect 10029 4082 10067 4098
rect 10029 4064 10031 4082
rect 9994 4048 10031 4064
rect 10065 4064 10067 4082
rect 10101 4082 10139 4098
rect 10101 4064 10103 4082
rect 10065 4048 10103 4064
rect 10137 4064 10139 4082
rect 10173 4064 10174 4098
rect 10137 4048 10174 4064
rect 9994 4025 10174 4048
rect 9994 3991 9995 4025
rect 10029 4014 10067 4025
rect 10029 3991 10031 4014
rect 9994 3980 10031 3991
rect 10065 3991 10067 4014
rect 10101 4014 10139 4025
rect 10101 3991 10103 4014
rect 10065 3980 10103 3991
rect 10137 3991 10139 4014
rect 10173 3991 10174 4025
rect 10137 3980 10174 3991
rect 9994 3952 10174 3980
rect 9994 3918 9995 3952
rect 10029 3946 10067 3952
rect 10029 3918 10031 3946
rect 9994 3912 10031 3918
rect 10065 3918 10067 3946
rect 10101 3946 10139 3952
rect 10101 3918 10103 3946
rect 10065 3912 10103 3918
rect 10137 3918 10139 3946
rect 10173 3918 10174 3952
rect 10137 3912 10174 3918
rect 9994 3879 10174 3912
rect 9994 3845 9995 3879
rect 10029 3878 10067 3879
rect 10029 3845 10031 3878
rect 9994 3844 10031 3845
rect 10065 3845 10067 3878
rect 10101 3878 10139 3879
rect 10101 3845 10103 3878
rect 10065 3844 10103 3845
rect 10137 3845 10139 3878
rect 10173 3845 10174 3879
rect 10137 3844 10174 3845
rect 9994 3810 10174 3844
rect 9994 3806 10031 3810
rect 9994 3772 9995 3806
rect 10029 3776 10031 3806
rect 10065 3806 10103 3810
rect 10065 3776 10067 3806
rect 10029 3772 10067 3776
rect 10101 3776 10103 3806
rect 10137 3806 10174 3810
rect 10137 3776 10139 3806
rect 10101 3772 10139 3776
rect 10173 3772 10174 3806
rect 9994 3742 10174 3772
rect 9994 3733 10031 3742
rect 9994 3699 9995 3733
rect 10029 3708 10031 3733
rect 10065 3733 10103 3742
rect 10065 3708 10067 3733
rect 10029 3699 10067 3708
rect 10101 3708 10103 3733
rect 10137 3733 10174 3742
rect 10137 3708 10139 3733
rect 10101 3699 10139 3708
rect 10173 3699 10174 3733
rect 9994 3674 10174 3699
rect 9994 3660 10031 3674
rect 9994 3626 9995 3660
rect 10029 3640 10031 3660
rect 10065 3660 10103 3674
rect 10065 3640 10067 3660
rect 10029 3626 10067 3640
rect 10101 3640 10103 3660
rect 10137 3660 10174 3674
rect 10137 3640 10139 3660
rect 10101 3626 10139 3640
rect 10173 3626 10174 3660
rect 9994 3606 10174 3626
rect 9994 3587 10031 3606
rect 9994 3553 9995 3587
rect 10029 3572 10031 3587
rect 10065 3587 10103 3606
rect 10065 3572 10067 3587
rect 10029 3553 10067 3572
rect 10101 3572 10103 3587
rect 10137 3587 10174 3606
rect 10137 3572 10139 3587
rect 10101 3553 10139 3572
rect 10173 3553 10174 3587
rect 9994 3538 10174 3553
rect 9994 3514 10031 3538
rect 9994 3480 9995 3514
rect 10029 3504 10031 3514
rect 10065 3514 10103 3538
rect 10065 3504 10067 3514
rect 10029 3480 10067 3504
rect 10101 3504 10103 3514
rect 10137 3514 10174 3538
rect 10137 3504 10139 3514
rect 10101 3480 10139 3504
rect 10173 3480 10174 3514
rect 9994 3470 10174 3480
rect 9994 3441 10031 3470
rect 9994 3407 9995 3441
rect 10029 3436 10031 3441
rect 10065 3441 10103 3470
rect 10065 3436 10067 3441
rect 10029 3407 10067 3436
rect 10101 3436 10103 3441
rect 10137 3441 10174 3470
rect 10137 3436 10139 3441
rect 10101 3407 10139 3436
rect 10173 3407 10174 3441
rect 9994 3402 10174 3407
rect 9994 3368 10031 3402
rect 10065 3368 10103 3402
rect 10137 3368 10174 3402
rect 9994 3334 9995 3368
rect 10029 3334 10067 3368
rect 10101 3334 10139 3368
rect 10173 3334 10174 3368
rect 9994 3300 10031 3334
rect 10065 3300 10103 3334
rect 10137 3300 10174 3334
rect 9994 3295 10174 3300
rect 9994 3261 9995 3295
rect 10029 3266 10067 3295
rect 10029 3261 10031 3266
rect 9994 3232 10031 3261
rect 10065 3261 10067 3266
rect 10101 3266 10139 3295
rect 10101 3261 10103 3266
rect 10065 3232 10103 3261
rect 10137 3261 10139 3266
rect 10173 3261 10174 3295
rect 10137 3232 10174 3261
rect 9994 3222 10174 3232
rect 9994 3188 9995 3222
rect 10029 3198 10067 3222
rect 10029 3188 10031 3198
rect 9994 3164 10031 3188
rect 10065 3188 10067 3198
rect 10101 3198 10139 3222
rect 10101 3188 10103 3198
rect 10065 3164 10103 3188
rect 10137 3188 10139 3198
rect 10173 3188 10174 3222
rect 10137 3164 10174 3188
rect 9994 3149 10174 3164
rect 9994 3115 9995 3149
rect 10029 3115 10067 3149
rect 10101 3115 10139 3149
rect 10173 3115 10174 3149
rect 9994 3076 10174 3115
rect 9994 3042 9995 3076
rect 10029 3042 10067 3076
rect 10101 3042 10139 3076
rect 10173 3042 10174 3076
rect 9994 3003 10174 3042
rect 9994 2969 9995 3003
rect 10029 2969 10067 3003
rect 10101 2969 10139 3003
rect 10173 2969 10174 3003
rect 9994 2930 10174 2969
rect 9994 2896 9995 2930
rect 10029 2896 10067 2930
rect 10101 2896 10139 2930
rect 10173 2896 10174 2930
rect 9994 2857 10174 2896
rect 9994 2823 9995 2857
rect 10029 2823 10067 2857
rect 10101 2823 10139 2857
rect 10173 2823 10174 2857
rect 9994 2784 10174 2823
rect 9994 2750 9995 2784
rect 10029 2750 10067 2784
rect 10101 2750 10139 2784
rect 10173 2750 10174 2784
rect 9994 2711 10174 2750
rect 9994 2677 9995 2711
rect 10029 2677 10067 2711
rect 10101 2677 10139 2711
rect 10173 2677 10174 2711
rect 9994 2638 10174 2677
rect 9994 2604 9995 2638
rect 10029 2604 10067 2638
rect 10101 2604 10139 2638
rect 10173 2604 10174 2638
rect 9994 2565 10174 2604
rect 9994 2531 9995 2565
rect 10029 2531 10067 2565
rect 10101 2531 10139 2565
rect 10173 2531 10174 2565
rect 9994 2492 10174 2531
rect 9994 2458 9995 2492
rect 10029 2482 10067 2492
rect 10029 2458 10031 2482
rect 9994 2448 10031 2458
rect 10065 2458 10067 2482
rect 10101 2482 10139 2492
rect 10101 2458 10103 2482
rect 10065 2448 10103 2458
rect 10137 2458 10139 2482
rect 10173 2458 10174 2492
rect 10137 2448 10174 2458
rect 9994 2419 10174 2448
rect 9994 2385 9995 2419
rect 10029 2414 10067 2419
rect 10029 2385 10031 2414
rect 9994 2380 10031 2385
rect 10065 2385 10067 2414
rect 10101 2414 10139 2419
rect 10101 2385 10103 2414
rect 10065 2380 10103 2385
rect 10137 2385 10139 2414
rect 10173 2385 10174 2419
rect 10137 2380 10174 2385
rect 9994 2346 10174 2380
rect 9994 2312 9995 2346
rect 10029 2312 10031 2346
rect 10065 2312 10067 2346
rect 10101 2312 10103 2346
rect 10137 2312 10139 2346
rect 10173 2312 10174 2346
rect 9994 2278 10174 2312
rect 9994 2273 10031 2278
rect 9994 2239 9995 2273
rect 10029 2244 10031 2273
rect 10065 2273 10103 2278
rect 10065 2244 10067 2273
rect 10029 2239 10067 2244
rect 10101 2244 10103 2273
rect 10137 2273 10174 2278
rect 10137 2244 10139 2273
rect 10101 2239 10139 2244
rect 10173 2239 10174 2273
rect 9994 2210 10174 2239
rect 9994 2200 10031 2210
rect 9994 2166 9995 2200
rect 10029 2176 10031 2200
rect 10065 2200 10103 2210
rect 10065 2176 10067 2200
rect 10029 2166 10067 2176
rect 10101 2176 10103 2200
rect 10137 2200 10174 2210
rect 10137 2176 10139 2200
rect 10101 2166 10139 2176
rect 10173 2166 10174 2200
rect 9994 2142 10174 2166
rect 9994 2126 10031 2142
rect 9994 2092 9995 2126
rect 10029 2108 10031 2126
rect 10065 2126 10103 2142
rect 10065 2108 10067 2126
rect 10029 2092 10067 2108
rect 10101 2108 10103 2126
rect 10137 2126 10174 2142
rect 10137 2108 10139 2126
rect 10101 2092 10139 2108
rect 10173 2092 10174 2126
rect 9994 2074 10174 2092
rect 9994 2052 10031 2074
rect 9994 2018 9995 2052
rect 10029 2040 10031 2052
rect 10065 2052 10103 2074
rect 10065 2040 10067 2052
rect 10029 2018 10067 2040
rect 10101 2040 10103 2052
rect 10137 2052 10174 2074
rect 10137 2040 10139 2052
rect 10101 2018 10139 2040
rect 10173 2018 10174 2052
rect 9994 2006 10174 2018
rect 9994 1978 10031 2006
rect 9994 1944 9995 1978
rect 10029 1972 10031 1978
rect 10065 1978 10103 2006
rect 10065 1972 10067 1978
rect 10029 1944 10067 1972
rect 10101 1972 10103 1978
rect 10137 1978 10174 2006
rect 10137 1972 10139 1978
rect 10101 1944 10139 1972
rect 10173 1944 10174 1978
rect 9994 1938 10174 1944
rect 9994 1904 10031 1938
rect 10065 1904 10103 1938
rect 10137 1904 10174 1938
rect 9994 1870 9995 1904
rect 10029 1870 10067 1904
rect 10101 1870 10139 1904
rect 10173 1870 10174 1904
rect 9994 1836 10031 1870
rect 10065 1836 10103 1870
rect 10137 1836 10174 1870
rect 9994 1830 10174 1836
rect 9994 1796 9995 1830
rect 10029 1802 10067 1830
rect 10029 1796 10031 1802
rect 9994 1768 10031 1796
rect 10065 1796 10067 1802
rect 10101 1802 10139 1830
rect 10101 1796 10103 1802
rect 10065 1768 10103 1796
rect 10137 1796 10139 1802
rect 10173 1796 10174 1830
rect 10137 1768 10174 1796
rect 9994 1756 10174 1768
rect 9994 1722 9995 1756
rect 10029 1734 10067 1756
rect 10029 1722 10031 1734
rect 9994 1700 10031 1722
rect 10065 1722 10067 1734
rect 10101 1734 10139 1756
rect 10101 1722 10103 1734
rect 10065 1700 10103 1722
rect 10137 1722 10139 1734
rect 10173 1722 10174 1756
rect 10137 1700 10174 1722
rect 9994 1682 10174 1700
rect 9994 1648 9995 1682
rect 10029 1666 10067 1682
rect 10029 1648 10031 1666
rect 9994 1632 10031 1648
rect 10065 1648 10067 1666
rect 10101 1666 10139 1682
rect 10101 1648 10103 1666
rect 10065 1632 10103 1648
rect 10137 1648 10139 1666
rect 10173 1648 10174 1682
rect 10137 1632 10174 1648
rect 9994 1608 10174 1632
rect 9994 1574 9995 1608
rect 10029 1598 10067 1608
rect 10029 1574 10031 1598
rect 9994 1564 10031 1574
rect 10065 1574 10067 1598
rect 10101 1598 10139 1608
rect 10101 1574 10103 1598
rect 10065 1564 10103 1574
rect 10137 1574 10139 1598
rect 10173 1574 10174 1608
rect 10137 1564 10174 1574
rect 9994 1548 10174 1564
rect 10239 3104 10359 4200
rect 10801 4308 10921 4324
rect 10801 4274 10844 4308
rect 10878 4274 10921 4308
rect 10801 4234 10921 4274
rect 10801 4200 10844 4234
rect 10878 4200 10921 4234
rect 10239 3070 10282 3104
rect 10316 3070 10359 3104
rect 10239 3026 10359 3070
rect 10239 2992 10282 3026
rect 10316 2992 10359 3026
rect 10239 2948 10359 2992
rect 10239 2914 10282 2948
rect 10316 2914 10359 2948
rect 10239 2870 10359 2914
rect 10239 2836 10282 2870
rect 10316 2836 10359 2870
rect 10239 2792 10359 2836
rect 10239 2758 10282 2792
rect 10316 2758 10359 2792
rect 10239 2713 10359 2758
rect 10239 2679 10282 2713
rect 10316 2679 10359 2713
rect 10239 2634 10359 2679
rect 10239 2600 10282 2634
rect 10316 2600 10359 2634
rect 9809 1470 9852 1504
rect 9886 1470 9929 1504
rect 9809 1430 9929 1470
rect 9809 1396 9852 1430
rect 9886 1396 9929 1430
rect 9809 1250 9929 1396
rect 9809 1144 9816 1250
rect 9922 1144 9929 1250
rect 10239 1504 10359 2600
rect 10461 4118 10699 4130
rect 10461 4092 10563 4118
rect 10597 4092 10699 4118
rect 10461 4082 10491 4092
rect 10669 4082 10699 4092
rect 10461 4014 10491 4048
rect 10669 4014 10699 4048
rect 10461 3946 10491 3980
rect 10669 3946 10699 3980
rect 10461 3878 10491 3912
rect 10669 3878 10699 3912
rect 10461 3810 10491 3844
rect 10669 3810 10699 3844
rect 10461 3742 10491 3776
rect 10669 3742 10699 3776
rect 10461 3674 10491 3708
rect 10669 3674 10699 3708
rect 10461 3606 10491 3640
rect 10669 3606 10699 3640
rect 10461 3538 10491 3572
rect 10669 3538 10699 3572
rect 10461 3470 10491 3504
rect 10669 3470 10699 3504
rect 10461 3402 10491 3436
rect 10669 3402 10699 3436
rect 10461 3334 10491 3368
rect 10669 3334 10699 3368
rect 10461 3266 10491 3300
rect 10669 3266 10699 3300
rect 10461 3198 10491 3232
rect 10669 3198 10699 3232
rect 10495 3164 10563 3194
rect 10597 3164 10665 3194
rect 10461 3148 10563 3164
rect 10597 3148 10699 3164
rect 10461 3108 10699 3148
rect 10461 3074 10491 3108
rect 10525 3074 10563 3108
rect 10597 3074 10635 3108
rect 10669 3074 10699 3108
rect 10461 3044 10699 3074
rect 10461 3028 10529 3044
rect 10461 2994 10491 3028
rect 10525 3010 10529 3028
rect 10563 3028 10597 3044
rect 10525 2994 10563 3010
rect 10631 3028 10699 3044
rect 10631 3010 10635 3028
rect 10597 2994 10635 3010
rect 10669 2994 10699 3028
rect 10461 2974 10699 2994
rect 10461 2948 10529 2974
rect 10461 2914 10491 2948
rect 10525 2940 10529 2948
rect 10563 2948 10597 2974
rect 10525 2914 10563 2940
rect 10631 2948 10699 2974
rect 10631 2940 10635 2948
rect 10597 2914 10635 2940
rect 10669 2914 10699 2948
rect 10461 2904 10699 2914
rect 10461 2870 10529 2904
rect 10563 2870 10597 2904
rect 10631 2870 10699 2904
rect 10461 2868 10699 2870
rect 10461 2834 10491 2868
rect 10525 2834 10563 2868
rect 10597 2834 10635 2868
rect 10669 2834 10699 2868
rect 10461 2800 10529 2834
rect 10563 2800 10597 2834
rect 10631 2800 10699 2834
rect 10461 2788 10699 2800
rect 10461 2754 10491 2788
rect 10525 2764 10563 2788
rect 10525 2754 10529 2764
rect 10461 2730 10529 2754
rect 10597 2764 10635 2788
rect 10563 2730 10597 2754
rect 10631 2754 10635 2764
rect 10669 2754 10699 2788
rect 10631 2730 10699 2754
rect 10461 2708 10699 2730
rect 10461 2674 10491 2708
rect 10525 2694 10563 2708
rect 10525 2674 10529 2694
rect 10461 2660 10529 2674
rect 10597 2694 10635 2708
rect 10563 2660 10597 2674
rect 10631 2674 10635 2694
rect 10669 2674 10699 2708
rect 10631 2660 10699 2674
rect 10461 2628 10699 2660
rect 10461 2594 10491 2628
rect 10525 2594 10563 2628
rect 10597 2594 10635 2628
rect 10669 2594 10699 2628
rect 10461 2556 10699 2594
rect 10461 2540 10563 2556
rect 10597 2540 10699 2556
rect 10495 2518 10563 2540
rect 10597 2518 10665 2540
rect 10461 2472 10491 2506
rect 10669 2472 10699 2506
rect 10461 2404 10491 2438
rect 10669 2404 10699 2438
rect 10461 2336 10491 2370
rect 10669 2336 10699 2370
rect 10461 2268 10491 2302
rect 10669 2268 10699 2302
rect 10461 2200 10491 2234
rect 10669 2200 10699 2234
rect 10461 2132 10491 2166
rect 10669 2132 10699 2166
rect 10461 2064 10491 2098
rect 10669 2064 10699 2098
rect 10461 1996 10491 2030
rect 10669 1996 10699 2030
rect 10461 1928 10491 1962
rect 10669 1928 10699 1962
rect 10461 1860 10491 1894
rect 10669 1860 10699 1894
rect 10461 1792 10491 1826
rect 10669 1792 10699 1826
rect 10461 1724 10491 1758
rect 10669 1724 10699 1758
rect 10461 1656 10491 1690
rect 10669 1656 10699 1690
rect 10461 1620 10491 1622
rect 10669 1620 10699 1622
rect 10461 1586 10563 1620
rect 10597 1586 10699 1620
rect 10461 1536 10699 1586
rect 10801 3104 10921 4200
rect 11231 4308 11351 4324
rect 11231 4274 11274 4308
rect 11308 4274 11351 4308
rect 11231 4234 11351 4274
rect 11231 4200 11274 4234
rect 11308 4200 11351 4234
rect 10801 3070 10844 3104
rect 10878 3070 10921 3104
rect 10801 3026 10921 3070
rect 10801 2992 10844 3026
rect 10878 2992 10921 3026
rect 10801 2948 10921 2992
rect 10801 2914 10844 2948
rect 10878 2914 10921 2948
rect 10801 2870 10921 2914
rect 10801 2836 10844 2870
rect 10878 2836 10921 2870
rect 10801 2792 10921 2836
rect 10801 2758 10844 2792
rect 10878 2758 10921 2792
rect 10801 2713 10921 2758
rect 10801 2679 10844 2713
rect 10878 2679 10921 2713
rect 10801 2634 10921 2679
rect 10801 2600 10844 2634
rect 10878 2600 10921 2634
rect 10239 1470 10282 1504
rect 10316 1470 10359 1504
rect 10239 1430 10359 1470
rect 10239 1396 10282 1430
rect 10316 1396 10359 1430
rect 10239 1250 10359 1396
rect 10239 1144 10246 1250
rect 10352 1144 10359 1250
rect 10801 1504 10921 2600
rect 10986 4064 10987 4098
rect 11021 4082 11059 4098
rect 11021 4064 11023 4082
rect 10986 4048 11023 4064
rect 11057 4064 11059 4082
rect 11093 4082 11131 4098
rect 11093 4064 11095 4082
rect 11057 4048 11095 4064
rect 11129 4064 11131 4082
rect 11165 4064 11166 4098
rect 11129 4048 11166 4064
rect 10986 4025 11166 4048
rect 10986 3991 10987 4025
rect 11021 4014 11059 4025
rect 11021 3991 11023 4014
rect 10986 3980 11023 3991
rect 11057 3991 11059 4014
rect 11093 4014 11131 4025
rect 11093 3991 11095 4014
rect 11057 3980 11095 3991
rect 11129 3991 11131 4014
rect 11165 3991 11166 4025
rect 11129 3980 11166 3991
rect 10986 3952 11166 3980
rect 10986 3918 10987 3952
rect 11021 3946 11059 3952
rect 11021 3918 11023 3946
rect 10986 3912 11023 3918
rect 11057 3918 11059 3946
rect 11093 3946 11131 3952
rect 11093 3918 11095 3946
rect 11057 3912 11095 3918
rect 11129 3918 11131 3946
rect 11165 3918 11166 3952
rect 11129 3912 11166 3918
rect 10986 3879 11166 3912
rect 10986 3845 10987 3879
rect 11021 3878 11059 3879
rect 11021 3845 11023 3878
rect 10986 3844 11023 3845
rect 11057 3845 11059 3878
rect 11093 3878 11131 3879
rect 11093 3845 11095 3878
rect 11057 3844 11095 3845
rect 11129 3845 11131 3878
rect 11165 3845 11166 3879
rect 11129 3844 11166 3845
rect 10986 3810 11166 3844
rect 10986 3806 11023 3810
rect 10986 3772 10987 3806
rect 11021 3776 11023 3806
rect 11057 3806 11095 3810
rect 11057 3776 11059 3806
rect 11021 3772 11059 3776
rect 11093 3776 11095 3806
rect 11129 3806 11166 3810
rect 11129 3776 11131 3806
rect 11093 3772 11131 3776
rect 11165 3772 11166 3806
rect 10986 3742 11166 3772
rect 10986 3733 11023 3742
rect 10986 3699 10987 3733
rect 11021 3708 11023 3733
rect 11057 3733 11095 3742
rect 11057 3708 11059 3733
rect 11021 3699 11059 3708
rect 11093 3708 11095 3733
rect 11129 3733 11166 3742
rect 11129 3708 11131 3733
rect 11093 3699 11131 3708
rect 11165 3699 11166 3733
rect 10986 3674 11166 3699
rect 10986 3660 11023 3674
rect 10986 3626 10987 3660
rect 11021 3640 11023 3660
rect 11057 3660 11095 3674
rect 11057 3640 11059 3660
rect 11021 3626 11059 3640
rect 11093 3640 11095 3660
rect 11129 3660 11166 3674
rect 11129 3640 11131 3660
rect 11093 3626 11131 3640
rect 11165 3626 11166 3660
rect 10986 3606 11166 3626
rect 10986 3587 11023 3606
rect 10986 3553 10987 3587
rect 11021 3572 11023 3587
rect 11057 3587 11095 3606
rect 11057 3572 11059 3587
rect 11021 3553 11059 3572
rect 11093 3572 11095 3587
rect 11129 3587 11166 3606
rect 11129 3572 11131 3587
rect 11093 3553 11131 3572
rect 11165 3553 11166 3587
rect 10986 3538 11166 3553
rect 10986 3514 11023 3538
rect 10986 3480 10987 3514
rect 11021 3504 11023 3514
rect 11057 3514 11095 3538
rect 11057 3504 11059 3514
rect 11021 3480 11059 3504
rect 11093 3504 11095 3514
rect 11129 3514 11166 3538
rect 11129 3504 11131 3514
rect 11093 3480 11131 3504
rect 11165 3480 11166 3514
rect 10986 3470 11166 3480
rect 10986 3441 11023 3470
rect 10986 3407 10987 3441
rect 11021 3436 11023 3441
rect 11057 3441 11095 3470
rect 11057 3436 11059 3441
rect 11021 3407 11059 3436
rect 11093 3436 11095 3441
rect 11129 3441 11166 3470
rect 11129 3436 11131 3441
rect 11093 3407 11131 3436
rect 11165 3407 11166 3441
rect 10986 3402 11166 3407
rect 10986 3368 11023 3402
rect 11057 3368 11095 3402
rect 11129 3368 11166 3402
rect 10986 3334 10987 3368
rect 11021 3334 11059 3368
rect 11093 3334 11131 3368
rect 11165 3334 11166 3368
rect 10986 3300 11023 3334
rect 11057 3300 11095 3334
rect 11129 3300 11166 3334
rect 10986 3295 11166 3300
rect 10986 3261 10987 3295
rect 11021 3266 11059 3295
rect 11021 3261 11023 3266
rect 10986 3232 11023 3261
rect 11057 3261 11059 3266
rect 11093 3266 11131 3295
rect 11093 3261 11095 3266
rect 11057 3232 11095 3261
rect 11129 3261 11131 3266
rect 11165 3261 11166 3295
rect 11129 3232 11166 3261
rect 10986 3222 11166 3232
rect 10986 3188 10987 3222
rect 11021 3198 11059 3222
rect 11021 3188 11023 3198
rect 10986 3164 11023 3188
rect 11057 3188 11059 3198
rect 11093 3198 11131 3222
rect 11093 3188 11095 3198
rect 11057 3164 11095 3188
rect 11129 3188 11131 3198
rect 11165 3188 11166 3222
rect 11129 3164 11166 3188
rect 10986 3149 11166 3164
rect 10986 3115 10987 3149
rect 11021 3115 11059 3149
rect 11093 3115 11131 3149
rect 11165 3115 11166 3149
rect 10986 3076 11166 3115
rect 10986 3042 10987 3076
rect 11021 3042 11059 3076
rect 11093 3042 11131 3076
rect 11165 3042 11166 3076
rect 10986 3003 11166 3042
rect 10986 2969 10987 3003
rect 11021 2969 11059 3003
rect 11093 2969 11131 3003
rect 11165 2969 11166 3003
rect 10986 2930 11166 2969
rect 10986 2896 10987 2930
rect 11021 2896 11059 2930
rect 11093 2896 11131 2930
rect 11165 2896 11166 2930
rect 10986 2857 11166 2896
rect 10986 2823 10987 2857
rect 11021 2823 11059 2857
rect 11093 2823 11131 2857
rect 11165 2823 11166 2857
rect 10986 2784 11166 2823
rect 10986 2750 10987 2784
rect 11021 2750 11059 2784
rect 11093 2750 11131 2784
rect 11165 2750 11166 2784
rect 10986 2711 11166 2750
rect 10986 2677 10987 2711
rect 11021 2677 11059 2711
rect 11093 2677 11131 2711
rect 11165 2677 11166 2711
rect 10986 2638 11166 2677
rect 10986 2604 10987 2638
rect 11021 2604 11059 2638
rect 11093 2604 11131 2638
rect 11165 2604 11166 2638
rect 10986 2565 11166 2604
rect 10986 2531 10987 2565
rect 11021 2531 11059 2565
rect 11093 2531 11131 2565
rect 11165 2531 11166 2565
rect 10986 2492 11166 2531
rect 10986 2458 10987 2492
rect 11021 2482 11059 2492
rect 11021 2458 11023 2482
rect 10986 2448 11023 2458
rect 11057 2458 11059 2482
rect 11093 2482 11131 2492
rect 11093 2458 11095 2482
rect 11057 2448 11095 2458
rect 11129 2458 11131 2482
rect 11165 2458 11166 2492
rect 11129 2448 11166 2458
rect 10986 2419 11166 2448
rect 10986 2385 10987 2419
rect 11021 2414 11059 2419
rect 11021 2385 11023 2414
rect 10986 2380 11023 2385
rect 11057 2385 11059 2414
rect 11093 2414 11131 2419
rect 11093 2385 11095 2414
rect 11057 2380 11095 2385
rect 11129 2385 11131 2414
rect 11165 2385 11166 2419
rect 11129 2380 11166 2385
rect 10986 2346 11166 2380
rect 10986 2312 10987 2346
rect 11021 2312 11023 2346
rect 11057 2312 11059 2346
rect 11093 2312 11095 2346
rect 11129 2312 11131 2346
rect 11165 2312 11166 2346
rect 10986 2278 11166 2312
rect 10986 2273 11023 2278
rect 10986 2239 10987 2273
rect 11021 2244 11023 2273
rect 11057 2273 11095 2278
rect 11057 2244 11059 2273
rect 11021 2239 11059 2244
rect 11093 2244 11095 2273
rect 11129 2273 11166 2278
rect 11129 2244 11131 2273
rect 11093 2239 11131 2244
rect 11165 2239 11166 2273
rect 10986 2210 11166 2239
rect 10986 2200 11023 2210
rect 10986 2166 10987 2200
rect 11021 2176 11023 2200
rect 11057 2200 11095 2210
rect 11057 2176 11059 2200
rect 11021 2166 11059 2176
rect 11093 2176 11095 2200
rect 11129 2200 11166 2210
rect 11129 2176 11131 2200
rect 11093 2166 11131 2176
rect 11165 2166 11166 2200
rect 10986 2142 11166 2166
rect 10986 2126 11023 2142
rect 10986 2092 10987 2126
rect 11021 2108 11023 2126
rect 11057 2126 11095 2142
rect 11057 2108 11059 2126
rect 11021 2092 11059 2108
rect 11093 2108 11095 2126
rect 11129 2126 11166 2142
rect 11129 2108 11131 2126
rect 11093 2092 11131 2108
rect 11165 2092 11166 2126
rect 10986 2074 11166 2092
rect 10986 2052 11023 2074
rect 10986 2018 10987 2052
rect 11021 2040 11023 2052
rect 11057 2052 11095 2074
rect 11057 2040 11059 2052
rect 11021 2018 11059 2040
rect 11093 2040 11095 2052
rect 11129 2052 11166 2074
rect 11129 2040 11131 2052
rect 11093 2018 11131 2040
rect 11165 2018 11166 2052
rect 10986 2006 11166 2018
rect 10986 1978 11023 2006
rect 10986 1944 10987 1978
rect 11021 1972 11023 1978
rect 11057 1978 11095 2006
rect 11057 1972 11059 1978
rect 11021 1944 11059 1972
rect 11093 1972 11095 1978
rect 11129 1978 11166 2006
rect 11129 1972 11131 1978
rect 11093 1944 11131 1972
rect 11165 1944 11166 1978
rect 10986 1938 11166 1944
rect 10986 1904 11023 1938
rect 11057 1904 11095 1938
rect 11129 1904 11166 1938
rect 10986 1870 10987 1904
rect 11021 1870 11059 1904
rect 11093 1870 11131 1904
rect 11165 1870 11166 1904
rect 10986 1836 11023 1870
rect 11057 1836 11095 1870
rect 11129 1836 11166 1870
rect 10986 1830 11166 1836
rect 10986 1796 10987 1830
rect 11021 1802 11059 1830
rect 11021 1796 11023 1802
rect 10986 1768 11023 1796
rect 11057 1796 11059 1802
rect 11093 1802 11131 1830
rect 11093 1796 11095 1802
rect 11057 1768 11095 1796
rect 11129 1796 11131 1802
rect 11165 1796 11166 1830
rect 11129 1768 11166 1796
rect 10986 1756 11166 1768
rect 10986 1722 10987 1756
rect 11021 1734 11059 1756
rect 11021 1722 11023 1734
rect 10986 1700 11023 1722
rect 11057 1722 11059 1734
rect 11093 1734 11131 1756
rect 11093 1722 11095 1734
rect 11057 1700 11095 1722
rect 11129 1722 11131 1734
rect 11165 1722 11166 1756
rect 11129 1700 11166 1722
rect 10986 1682 11166 1700
rect 10986 1648 10987 1682
rect 11021 1666 11059 1682
rect 11021 1648 11023 1666
rect 10986 1632 11023 1648
rect 11057 1648 11059 1666
rect 11093 1666 11131 1682
rect 11093 1648 11095 1666
rect 11057 1632 11095 1648
rect 11129 1648 11131 1666
rect 11165 1648 11166 1682
rect 11129 1632 11166 1648
rect 10986 1608 11166 1632
rect 10986 1574 10987 1608
rect 11021 1598 11059 1608
rect 11021 1574 11023 1598
rect 10986 1564 11023 1574
rect 11057 1574 11059 1598
rect 11093 1598 11131 1608
rect 11093 1574 11095 1598
rect 11057 1564 11095 1574
rect 11129 1574 11131 1598
rect 11165 1574 11166 1608
rect 11129 1564 11166 1574
rect 10986 1548 11166 1564
rect 11231 3104 11351 4200
rect 11793 4308 11913 4324
rect 11793 4274 11836 4308
rect 11870 4274 11913 4308
rect 11793 4234 11913 4274
rect 11793 4200 11836 4234
rect 11870 4200 11913 4234
rect 11231 3070 11274 3104
rect 11308 3070 11351 3104
rect 11231 3026 11351 3070
rect 11231 2992 11274 3026
rect 11308 2992 11351 3026
rect 11231 2948 11351 2992
rect 11231 2914 11274 2948
rect 11308 2914 11351 2948
rect 11231 2870 11351 2914
rect 11231 2836 11274 2870
rect 11308 2836 11351 2870
rect 11231 2792 11351 2836
rect 11231 2758 11274 2792
rect 11308 2758 11351 2792
rect 11231 2713 11351 2758
rect 11231 2679 11274 2713
rect 11308 2679 11351 2713
rect 11231 2634 11351 2679
rect 11231 2600 11274 2634
rect 11308 2600 11351 2634
rect 10801 1470 10844 1504
rect 10878 1470 10921 1504
rect 10801 1430 10921 1470
rect 10801 1396 10844 1430
rect 10878 1396 10921 1430
rect 10801 1250 10921 1396
rect 10801 1144 10808 1250
rect 10914 1144 10921 1250
rect 11231 1504 11351 2600
rect 11453 4092 11555 4118
rect 11589 4092 11691 4118
rect 11453 4082 11483 4092
rect 11661 4082 11691 4092
rect 11453 4014 11483 4048
rect 11661 4014 11691 4048
rect 11453 3946 11483 3980
rect 11661 3946 11691 3980
rect 11453 3878 11483 3912
rect 11661 3878 11691 3912
rect 11453 3810 11483 3844
rect 11661 3810 11691 3844
rect 11453 3742 11483 3776
rect 11661 3742 11691 3776
rect 11453 3674 11483 3708
rect 11661 3674 11691 3708
rect 11453 3606 11483 3640
rect 11661 3606 11691 3640
rect 11453 3538 11483 3572
rect 11661 3538 11691 3572
rect 11453 3470 11483 3504
rect 11661 3470 11691 3504
rect 11453 3402 11483 3436
rect 11661 3402 11691 3436
rect 11453 3334 11483 3368
rect 11661 3334 11691 3368
rect 11453 3266 11483 3300
rect 11661 3266 11691 3300
rect 11453 3198 11483 3232
rect 11661 3198 11691 3232
rect 11487 3164 11555 3194
rect 11589 3164 11657 3194
rect 11453 3148 11555 3164
rect 11589 3148 11691 3164
rect 11453 3108 11691 3148
rect 11453 3074 11483 3108
rect 11517 3074 11555 3108
rect 11589 3074 11627 3108
rect 11661 3074 11691 3108
rect 11453 3044 11691 3074
rect 11453 3028 11521 3044
rect 11453 2994 11483 3028
rect 11517 3010 11521 3028
rect 11555 3028 11589 3044
rect 11517 2994 11555 3010
rect 11623 3028 11691 3044
rect 11623 3010 11627 3028
rect 11589 2994 11627 3010
rect 11661 2994 11691 3028
rect 11453 2974 11691 2994
rect 11453 2948 11521 2974
rect 11453 2914 11483 2948
rect 11517 2940 11521 2948
rect 11555 2948 11589 2974
rect 11517 2914 11555 2940
rect 11623 2948 11691 2974
rect 11623 2940 11627 2948
rect 11589 2914 11627 2940
rect 11661 2914 11691 2948
rect 11453 2904 11691 2914
rect 11453 2870 11521 2904
rect 11555 2870 11589 2904
rect 11623 2870 11691 2904
rect 11453 2868 11691 2870
rect 11453 2834 11483 2868
rect 11517 2834 11555 2868
rect 11589 2834 11627 2868
rect 11661 2834 11691 2868
rect 11453 2800 11521 2834
rect 11555 2800 11589 2834
rect 11623 2800 11691 2834
rect 11453 2788 11691 2800
rect 11453 2754 11483 2788
rect 11517 2764 11555 2788
rect 11517 2754 11521 2764
rect 11453 2730 11521 2754
rect 11589 2764 11627 2788
rect 11555 2730 11589 2754
rect 11623 2754 11627 2764
rect 11661 2754 11691 2788
rect 11623 2730 11691 2754
rect 11453 2708 11691 2730
rect 11453 2674 11483 2708
rect 11517 2694 11555 2708
rect 11517 2674 11521 2694
rect 11453 2660 11521 2674
rect 11589 2694 11627 2708
rect 11555 2660 11589 2674
rect 11623 2674 11627 2694
rect 11661 2674 11691 2708
rect 11623 2660 11691 2674
rect 11453 2628 11691 2660
rect 11453 2594 11483 2628
rect 11517 2594 11555 2628
rect 11589 2594 11627 2628
rect 11661 2594 11691 2628
rect 11453 2556 11691 2594
rect 11453 2540 11555 2556
rect 11589 2540 11691 2556
rect 11487 2518 11555 2540
rect 11589 2518 11657 2540
rect 11453 2472 11483 2506
rect 11661 2472 11691 2506
rect 11453 2404 11483 2438
rect 11661 2404 11691 2438
rect 11453 2336 11483 2370
rect 11661 2336 11691 2370
rect 11453 2268 11483 2302
rect 11661 2268 11691 2302
rect 11453 2200 11483 2234
rect 11661 2200 11691 2234
rect 11453 2132 11483 2166
rect 11661 2132 11691 2166
rect 11453 2064 11483 2098
rect 11661 2064 11691 2098
rect 11453 1996 11483 2030
rect 11661 1996 11691 2030
rect 11453 1928 11483 1962
rect 11661 1928 11691 1962
rect 11453 1860 11483 1894
rect 11661 1860 11691 1894
rect 11453 1792 11483 1826
rect 11661 1792 11691 1826
rect 11453 1724 11483 1758
rect 11661 1724 11691 1758
rect 11453 1656 11483 1690
rect 11661 1656 11691 1690
rect 11453 1620 11483 1622
rect 11661 1620 11691 1622
rect 11453 1586 11555 1620
rect 11589 1586 11691 1620
rect 11453 1536 11691 1586
rect 11793 3104 11913 4200
rect 12223 4308 12343 4324
rect 12223 4274 12266 4308
rect 12300 4274 12343 4308
rect 12223 4234 12343 4274
rect 12223 4200 12266 4234
rect 12300 4200 12343 4234
rect 11793 3070 11836 3104
rect 11870 3070 11913 3104
rect 11793 3026 11913 3070
rect 11793 2992 11836 3026
rect 11870 2992 11913 3026
rect 11793 2948 11913 2992
rect 11793 2914 11836 2948
rect 11870 2914 11913 2948
rect 11793 2870 11913 2914
rect 11793 2836 11836 2870
rect 11870 2836 11913 2870
rect 11793 2792 11913 2836
rect 11793 2758 11836 2792
rect 11870 2758 11913 2792
rect 11793 2713 11913 2758
rect 11793 2679 11836 2713
rect 11870 2679 11913 2713
rect 11793 2634 11913 2679
rect 11793 2600 11836 2634
rect 11870 2600 11913 2634
rect 11231 1470 11274 1504
rect 11308 1470 11351 1504
rect 11231 1430 11351 1470
rect 11231 1396 11274 1430
rect 11308 1396 11351 1430
rect 11231 1250 11351 1396
rect 11231 1144 11238 1250
rect 11344 1144 11351 1250
rect 11793 1504 11913 2600
rect 11978 4064 11979 4098
rect 12013 4082 12051 4098
rect 12013 4064 12015 4082
rect 11978 4048 12015 4064
rect 12049 4064 12051 4082
rect 12085 4082 12123 4098
rect 12085 4064 12087 4082
rect 12049 4048 12087 4064
rect 12121 4064 12123 4082
rect 12157 4064 12158 4098
rect 12121 4048 12158 4064
rect 11978 4025 12158 4048
rect 11978 3991 11979 4025
rect 12013 4014 12051 4025
rect 12013 3991 12015 4014
rect 11978 3980 12015 3991
rect 12049 3991 12051 4014
rect 12085 4014 12123 4025
rect 12085 3991 12087 4014
rect 12049 3980 12087 3991
rect 12121 3991 12123 4014
rect 12157 3991 12158 4025
rect 12121 3980 12158 3991
rect 11978 3952 12158 3980
rect 11978 3918 11979 3952
rect 12013 3946 12051 3952
rect 12013 3918 12015 3946
rect 11978 3912 12015 3918
rect 12049 3918 12051 3946
rect 12085 3946 12123 3952
rect 12085 3918 12087 3946
rect 12049 3912 12087 3918
rect 12121 3918 12123 3946
rect 12157 3918 12158 3952
rect 12121 3912 12158 3918
rect 11978 3879 12158 3912
rect 11978 3845 11979 3879
rect 12013 3878 12051 3879
rect 12013 3845 12015 3878
rect 11978 3844 12015 3845
rect 12049 3845 12051 3878
rect 12085 3878 12123 3879
rect 12085 3845 12087 3878
rect 12049 3844 12087 3845
rect 12121 3845 12123 3878
rect 12157 3845 12158 3879
rect 12121 3844 12158 3845
rect 11978 3810 12158 3844
rect 11978 3806 12015 3810
rect 11978 3772 11979 3806
rect 12013 3776 12015 3806
rect 12049 3806 12087 3810
rect 12049 3776 12051 3806
rect 12013 3772 12051 3776
rect 12085 3776 12087 3806
rect 12121 3806 12158 3810
rect 12121 3776 12123 3806
rect 12085 3772 12123 3776
rect 12157 3772 12158 3806
rect 11978 3742 12158 3772
rect 11978 3733 12015 3742
rect 11978 3699 11979 3733
rect 12013 3708 12015 3733
rect 12049 3733 12087 3742
rect 12049 3708 12051 3733
rect 12013 3699 12051 3708
rect 12085 3708 12087 3733
rect 12121 3733 12158 3742
rect 12121 3708 12123 3733
rect 12085 3699 12123 3708
rect 12157 3699 12158 3733
rect 11978 3674 12158 3699
rect 11978 3660 12015 3674
rect 11978 3626 11979 3660
rect 12013 3640 12015 3660
rect 12049 3660 12087 3674
rect 12049 3640 12051 3660
rect 12013 3626 12051 3640
rect 12085 3640 12087 3660
rect 12121 3660 12158 3674
rect 12121 3640 12123 3660
rect 12085 3626 12123 3640
rect 12157 3626 12158 3660
rect 11978 3606 12158 3626
rect 11978 3587 12015 3606
rect 11978 3553 11979 3587
rect 12013 3572 12015 3587
rect 12049 3587 12087 3606
rect 12049 3572 12051 3587
rect 12013 3553 12051 3572
rect 12085 3572 12087 3587
rect 12121 3587 12158 3606
rect 12121 3572 12123 3587
rect 12085 3553 12123 3572
rect 12157 3553 12158 3587
rect 11978 3538 12158 3553
rect 11978 3514 12015 3538
rect 11978 3480 11979 3514
rect 12013 3504 12015 3514
rect 12049 3514 12087 3538
rect 12049 3504 12051 3514
rect 12013 3480 12051 3504
rect 12085 3504 12087 3514
rect 12121 3514 12158 3538
rect 12121 3504 12123 3514
rect 12085 3480 12123 3504
rect 12157 3480 12158 3514
rect 11978 3470 12158 3480
rect 11978 3441 12015 3470
rect 11978 3407 11979 3441
rect 12013 3436 12015 3441
rect 12049 3441 12087 3470
rect 12049 3436 12051 3441
rect 12013 3407 12051 3436
rect 12085 3436 12087 3441
rect 12121 3441 12158 3470
rect 12121 3436 12123 3441
rect 12085 3407 12123 3436
rect 12157 3407 12158 3441
rect 11978 3402 12158 3407
rect 11978 3368 12015 3402
rect 12049 3368 12087 3402
rect 12121 3368 12158 3402
rect 11978 3334 11979 3368
rect 12013 3334 12051 3368
rect 12085 3334 12123 3368
rect 12157 3334 12158 3368
rect 11978 3300 12015 3334
rect 12049 3300 12087 3334
rect 12121 3300 12158 3334
rect 11978 3295 12158 3300
rect 11978 3261 11979 3295
rect 12013 3266 12051 3295
rect 12013 3261 12015 3266
rect 11978 3232 12015 3261
rect 12049 3261 12051 3266
rect 12085 3266 12123 3295
rect 12085 3261 12087 3266
rect 12049 3232 12087 3261
rect 12121 3261 12123 3266
rect 12157 3261 12158 3295
rect 12121 3232 12158 3261
rect 11978 3222 12158 3232
rect 11978 3188 11979 3222
rect 12013 3198 12051 3222
rect 12013 3188 12015 3198
rect 11978 3164 12015 3188
rect 12049 3188 12051 3198
rect 12085 3198 12123 3222
rect 12085 3188 12087 3198
rect 12049 3164 12087 3188
rect 12121 3188 12123 3198
rect 12157 3188 12158 3222
rect 12121 3164 12158 3188
rect 11978 3149 12158 3164
rect 11978 3115 11979 3149
rect 12013 3115 12051 3149
rect 12085 3115 12123 3149
rect 12157 3115 12158 3149
rect 11978 3076 12158 3115
rect 11978 3042 11979 3076
rect 12013 3042 12051 3076
rect 12085 3042 12123 3076
rect 12157 3042 12158 3076
rect 11978 3003 12158 3042
rect 11978 2969 11979 3003
rect 12013 2969 12051 3003
rect 12085 2969 12123 3003
rect 12157 2969 12158 3003
rect 11978 2930 12158 2969
rect 11978 2896 11979 2930
rect 12013 2896 12051 2930
rect 12085 2896 12123 2930
rect 12157 2896 12158 2930
rect 11978 2857 12158 2896
rect 11978 2823 11979 2857
rect 12013 2823 12051 2857
rect 12085 2823 12123 2857
rect 12157 2823 12158 2857
rect 11978 2784 12158 2823
rect 11978 2750 11979 2784
rect 12013 2750 12051 2784
rect 12085 2750 12123 2784
rect 12157 2750 12158 2784
rect 11978 2711 12158 2750
rect 11978 2677 11979 2711
rect 12013 2677 12051 2711
rect 12085 2677 12123 2711
rect 12157 2677 12158 2711
rect 11978 2638 12158 2677
rect 11978 2604 11979 2638
rect 12013 2604 12051 2638
rect 12085 2604 12123 2638
rect 12157 2604 12158 2638
rect 11978 2565 12158 2604
rect 11978 2531 11979 2565
rect 12013 2531 12051 2565
rect 12085 2531 12123 2565
rect 12157 2531 12158 2565
rect 11978 2492 12158 2531
rect 11978 2458 11979 2492
rect 12013 2482 12051 2492
rect 12013 2458 12015 2482
rect 11978 2448 12015 2458
rect 12049 2458 12051 2482
rect 12085 2482 12123 2492
rect 12085 2458 12087 2482
rect 12049 2448 12087 2458
rect 12121 2458 12123 2482
rect 12157 2458 12158 2492
rect 12121 2448 12158 2458
rect 11978 2419 12158 2448
rect 11978 2385 11979 2419
rect 12013 2414 12051 2419
rect 12013 2385 12015 2414
rect 11978 2380 12015 2385
rect 12049 2385 12051 2414
rect 12085 2414 12123 2419
rect 12085 2385 12087 2414
rect 12049 2380 12087 2385
rect 12121 2385 12123 2414
rect 12157 2385 12158 2419
rect 12121 2380 12158 2385
rect 11978 2346 12158 2380
rect 11978 2312 11979 2346
rect 12013 2312 12015 2346
rect 12049 2312 12051 2346
rect 12085 2312 12087 2346
rect 12121 2312 12123 2346
rect 12157 2312 12158 2346
rect 11978 2278 12158 2312
rect 11978 2273 12015 2278
rect 11978 2239 11979 2273
rect 12013 2244 12015 2273
rect 12049 2273 12087 2278
rect 12049 2244 12051 2273
rect 12013 2239 12051 2244
rect 12085 2244 12087 2273
rect 12121 2273 12158 2278
rect 12121 2244 12123 2273
rect 12085 2239 12123 2244
rect 12157 2239 12158 2273
rect 11978 2210 12158 2239
rect 11978 2200 12015 2210
rect 11978 2166 11979 2200
rect 12013 2176 12015 2200
rect 12049 2200 12087 2210
rect 12049 2176 12051 2200
rect 12013 2166 12051 2176
rect 12085 2176 12087 2200
rect 12121 2200 12158 2210
rect 12121 2176 12123 2200
rect 12085 2166 12123 2176
rect 12157 2166 12158 2200
rect 11978 2142 12158 2166
rect 11978 2126 12015 2142
rect 11978 2092 11979 2126
rect 12013 2108 12015 2126
rect 12049 2126 12087 2142
rect 12049 2108 12051 2126
rect 12013 2092 12051 2108
rect 12085 2108 12087 2126
rect 12121 2126 12158 2142
rect 12121 2108 12123 2126
rect 12085 2092 12123 2108
rect 12157 2092 12158 2126
rect 11978 2074 12158 2092
rect 11978 2052 12015 2074
rect 11978 2018 11979 2052
rect 12013 2040 12015 2052
rect 12049 2052 12087 2074
rect 12049 2040 12051 2052
rect 12013 2018 12051 2040
rect 12085 2040 12087 2052
rect 12121 2052 12158 2074
rect 12121 2040 12123 2052
rect 12085 2018 12123 2040
rect 12157 2018 12158 2052
rect 11978 2006 12158 2018
rect 11978 1978 12015 2006
rect 11978 1944 11979 1978
rect 12013 1972 12015 1978
rect 12049 1978 12087 2006
rect 12049 1972 12051 1978
rect 12013 1944 12051 1972
rect 12085 1972 12087 1978
rect 12121 1978 12158 2006
rect 12121 1972 12123 1978
rect 12085 1944 12123 1972
rect 12157 1944 12158 1978
rect 11978 1938 12158 1944
rect 11978 1904 12015 1938
rect 12049 1904 12087 1938
rect 12121 1904 12158 1938
rect 11978 1870 11979 1904
rect 12013 1870 12051 1904
rect 12085 1870 12123 1904
rect 12157 1870 12158 1904
rect 11978 1836 12015 1870
rect 12049 1836 12087 1870
rect 12121 1836 12158 1870
rect 11978 1830 12158 1836
rect 11978 1796 11979 1830
rect 12013 1802 12051 1830
rect 12013 1796 12015 1802
rect 11978 1768 12015 1796
rect 12049 1796 12051 1802
rect 12085 1802 12123 1830
rect 12085 1796 12087 1802
rect 12049 1768 12087 1796
rect 12121 1796 12123 1802
rect 12157 1796 12158 1830
rect 12121 1768 12158 1796
rect 11978 1756 12158 1768
rect 11978 1722 11979 1756
rect 12013 1734 12051 1756
rect 12013 1722 12015 1734
rect 11978 1700 12015 1722
rect 12049 1722 12051 1734
rect 12085 1734 12123 1756
rect 12085 1722 12087 1734
rect 12049 1700 12087 1722
rect 12121 1722 12123 1734
rect 12157 1722 12158 1756
rect 12121 1700 12158 1722
rect 11978 1682 12158 1700
rect 11978 1648 11979 1682
rect 12013 1666 12051 1682
rect 12013 1648 12015 1666
rect 11978 1632 12015 1648
rect 12049 1648 12051 1666
rect 12085 1666 12123 1682
rect 12085 1648 12087 1666
rect 12049 1632 12087 1648
rect 12121 1648 12123 1666
rect 12157 1648 12158 1682
rect 12121 1632 12158 1648
rect 11978 1608 12158 1632
rect 11978 1574 11979 1608
rect 12013 1598 12051 1608
rect 12013 1574 12015 1598
rect 11978 1564 12015 1574
rect 12049 1574 12051 1598
rect 12085 1598 12123 1608
rect 12085 1574 12087 1598
rect 12049 1564 12087 1574
rect 12121 1574 12123 1598
rect 12157 1574 12158 1608
rect 12121 1564 12158 1574
rect 11978 1548 12158 1564
rect 12223 3104 12343 4200
rect 12785 4308 12905 4324
rect 12785 4274 12828 4308
rect 12862 4274 12905 4308
rect 12785 4234 12905 4274
rect 12785 4200 12828 4234
rect 12862 4200 12905 4234
rect 12223 3070 12266 3104
rect 12300 3070 12343 3104
rect 12223 3026 12343 3070
rect 12223 2992 12266 3026
rect 12300 2992 12343 3026
rect 12223 2948 12343 2992
rect 12223 2914 12266 2948
rect 12300 2914 12343 2948
rect 12223 2870 12343 2914
rect 12223 2836 12266 2870
rect 12300 2836 12343 2870
rect 12223 2792 12343 2836
rect 12223 2758 12266 2792
rect 12300 2758 12343 2792
rect 12223 2713 12343 2758
rect 12223 2679 12266 2713
rect 12300 2679 12343 2713
rect 12223 2634 12343 2679
rect 12223 2600 12266 2634
rect 12300 2600 12343 2634
rect 11793 1470 11836 1504
rect 11870 1470 11913 1504
rect 11793 1430 11913 1470
rect 11793 1396 11836 1430
rect 11870 1396 11913 1430
rect 11793 1250 11913 1396
rect 11793 1144 11800 1250
rect 11906 1144 11913 1250
rect 12223 1504 12343 2600
rect 12445 4092 12547 4118
rect 12581 4092 12683 4118
rect 12445 4082 12475 4092
rect 12653 4082 12683 4092
rect 12445 4014 12475 4048
rect 12653 4014 12683 4048
rect 12445 3946 12475 3980
rect 12653 3946 12683 3980
rect 12445 3878 12475 3912
rect 12653 3878 12683 3912
rect 12445 3810 12475 3844
rect 12653 3810 12683 3844
rect 12445 3742 12475 3776
rect 12653 3742 12683 3776
rect 12445 3674 12475 3708
rect 12653 3674 12683 3708
rect 12445 3606 12475 3640
rect 12653 3606 12683 3640
rect 12445 3538 12475 3572
rect 12653 3538 12683 3572
rect 12445 3470 12475 3504
rect 12653 3470 12683 3504
rect 12445 3402 12475 3436
rect 12653 3402 12683 3436
rect 12445 3334 12475 3368
rect 12653 3334 12683 3368
rect 12445 3266 12475 3300
rect 12653 3266 12683 3300
rect 12445 3198 12475 3232
rect 12653 3198 12683 3232
rect 12479 3164 12547 3194
rect 12581 3164 12649 3194
rect 12445 3148 12547 3164
rect 12581 3148 12683 3164
rect 12445 3108 12683 3148
rect 12445 3074 12475 3108
rect 12509 3074 12547 3108
rect 12581 3074 12619 3108
rect 12653 3074 12683 3108
rect 12445 3044 12683 3074
rect 12445 3028 12513 3044
rect 12445 2994 12475 3028
rect 12509 3010 12513 3028
rect 12547 3028 12581 3044
rect 12509 2994 12547 3010
rect 12615 3028 12683 3044
rect 12615 3010 12619 3028
rect 12581 2994 12619 3010
rect 12653 2994 12683 3028
rect 12445 2974 12683 2994
rect 12445 2948 12513 2974
rect 12445 2914 12475 2948
rect 12509 2940 12513 2948
rect 12547 2948 12581 2974
rect 12509 2914 12547 2940
rect 12615 2948 12683 2974
rect 12615 2940 12619 2948
rect 12581 2914 12619 2940
rect 12653 2914 12683 2948
rect 12445 2904 12683 2914
rect 12445 2870 12513 2904
rect 12547 2870 12581 2904
rect 12615 2870 12683 2904
rect 12445 2868 12683 2870
rect 12445 2834 12475 2868
rect 12509 2834 12547 2868
rect 12581 2834 12619 2868
rect 12653 2834 12683 2868
rect 12445 2800 12513 2834
rect 12547 2800 12581 2834
rect 12615 2800 12683 2834
rect 12445 2788 12683 2800
rect 12445 2754 12475 2788
rect 12509 2764 12547 2788
rect 12509 2754 12513 2764
rect 12445 2730 12513 2754
rect 12581 2764 12619 2788
rect 12547 2730 12581 2754
rect 12615 2754 12619 2764
rect 12653 2754 12683 2788
rect 12615 2730 12683 2754
rect 12445 2708 12683 2730
rect 12445 2674 12475 2708
rect 12509 2694 12547 2708
rect 12509 2674 12513 2694
rect 12445 2660 12513 2674
rect 12581 2694 12619 2708
rect 12547 2660 12581 2674
rect 12615 2674 12619 2694
rect 12653 2674 12683 2708
rect 12615 2660 12683 2674
rect 12445 2628 12683 2660
rect 12445 2594 12475 2628
rect 12509 2594 12547 2628
rect 12581 2594 12619 2628
rect 12653 2594 12683 2628
rect 12445 2556 12683 2594
rect 12445 2540 12547 2556
rect 12581 2540 12683 2556
rect 12479 2518 12547 2540
rect 12581 2518 12649 2540
rect 12445 2472 12475 2506
rect 12653 2472 12683 2506
rect 12445 2404 12475 2438
rect 12653 2404 12683 2438
rect 12445 2336 12475 2370
rect 12653 2336 12683 2370
rect 12445 2268 12475 2302
rect 12653 2268 12683 2302
rect 12445 2200 12475 2234
rect 12653 2200 12683 2234
rect 12445 2132 12475 2166
rect 12653 2132 12683 2166
rect 12445 2064 12475 2098
rect 12653 2064 12683 2098
rect 12445 1996 12475 2030
rect 12653 1996 12683 2030
rect 12445 1928 12475 1962
rect 12653 1928 12683 1962
rect 12445 1860 12475 1894
rect 12653 1860 12683 1894
rect 12445 1792 12475 1826
rect 12653 1792 12683 1826
rect 12445 1724 12475 1758
rect 12653 1724 12683 1758
rect 12445 1656 12475 1690
rect 12653 1656 12683 1690
rect 12445 1620 12475 1622
rect 12653 1620 12683 1622
rect 12445 1586 12547 1620
rect 12581 1586 12683 1620
rect 12445 1536 12683 1586
rect 12785 3104 12905 4200
rect 13215 4308 13335 4324
rect 13215 4274 13258 4308
rect 13292 4274 13335 4308
rect 13215 4234 13335 4274
rect 13215 4200 13258 4234
rect 13292 4200 13335 4234
rect 12785 3070 12828 3104
rect 12862 3070 12905 3104
rect 12785 3026 12905 3070
rect 12785 2992 12828 3026
rect 12862 2992 12905 3026
rect 12785 2948 12905 2992
rect 12785 2914 12828 2948
rect 12862 2914 12905 2948
rect 12785 2870 12905 2914
rect 12785 2836 12828 2870
rect 12862 2836 12905 2870
rect 12785 2792 12905 2836
rect 12785 2758 12828 2792
rect 12862 2758 12905 2792
rect 12785 2713 12905 2758
rect 12785 2679 12828 2713
rect 12862 2679 12905 2713
rect 12785 2634 12905 2679
rect 12785 2600 12828 2634
rect 12862 2600 12905 2634
rect 12223 1470 12266 1504
rect 12300 1470 12343 1504
rect 12223 1430 12343 1470
rect 12223 1396 12266 1430
rect 12300 1396 12343 1430
rect 12223 1250 12343 1396
rect 12223 1144 12230 1250
rect 12336 1144 12343 1250
rect 12785 1504 12905 2600
rect 12970 4064 12971 4098
rect 13005 4082 13043 4098
rect 13005 4064 13007 4082
rect 12970 4048 13007 4064
rect 13041 4064 13043 4082
rect 13077 4082 13115 4098
rect 13077 4064 13079 4082
rect 13041 4048 13079 4064
rect 13113 4064 13115 4082
rect 13149 4064 13150 4098
rect 13113 4048 13150 4064
rect 12970 4025 13150 4048
rect 12970 3991 12971 4025
rect 13005 4014 13043 4025
rect 13005 3991 13007 4014
rect 12970 3980 13007 3991
rect 13041 3991 13043 4014
rect 13077 4014 13115 4025
rect 13077 3991 13079 4014
rect 13041 3980 13079 3991
rect 13113 3991 13115 4014
rect 13149 3991 13150 4025
rect 13113 3980 13150 3991
rect 12970 3952 13150 3980
rect 12970 3918 12971 3952
rect 13005 3946 13043 3952
rect 13005 3918 13007 3946
rect 12970 3912 13007 3918
rect 13041 3918 13043 3946
rect 13077 3946 13115 3952
rect 13077 3918 13079 3946
rect 13041 3912 13079 3918
rect 13113 3918 13115 3946
rect 13149 3918 13150 3952
rect 13113 3912 13150 3918
rect 12970 3879 13150 3912
rect 12970 3845 12971 3879
rect 13005 3878 13043 3879
rect 13005 3845 13007 3878
rect 12970 3844 13007 3845
rect 13041 3845 13043 3878
rect 13077 3878 13115 3879
rect 13077 3845 13079 3878
rect 13041 3844 13079 3845
rect 13113 3845 13115 3878
rect 13149 3845 13150 3879
rect 13113 3844 13150 3845
rect 12970 3810 13150 3844
rect 12970 3806 13007 3810
rect 12970 3772 12971 3806
rect 13005 3776 13007 3806
rect 13041 3806 13079 3810
rect 13041 3776 13043 3806
rect 13005 3772 13043 3776
rect 13077 3776 13079 3806
rect 13113 3806 13150 3810
rect 13113 3776 13115 3806
rect 13077 3772 13115 3776
rect 13149 3772 13150 3806
rect 12970 3742 13150 3772
rect 12970 3733 13007 3742
rect 12970 3699 12971 3733
rect 13005 3708 13007 3733
rect 13041 3733 13079 3742
rect 13041 3708 13043 3733
rect 13005 3699 13043 3708
rect 13077 3708 13079 3733
rect 13113 3733 13150 3742
rect 13113 3708 13115 3733
rect 13077 3699 13115 3708
rect 13149 3699 13150 3733
rect 12970 3674 13150 3699
rect 12970 3660 13007 3674
rect 12970 3626 12971 3660
rect 13005 3640 13007 3660
rect 13041 3660 13079 3674
rect 13041 3640 13043 3660
rect 13005 3626 13043 3640
rect 13077 3640 13079 3660
rect 13113 3660 13150 3674
rect 13113 3640 13115 3660
rect 13077 3626 13115 3640
rect 13149 3626 13150 3660
rect 12970 3606 13150 3626
rect 12970 3587 13007 3606
rect 12970 3553 12971 3587
rect 13005 3572 13007 3587
rect 13041 3587 13079 3606
rect 13041 3572 13043 3587
rect 13005 3553 13043 3572
rect 13077 3572 13079 3587
rect 13113 3587 13150 3606
rect 13113 3572 13115 3587
rect 13077 3553 13115 3572
rect 13149 3553 13150 3587
rect 12970 3538 13150 3553
rect 12970 3514 13007 3538
rect 12970 3480 12971 3514
rect 13005 3504 13007 3514
rect 13041 3514 13079 3538
rect 13041 3504 13043 3514
rect 13005 3480 13043 3504
rect 13077 3504 13079 3514
rect 13113 3514 13150 3538
rect 13113 3504 13115 3514
rect 13077 3480 13115 3504
rect 13149 3480 13150 3514
rect 12970 3470 13150 3480
rect 12970 3441 13007 3470
rect 12970 3407 12971 3441
rect 13005 3436 13007 3441
rect 13041 3441 13079 3470
rect 13041 3436 13043 3441
rect 13005 3407 13043 3436
rect 13077 3436 13079 3441
rect 13113 3441 13150 3470
rect 13113 3436 13115 3441
rect 13077 3407 13115 3436
rect 13149 3407 13150 3441
rect 12970 3402 13150 3407
rect 12970 3368 13007 3402
rect 13041 3368 13079 3402
rect 13113 3368 13150 3402
rect 12970 3334 12971 3368
rect 13005 3334 13043 3368
rect 13077 3334 13115 3368
rect 13149 3334 13150 3368
rect 12970 3300 13007 3334
rect 13041 3300 13079 3334
rect 13113 3300 13150 3334
rect 12970 3295 13150 3300
rect 12970 3261 12971 3295
rect 13005 3266 13043 3295
rect 13005 3261 13007 3266
rect 12970 3232 13007 3261
rect 13041 3261 13043 3266
rect 13077 3266 13115 3295
rect 13077 3261 13079 3266
rect 13041 3232 13079 3261
rect 13113 3261 13115 3266
rect 13149 3261 13150 3295
rect 13113 3232 13150 3261
rect 12970 3222 13150 3232
rect 12970 3188 12971 3222
rect 13005 3198 13043 3222
rect 13005 3188 13007 3198
rect 12970 3164 13007 3188
rect 13041 3188 13043 3198
rect 13077 3198 13115 3222
rect 13077 3188 13079 3198
rect 13041 3164 13079 3188
rect 13113 3188 13115 3198
rect 13149 3188 13150 3222
rect 13113 3164 13150 3188
rect 12970 3149 13150 3164
rect 12970 3115 12971 3149
rect 13005 3115 13043 3149
rect 13077 3115 13115 3149
rect 13149 3115 13150 3149
rect 12970 3076 13150 3115
rect 12970 3042 12971 3076
rect 13005 3042 13043 3076
rect 13077 3042 13115 3076
rect 13149 3042 13150 3076
rect 12970 3003 13150 3042
rect 12970 2969 12971 3003
rect 13005 2969 13043 3003
rect 13077 2969 13115 3003
rect 13149 2969 13150 3003
rect 12970 2930 13150 2969
rect 12970 2896 12971 2930
rect 13005 2896 13043 2930
rect 13077 2896 13115 2930
rect 13149 2896 13150 2930
rect 12970 2857 13150 2896
rect 12970 2823 12971 2857
rect 13005 2823 13043 2857
rect 13077 2823 13115 2857
rect 13149 2823 13150 2857
rect 12970 2784 13150 2823
rect 12970 2750 12971 2784
rect 13005 2750 13043 2784
rect 13077 2750 13115 2784
rect 13149 2750 13150 2784
rect 12970 2711 13150 2750
rect 12970 2677 12971 2711
rect 13005 2677 13043 2711
rect 13077 2677 13115 2711
rect 13149 2677 13150 2711
rect 12970 2638 13150 2677
rect 12970 2604 12971 2638
rect 13005 2604 13043 2638
rect 13077 2604 13115 2638
rect 13149 2604 13150 2638
rect 12970 2565 13150 2604
rect 12970 2531 12971 2565
rect 13005 2531 13043 2565
rect 13077 2531 13115 2565
rect 13149 2531 13150 2565
rect 12970 2492 13150 2531
rect 12970 2458 12971 2492
rect 13005 2482 13043 2492
rect 13005 2458 13007 2482
rect 12970 2448 13007 2458
rect 13041 2458 13043 2482
rect 13077 2482 13115 2492
rect 13077 2458 13079 2482
rect 13041 2448 13079 2458
rect 13113 2458 13115 2482
rect 13149 2458 13150 2492
rect 13113 2448 13150 2458
rect 12970 2419 13150 2448
rect 12970 2385 12971 2419
rect 13005 2414 13043 2419
rect 13005 2385 13007 2414
rect 12970 2380 13007 2385
rect 13041 2385 13043 2414
rect 13077 2414 13115 2419
rect 13077 2385 13079 2414
rect 13041 2380 13079 2385
rect 13113 2385 13115 2414
rect 13149 2385 13150 2419
rect 13113 2380 13150 2385
rect 12970 2346 13150 2380
rect 12970 2312 12971 2346
rect 13005 2312 13007 2346
rect 13041 2312 13043 2346
rect 13077 2312 13079 2346
rect 13113 2312 13115 2346
rect 13149 2312 13150 2346
rect 12970 2278 13150 2312
rect 12970 2273 13007 2278
rect 12970 2239 12971 2273
rect 13005 2244 13007 2273
rect 13041 2273 13079 2278
rect 13041 2244 13043 2273
rect 13005 2239 13043 2244
rect 13077 2244 13079 2273
rect 13113 2273 13150 2278
rect 13113 2244 13115 2273
rect 13077 2239 13115 2244
rect 13149 2239 13150 2273
rect 12970 2210 13150 2239
rect 12970 2200 13007 2210
rect 12970 2166 12971 2200
rect 13005 2176 13007 2200
rect 13041 2200 13079 2210
rect 13041 2176 13043 2200
rect 13005 2166 13043 2176
rect 13077 2176 13079 2200
rect 13113 2200 13150 2210
rect 13113 2176 13115 2200
rect 13077 2166 13115 2176
rect 13149 2166 13150 2200
rect 12970 2142 13150 2166
rect 12970 2126 13007 2142
rect 12970 2092 12971 2126
rect 13005 2108 13007 2126
rect 13041 2126 13079 2142
rect 13041 2108 13043 2126
rect 13005 2092 13043 2108
rect 13077 2108 13079 2126
rect 13113 2126 13150 2142
rect 13113 2108 13115 2126
rect 13077 2092 13115 2108
rect 13149 2092 13150 2126
rect 12970 2074 13150 2092
rect 12970 2052 13007 2074
rect 12970 2018 12971 2052
rect 13005 2040 13007 2052
rect 13041 2052 13079 2074
rect 13041 2040 13043 2052
rect 13005 2018 13043 2040
rect 13077 2040 13079 2052
rect 13113 2052 13150 2074
rect 13113 2040 13115 2052
rect 13077 2018 13115 2040
rect 13149 2018 13150 2052
rect 12970 2006 13150 2018
rect 12970 1978 13007 2006
rect 12970 1944 12971 1978
rect 13005 1972 13007 1978
rect 13041 1978 13079 2006
rect 13041 1972 13043 1978
rect 13005 1944 13043 1972
rect 13077 1972 13079 1978
rect 13113 1978 13150 2006
rect 13113 1972 13115 1978
rect 13077 1944 13115 1972
rect 13149 1944 13150 1978
rect 12970 1938 13150 1944
rect 12970 1904 13007 1938
rect 13041 1904 13079 1938
rect 13113 1904 13150 1938
rect 12970 1870 12971 1904
rect 13005 1870 13043 1904
rect 13077 1870 13115 1904
rect 13149 1870 13150 1904
rect 12970 1836 13007 1870
rect 13041 1836 13079 1870
rect 13113 1836 13150 1870
rect 12970 1830 13150 1836
rect 12970 1796 12971 1830
rect 13005 1802 13043 1830
rect 13005 1796 13007 1802
rect 12970 1768 13007 1796
rect 13041 1796 13043 1802
rect 13077 1802 13115 1830
rect 13077 1796 13079 1802
rect 13041 1768 13079 1796
rect 13113 1796 13115 1802
rect 13149 1796 13150 1830
rect 13113 1768 13150 1796
rect 12970 1756 13150 1768
rect 12970 1722 12971 1756
rect 13005 1734 13043 1756
rect 13005 1722 13007 1734
rect 12970 1700 13007 1722
rect 13041 1722 13043 1734
rect 13077 1734 13115 1756
rect 13077 1722 13079 1734
rect 13041 1700 13079 1722
rect 13113 1722 13115 1734
rect 13149 1722 13150 1756
rect 13113 1700 13150 1722
rect 12970 1682 13150 1700
rect 12970 1648 12971 1682
rect 13005 1666 13043 1682
rect 13005 1648 13007 1666
rect 12970 1632 13007 1648
rect 13041 1648 13043 1666
rect 13077 1666 13115 1682
rect 13077 1648 13079 1666
rect 13041 1632 13079 1648
rect 13113 1648 13115 1666
rect 13149 1648 13150 1682
rect 13113 1632 13150 1648
rect 12970 1608 13150 1632
rect 12970 1574 12971 1608
rect 13005 1598 13043 1608
rect 13005 1574 13007 1598
rect 12970 1564 13007 1574
rect 13041 1574 13043 1598
rect 13077 1598 13115 1608
rect 13077 1574 13079 1598
rect 13041 1564 13079 1574
rect 13113 1574 13115 1598
rect 13149 1574 13150 1608
rect 13113 1564 13150 1574
rect 12970 1548 13150 1564
rect 13215 3104 13335 4200
rect 13777 4308 13897 4324
rect 13777 4274 13820 4308
rect 13854 4274 13897 4308
rect 13777 4234 13897 4274
rect 13777 4200 13820 4234
rect 13854 4200 13897 4234
rect 13215 3070 13258 3104
rect 13292 3070 13335 3104
rect 13215 3026 13335 3070
rect 13215 2992 13258 3026
rect 13292 2992 13335 3026
rect 13215 2948 13335 2992
rect 13215 2914 13258 2948
rect 13292 2914 13335 2948
rect 13215 2870 13335 2914
rect 13215 2836 13258 2870
rect 13292 2836 13335 2870
rect 13215 2792 13335 2836
rect 13215 2758 13258 2792
rect 13292 2758 13335 2792
rect 13215 2713 13335 2758
rect 13215 2679 13258 2713
rect 13292 2679 13335 2713
rect 13215 2634 13335 2679
rect 13215 2600 13258 2634
rect 13292 2600 13335 2634
rect 12785 1470 12828 1504
rect 12862 1470 12905 1504
rect 12785 1430 12905 1470
rect 12785 1396 12828 1430
rect 12862 1396 12905 1430
rect 12785 1250 12905 1396
rect 12785 1144 12792 1250
rect 12898 1144 12905 1250
rect 13215 1504 13335 2600
rect 13437 4092 13539 4118
rect 13573 4092 13675 4118
rect 13437 4082 13467 4092
rect 13645 4082 13675 4092
rect 13437 4014 13467 4048
rect 13645 4014 13675 4048
rect 13437 3946 13467 3980
rect 13645 3946 13675 3980
rect 13437 3878 13467 3912
rect 13645 3878 13675 3912
rect 13437 3810 13467 3844
rect 13645 3810 13675 3844
rect 13437 3742 13467 3776
rect 13645 3742 13675 3776
rect 13437 3674 13467 3708
rect 13645 3674 13675 3708
rect 13437 3606 13467 3640
rect 13645 3606 13675 3640
rect 13437 3538 13467 3572
rect 13645 3538 13675 3572
rect 13437 3470 13467 3504
rect 13645 3470 13675 3504
rect 13437 3402 13467 3436
rect 13645 3402 13675 3436
rect 13437 3334 13467 3368
rect 13645 3334 13675 3368
rect 13437 3266 13467 3300
rect 13645 3266 13675 3300
rect 13437 3198 13467 3232
rect 13645 3198 13675 3232
rect 13471 3164 13539 3194
rect 13573 3164 13641 3194
rect 13437 3148 13539 3164
rect 13573 3148 13675 3164
rect 13437 3108 13675 3148
rect 13437 3074 13467 3108
rect 13501 3074 13539 3108
rect 13573 3074 13611 3108
rect 13645 3074 13675 3108
rect 13437 3044 13675 3074
rect 13437 3028 13505 3044
rect 13437 2994 13467 3028
rect 13501 3010 13505 3028
rect 13539 3028 13573 3044
rect 13501 2994 13539 3010
rect 13607 3028 13675 3044
rect 13607 3010 13611 3028
rect 13573 2994 13611 3010
rect 13645 2994 13675 3028
rect 13437 2974 13675 2994
rect 13437 2948 13505 2974
rect 13437 2914 13467 2948
rect 13501 2940 13505 2948
rect 13539 2948 13573 2974
rect 13501 2914 13539 2940
rect 13607 2948 13675 2974
rect 13607 2940 13611 2948
rect 13573 2914 13611 2940
rect 13645 2914 13675 2948
rect 13437 2904 13675 2914
rect 13437 2870 13505 2904
rect 13539 2870 13573 2904
rect 13607 2870 13675 2904
rect 13437 2868 13675 2870
rect 13437 2834 13467 2868
rect 13501 2834 13539 2868
rect 13573 2834 13611 2868
rect 13645 2834 13675 2868
rect 13437 2800 13505 2834
rect 13539 2800 13573 2834
rect 13607 2800 13675 2834
rect 13437 2788 13675 2800
rect 13437 2754 13467 2788
rect 13501 2764 13539 2788
rect 13501 2754 13505 2764
rect 13437 2730 13505 2754
rect 13573 2764 13611 2788
rect 13539 2730 13573 2754
rect 13607 2754 13611 2764
rect 13645 2754 13675 2788
rect 13607 2730 13675 2754
rect 13437 2708 13675 2730
rect 13437 2674 13467 2708
rect 13501 2694 13539 2708
rect 13501 2674 13505 2694
rect 13437 2660 13505 2674
rect 13573 2694 13611 2708
rect 13539 2660 13573 2674
rect 13607 2674 13611 2694
rect 13645 2674 13675 2708
rect 13607 2660 13675 2674
rect 13437 2628 13675 2660
rect 13437 2594 13467 2628
rect 13501 2594 13539 2628
rect 13573 2594 13611 2628
rect 13645 2594 13675 2628
rect 13437 2556 13675 2594
rect 13437 2540 13539 2556
rect 13573 2540 13675 2556
rect 13471 2518 13539 2540
rect 13573 2518 13641 2540
rect 13437 2472 13467 2506
rect 13645 2472 13675 2506
rect 13437 2404 13467 2438
rect 13645 2404 13675 2438
rect 13437 2336 13467 2370
rect 13645 2336 13675 2370
rect 13437 2268 13467 2302
rect 13645 2268 13675 2302
rect 13437 2200 13467 2234
rect 13645 2200 13675 2234
rect 13437 2132 13467 2166
rect 13645 2132 13675 2166
rect 13437 2064 13467 2098
rect 13645 2064 13675 2098
rect 13437 1996 13467 2030
rect 13645 1996 13675 2030
rect 13437 1928 13467 1962
rect 13645 1928 13675 1962
rect 13437 1860 13467 1894
rect 13645 1860 13675 1894
rect 13437 1792 13467 1826
rect 13645 1792 13675 1826
rect 13437 1724 13467 1758
rect 13645 1724 13675 1758
rect 13437 1656 13467 1690
rect 13645 1656 13675 1690
rect 13437 1620 13467 1622
rect 13645 1620 13675 1622
rect 13437 1586 13539 1620
rect 13573 1586 13675 1620
rect 13437 1536 13675 1586
rect 13777 3104 13897 4200
rect 14135 4308 14255 4324
rect 14135 4274 14178 4308
rect 14212 4274 14255 4308
rect 14135 4234 14255 4274
rect 14135 4200 14178 4234
rect 14212 4200 14255 4234
rect 13777 3070 13820 3104
rect 13854 3070 13897 3104
rect 13777 3026 13897 3070
rect 13777 2992 13820 3026
rect 13854 2992 13897 3026
rect 13777 2948 13897 2992
rect 13777 2914 13820 2948
rect 13854 2914 13897 2948
rect 13777 2870 13897 2914
rect 13777 2836 13820 2870
rect 13854 2836 13897 2870
rect 13777 2792 13897 2836
rect 13777 2758 13820 2792
rect 13854 2758 13897 2792
rect 13777 2713 13897 2758
rect 13777 2679 13820 2713
rect 13854 2679 13897 2713
rect 13777 2634 13897 2679
rect 13777 2600 13820 2634
rect 13854 2600 13897 2634
rect 13215 1470 13258 1504
rect 13292 1470 13335 1504
rect 13215 1430 13335 1470
rect 13215 1396 13258 1430
rect 13292 1396 13335 1430
rect 13215 1250 13335 1396
rect 13215 1144 13222 1250
rect 13328 1144 13335 1250
rect 13777 1504 13897 2600
rect 13997 4082 14035 4098
rect 13997 4064 13999 4082
rect 13963 4048 13999 4064
rect 14033 4064 14035 4082
rect 14033 4048 14069 4064
rect 13963 4024 14069 4048
rect 13997 4014 14035 4024
rect 13997 3990 13999 4014
rect 13963 3980 13999 3990
rect 14033 3990 14035 4014
rect 14033 3980 14069 3990
rect 13963 3950 14069 3980
rect 13997 3946 14035 3950
rect 13997 3916 13999 3946
rect 13963 3912 13999 3916
rect 14033 3916 14035 3946
rect 14033 3912 14069 3916
rect 13963 3878 14069 3912
rect 13963 3876 13999 3878
rect 13997 3844 13999 3876
rect 14033 3876 14069 3878
rect 14033 3844 14035 3876
rect 13997 3842 14035 3844
rect 13963 3810 14069 3842
rect 13963 3802 13999 3810
rect 13997 3776 13999 3802
rect 14033 3802 14069 3810
rect 14033 3776 14035 3802
rect 13997 3768 14035 3776
rect 13963 3742 14069 3768
rect 13963 3728 13999 3742
rect 13997 3708 13999 3728
rect 14033 3728 14069 3742
rect 14033 3708 14035 3728
rect 13997 3694 14035 3708
rect 13963 3674 14069 3694
rect 13963 3654 13999 3674
rect 13997 3640 13999 3654
rect 14033 3654 14069 3674
rect 14033 3640 14035 3654
rect 13997 3620 14035 3640
rect 13963 3606 14069 3620
rect 13963 3580 13999 3606
rect 13997 3572 13999 3580
rect 14033 3580 14069 3606
rect 14033 3572 14035 3580
rect 13997 3546 14035 3572
rect 13963 3538 14069 3546
rect 13963 3506 13999 3538
rect 13997 3504 13999 3506
rect 14033 3506 14069 3538
rect 14033 3504 14035 3506
rect 13997 3472 14035 3504
rect 13963 3470 14069 3472
rect 13963 3436 13999 3470
rect 14033 3436 14069 3470
rect 13963 3432 14069 3436
rect 13997 3402 14035 3432
rect 13997 3398 13999 3402
rect 13963 3368 13999 3398
rect 14033 3398 14035 3402
rect 14033 3368 14069 3398
rect 13963 3358 14069 3368
rect 13997 3334 14035 3358
rect 13997 3324 13999 3334
rect 13963 3300 13999 3324
rect 14033 3324 14035 3334
rect 14033 3300 14069 3324
rect 13963 3284 14069 3300
rect 13997 3266 14035 3284
rect 13997 3250 13999 3266
rect 13963 3232 13999 3250
rect 14033 3250 14035 3266
rect 14033 3232 14069 3250
rect 13963 3210 14069 3232
rect 13997 3198 14035 3210
rect 13997 3176 13999 3198
rect 13963 3164 13999 3176
rect 14033 3176 14035 3198
rect 14033 3164 14069 3176
rect 13963 3136 14069 3164
rect 13997 3102 14035 3136
rect 13963 3062 14069 3102
rect 13997 3028 14035 3062
rect 13963 2988 14069 3028
rect 13997 2954 14035 2988
rect 13963 2914 14069 2954
rect 13997 2880 14035 2914
rect 13963 2840 14069 2880
rect 13997 2806 14035 2840
rect 13963 2766 14069 2806
rect 13997 2732 14035 2766
rect 13963 2692 14069 2732
rect 13997 2658 14035 2692
rect 13963 2618 14069 2658
rect 13997 2584 14035 2618
rect 13963 2544 14069 2584
rect 13997 2510 14035 2544
rect 13963 2482 14069 2510
rect 13963 2470 13999 2482
rect 13997 2448 13999 2470
rect 14033 2470 14069 2482
rect 14033 2448 14035 2470
rect 13997 2436 14035 2448
rect 13963 2414 14069 2436
rect 13963 2396 13999 2414
rect 13997 2380 13999 2396
rect 14033 2396 14069 2414
rect 14033 2380 14035 2396
rect 13997 2362 14035 2380
rect 13963 2346 14069 2362
rect 13963 2322 13999 2346
rect 13997 2312 13999 2322
rect 14033 2322 14069 2346
rect 14033 2312 14035 2322
rect 13997 2288 14035 2312
rect 13963 2278 14069 2288
rect 13963 2248 13999 2278
rect 13997 2244 13999 2248
rect 14033 2248 14069 2278
rect 14033 2244 14035 2248
rect 13997 2214 14035 2244
rect 13963 2210 14069 2214
rect 13963 2176 13999 2210
rect 14033 2176 14069 2210
rect 13963 2174 14069 2176
rect 13997 2142 14035 2174
rect 13997 2140 13999 2142
rect 13963 2108 13999 2140
rect 14033 2140 14035 2142
rect 14033 2108 14069 2140
rect 13963 2100 14069 2108
rect 13997 2074 14035 2100
rect 13997 2066 13999 2074
rect 13963 2040 13999 2066
rect 14033 2066 14035 2074
rect 14033 2040 14069 2066
rect 13963 2026 14069 2040
rect 13997 2006 14035 2026
rect 13997 1992 13999 2006
rect 13963 1972 13999 1992
rect 14033 1992 14035 2006
rect 14033 1972 14069 1992
rect 13963 1952 14069 1972
rect 13997 1938 14035 1952
rect 13997 1918 13999 1938
rect 13963 1904 13999 1918
rect 14033 1918 14035 1938
rect 14033 1904 14069 1918
rect 13963 1878 14069 1904
rect 13997 1870 14035 1878
rect 13997 1844 13999 1870
rect 13963 1836 13999 1844
rect 14033 1844 14035 1870
rect 14033 1836 14069 1844
rect 13963 1804 14069 1836
rect 13997 1802 14035 1804
rect 13997 1770 13999 1802
rect 13963 1768 13999 1770
rect 14033 1770 14035 1802
rect 14033 1768 14069 1770
rect 13963 1734 14069 1768
rect 13963 1730 13999 1734
rect 13997 1700 13999 1730
rect 14033 1730 14069 1734
rect 14033 1700 14035 1730
rect 13997 1696 14035 1700
rect 13963 1666 14069 1696
rect 13963 1656 13999 1666
rect 13997 1632 13999 1656
rect 14033 1656 14069 1666
rect 14033 1632 14035 1656
rect 13997 1622 14035 1632
rect 13963 1598 14069 1622
rect 13963 1582 13999 1598
rect 13997 1564 13999 1582
rect 14033 1582 14069 1598
rect 14033 1564 14035 1582
rect 13997 1548 14035 1564
rect 14135 3104 14255 4200
rect 14135 3070 14178 3104
rect 14212 3070 14255 3104
rect 14135 3026 14255 3070
rect 14135 2992 14178 3026
rect 14212 2992 14255 3026
rect 14135 2948 14255 2992
rect 14135 2914 14178 2948
rect 14212 2914 14255 2948
rect 14135 2870 14255 2914
rect 14135 2836 14178 2870
rect 14212 2836 14255 2870
rect 14135 2792 14255 2836
rect 14135 2758 14178 2792
rect 14212 2758 14255 2792
rect 14135 2713 14255 2758
rect 14135 2679 14178 2713
rect 14212 2679 14255 2713
rect 14135 2634 14255 2679
rect 14135 2600 14178 2634
rect 14212 2600 14255 2634
rect 13777 1470 13820 1504
rect 13854 1470 13897 1504
rect 13777 1430 13897 1470
rect 13777 1396 13820 1430
rect 13854 1396 13897 1430
rect 13777 1250 13897 1396
rect 13777 1144 13784 1250
rect 13890 1144 13897 1250
rect 14135 1504 14255 2600
rect 14135 1470 14178 1504
rect 14212 1470 14255 1504
rect 14135 1430 14255 1470
rect 14135 1396 14178 1430
rect 14212 1396 14255 1430
rect 14135 1250 14255 1396
rect 14135 1144 14142 1250
rect 14248 1144 14255 1250
rect 14356 4286 14428 4325
rect 14390 4252 14428 4286
rect 14356 4213 14428 4252
rect 14390 4179 14428 4213
rect 14356 4140 14428 4179
rect 14390 4106 14428 4140
rect 14356 4082 14428 4106
rect 14390 4033 14428 4082
rect 14356 4014 14428 4033
rect 14390 3960 14428 4014
rect 14356 3957 14536 3960
rect 14356 3952 14468 3957
rect 14356 3946 14428 3952
rect 14390 3918 14428 3946
rect 14462 3923 14468 3952
rect 14502 3924 14536 3957
rect 14502 3923 14604 3924
rect 14462 3921 14604 3923
rect 14462 3918 14500 3921
rect 14390 3888 14500 3918
rect 14534 3889 14572 3921
rect 14638 3905 14653 4551
rect 14390 3887 14468 3888
rect 14534 3887 14536 3889
rect 14356 3880 14468 3887
rect 14356 3878 14428 3880
rect 14390 3846 14428 3878
rect 14462 3854 14468 3880
rect 14502 3855 14536 3887
rect 14570 3887 14572 3889
rect 14606 3887 14653 3905
rect 14570 3871 14653 3887
rect 14570 3855 14604 3871
rect 14502 3854 14604 3855
rect 14462 3848 14604 3854
rect 14462 3846 14500 3848
rect 14390 3819 14500 3846
rect 14534 3820 14572 3848
rect 14638 3837 14653 3871
rect 14390 3814 14468 3819
rect 14534 3814 14536 3820
rect 14356 3810 14468 3814
rect 14390 3808 14468 3810
rect 14390 3776 14428 3808
rect 14356 3775 14428 3776
rect 14390 3774 14428 3775
rect 14462 3785 14468 3808
rect 14502 3786 14536 3814
rect 14570 3814 14572 3820
rect 14606 3814 14653 3837
rect 14570 3803 14653 3814
rect 14570 3786 14604 3803
rect 14502 3785 14604 3786
rect 14462 3775 14604 3785
rect 14462 3774 14500 3775
rect 14390 3750 14500 3774
rect 14534 3751 14572 3775
rect 14638 3769 14653 3803
rect 14390 3736 14468 3750
rect 14534 3741 14536 3751
rect 14390 3708 14428 3736
rect 14356 3702 14428 3708
rect 14462 3716 14468 3736
rect 14502 3717 14536 3741
rect 14570 3741 14572 3751
rect 14606 3741 14653 3769
rect 14570 3735 14653 3741
rect 14570 3717 14604 3735
rect 14502 3716 14604 3717
rect 14462 3702 14604 3716
rect 14390 3681 14500 3702
rect 14534 3682 14572 3702
rect 14638 3701 14653 3735
rect 14390 3664 14468 3681
rect 14534 3668 14536 3682
rect 14390 3640 14428 3664
rect 14356 3630 14428 3640
rect 14462 3647 14468 3664
rect 14502 3648 14536 3668
rect 14570 3668 14572 3682
rect 14606 3668 14653 3701
rect 14570 3667 14653 3668
rect 14570 3648 14604 3667
rect 14502 3647 14604 3648
rect 14462 3633 14604 3647
rect 14638 3633 14653 3667
rect 14462 3630 14653 3633
rect 14356 3629 14653 3630
rect 14390 3612 14500 3629
rect 14534 3613 14572 3629
rect 14390 3592 14468 3612
rect 14534 3595 14536 3613
rect 14390 3572 14428 3592
rect 14356 3558 14428 3572
rect 14462 3578 14468 3592
rect 14502 3579 14536 3595
rect 14570 3595 14572 3613
rect 14606 3599 14653 3629
rect 14570 3579 14604 3595
rect 14502 3578 14604 3579
rect 14462 3565 14604 3578
rect 14638 3565 14653 3599
rect 14462 3558 14653 3565
rect 14356 3556 14653 3558
rect 14390 3543 14500 3556
rect 14534 3544 14572 3556
rect 14390 3520 14468 3543
rect 14534 3522 14536 3544
rect 14390 3504 14428 3520
rect 14356 3486 14428 3504
rect 14462 3509 14468 3520
rect 14502 3510 14536 3522
rect 14570 3522 14572 3544
rect 14606 3531 14653 3556
rect 14570 3510 14604 3522
rect 14502 3509 14604 3510
rect 14462 3497 14604 3509
rect 14638 3497 14653 3531
rect 14462 3486 14653 3497
rect 14356 3483 14653 3486
rect 14390 3474 14500 3483
rect 14534 3475 14572 3483
rect 14390 3448 14468 3474
rect 14534 3449 14536 3475
rect 14390 3436 14428 3448
rect 14356 3414 14428 3436
rect 14462 3440 14468 3448
rect 14502 3441 14536 3449
rect 14570 3449 14572 3475
rect 14606 3463 14653 3483
rect 14570 3441 14604 3449
rect 14502 3440 14604 3441
rect 14462 3429 14604 3440
rect 14638 3429 14653 3463
rect 14462 3414 14653 3429
rect 14356 3410 14653 3414
rect 14390 3405 14500 3410
rect 14534 3406 14572 3410
rect 14390 3376 14468 3405
rect 14534 3376 14536 3406
rect 14390 3368 14428 3376
rect 14356 3342 14428 3368
rect 14462 3371 14468 3376
rect 14502 3372 14536 3376
rect 14570 3376 14572 3406
rect 14606 3395 14653 3410
rect 14570 3372 14604 3376
rect 14502 3371 14604 3372
rect 14462 3361 14604 3371
rect 14638 3361 14653 3395
rect 14462 3342 14653 3361
rect 14356 3337 14653 3342
rect 14390 3336 14500 3337
rect 14390 3304 14468 3336
rect 14390 3300 14428 3304
rect 14356 3270 14428 3300
rect 14462 3302 14468 3304
rect 14534 3303 14536 3337
rect 14570 3303 14572 3337
rect 14606 3327 14653 3337
rect 14502 3302 14604 3303
rect 14462 3293 14604 3302
rect 14638 3293 14653 3327
rect 14462 3270 14653 3293
rect 14356 3268 14653 3270
rect 14356 3267 14536 3268
rect 14356 3266 14468 3267
rect 14390 3233 14468 3266
rect 14502 3264 14536 3267
rect 14534 3234 14536 3264
rect 14570 3264 14653 3268
rect 14570 3234 14572 3264
rect 14606 3259 14653 3264
rect 14390 3232 14500 3233
rect 14390 3230 14428 3232
rect 14356 3198 14428 3230
rect 14462 3230 14500 3232
rect 14534 3230 14572 3234
rect 14462 3225 14604 3230
rect 14638 3225 14653 3259
rect 14462 3199 14653 3225
rect 14462 3198 14536 3199
rect 14390 3164 14468 3198
rect 14502 3191 14536 3198
rect 14534 3165 14536 3191
rect 14570 3191 14653 3199
rect 14570 3165 14572 3191
rect 14390 3160 14500 3164
rect 14390 3157 14428 3160
rect 14356 3126 14428 3157
rect 14462 3157 14500 3160
rect 14534 3157 14572 3165
rect 14638 3157 14653 3191
rect 14462 3130 14653 3157
rect 14462 3129 14536 3130
rect 14462 3126 14468 3129
rect 14356 3118 14468 3126
rect 14502 3118 14536 3129
rect 14390 3095 14468 3118
rect 14534 3096 14536 3118
rect 14570 3123 14653 3130
rect 14570 3118 14604 3123
rect 14570 3096 14572 3118
rect 14390 3088 14500 3095
rect 14390 3084 14428 3088
rect 14356 3054 14428 3084
rect 14462 3084 14500 3088
rect 14534 3084 14572 3096
rect 14638 3089 14653 3123
rect 14606 3084 14653 3089
rect 14462 3061 14653 3084
rect 14462 3060 14536 3061
rect 14462 3054 14468 3060
rect 14356 3045 14468 3054
rect 14502 3045 14536 3060
rect 14390 3026 14468 3045
rect 14534 3027 14536 3045
rect 14570 3055 14653 3061
rect 14570 3045 14604 3055
rect 14570 3027 14572 3045
rect 14390 3016 14500 3026
rect 14390 3011 14428 3016
rect 14356 2982 14428 3011
rect 14462 3011 14500 3016
rect 14534 3011 14572 3027
rect 14638 3021 14653 3055
rect 14606 3011 14653 3021
rect 14462 2992 14653 3011
rect 14462 2991 14536 2992
rect 14462 2982 14468 2991
rect 14356 2972 14468 2982
rect 14502 2972 14536 2991
rect 14390 2957 14468 2972
rect 14534 2958 14536 2972
rect 14570 2987 14653 2992
rect 14570 2972 14604 2987
rect 14570 2958 14572 2972
rect 14390 2944 14500 2957
rect 14390 2938 14428 2944
rect 14356 2910 14428 2938
rect 14462 2938 14500 2944
rect 14534 2938 14572 2958
rect 14638 2953 14653 2987
rect 14606 2938 14653 2953
rect 14462 2923 14653 2938
rect 14462 2922 14536 2923
rect 14462 2910 14468 2922
rect 14356 2899 14468 2910
rect 14502 2899 14536 2922
rect 14390 2888 14468 2899
rect 14534 2889 14536 2899
rect 14570 2919 14653 2923
rect 14570 2899 14604 2919
rect 14570 2889 14572 2899
rect 14390 2872 14500 2888
rect 14390 2865 14428 2872
rect 14356 2838 14428 2865
rect 14462 2865 14500 2872
rect 14534 2865 14572 2889
rect 14638 2885 14653 2919
rect 14606 2865 14653 2885
rect 14462 2854 14653 2865
rect 14462 2853 14536 2854
rect 14462 2838 14468 2853
rect 14356 2826 14468 2838
rect 14502 2826 14536 2853
rect 14390 2819 14468 2826
rect 14534 2820 14536 2826
rect 14570 2851 14653 2854
rect 14570 2826 14604 2851
rect 14570 2820 14572 2826
rect 14390 2800 14500 2819
rect 14390 2792 14428 2800
rect 14356 2766 14428 2792
rect 14462 2792 14500 2800
rect 14534 2792 14572 2820
rect 14638 2817 14653 2851
rect 14606 2792 14653 2817
rect 14462 2785 14653 2792
rect 14462 2784 14536 2785
rect 14462 2766 14468 2784
rect 14356 2753 14468 2766
rect 14502 2753 14536 2784
rect 14390 2750 14468 2753
rect 14534 2751 14536 2753
rect 14570 2783 14653 2785
rect 14570 2753 14604 2783
rect 14570 2751 14572 2753
rect 14390 2728 14500 2750
rect 14390 2719 14428 2728
rect 14356 2694 14428 2719
rect 14462 2719 14500 2728
rect 14534 2719 14572 2751
rect 14638 2749 14653 2783
rect 14606 2719 14653 2749
rect 14462 2716 14653 2719
rect 14462 2715 14536 2716
rect 14462 2694 14468 2715
rect 14356 2681 14468 2694
rect 14502 2682 14536 2715
rect 14570 2715 14653 2716
rect 14570 2682 14604 2715
rect 14502 2681 14604 2682
rect 14638 2681 14653 2715
rect 14356 2680 14653 2681
rect 14390 2656 14500 2680
rect 14390 2646 14428 2656
rect 14356 2622 14428 2646
rect 14462 2646 14500 2656
rect 14534 2647 14572 2680
rect 14606 2647 14653 2680
rect 14534 2646 14536 2647
rect 14462 2622 14468 2646
rect 14356 2612 14468 2622
rect 14502 2613 14536 2646
rect 14570 2646 14572 2647
rect 14570 2613 14604 2646
rect 14638 2613 14653 2647
rect 14502 2612 14653 2613
rect 14356 2607 14653 2612
rect 14390 2584 14500 2607
rect 14390 2573 14428 2584
rect 14356 2550 14428 2573
rect 14462 2577 14500 2584
rect 14534 2578 14572 2607
rect 14606 2579 14653 2607
rect 14462 2550 14468 2577
rect 14534 2573 14536 2578
rect 14356 2543 14468 2550
rect 14502 2544 14536 2573
rect 14570 2573 14572 2578
rect 14570 2545 14604 2573
rect 14638 2545 14653 2579
rect 14570 2544 14653 2545
rect 14502 2543 14653 2544
rect 14356 2534 14653 2543
rect 14390 2512 14500 2534
rect 14390 2500 14428 2512
rect 14356 2482 14428 2500
rect 14390 2478 14428 2482
rect 14462 2508 14500 2512
rect 14534 2509 14572 2534
rect 14606 2511 14653 2534
rect 14462 2478 14468 2508
rect 14534 2500 14536 2509
rect 14390 2474 14468 2478
rect 14502 2475 14536 2500
rect 14570 2500 14572 2509
rect 14570 2477 14604 2500
rect 14638 2477 14653 2511
rect 14570 2475 14653 2477
rect 14502 2474 14653 2475
rect 14390 2461 14653 2474
rect 14390 2440 14500 2461
rect 14390 2427 14428 2440
rect 14356 2414 14428 2427
rect 14390 2406 14428 2414
rect 14462 2439 14500 2440
rect 14534 2440 14572 2461
rect 14606 2443 14653 2461
rect 14462 2406 14468 2439
rect 14534 2427 14536 2440
rect 14390 2405 14468 2406
rect 14502 2406 14536 2427
rect 14570 2427 14572 2440
rect 14570 2409 14604 2427
rect 14638 2409 14653 2443
rect 14570 2406 14653 2409
rect 14502 2405 14653 2406
rect 14390 2388 14653 2405
rect 14390 2370 14500 2388
rect 14534 2371 14572 2388
rect 14606 2375 14653 2388
rect 14390 2368 14468 2370
rect 14390 2354 14428 2368
rect 14356 2346 14428 2354
rect 14390 2334 14428 2346
rect 14462 2336 14468 2368
rect 14534 2354 14536 2371
rect 14502 2337 14536 2354
rect 14570 2354 14572 2371
rect 14570 2341 14604 2354
rect 14638 2341 14653 2375
rect 14570 2337 14653 2341
rect 14502 2336 14653 2337
rect 14462 2334 14653 2336
rect 14390 2315 14653 2334
rect 14390 2301 14500 2315
rect 14534 2302 14572 2315
rect 14606 2307 14653 2315
rect 14390 2296 14468 2301
rect 14390 2281 14428 2296
rect 14356 2278 14428 2281
rect 14390 2262 14428 2278
rect 14462 2267 14468 2296
rect 14534 2281 14536 2302
rect 14502 2268 14536 2281
rect 14570 2281 14572 2302
rect 14570 2273 14604 2281
rect 14638 2273 14653 2307
rect 14570 2268 14653 2273
rect 14502 2267 14653 2268
rect 14462 2262 14653 2267
rect 14390 2244 14653 2262
rect 14356 2242 14653 2244
rect 14390 2232 14500 2242
rect 14534 2233 14572 2242
rect 14606 2239 14653 2242
rect 14390 2224 14468 2232
rect 14390 2190 14428 2224
rect 14462 2198 14468 2224
rect 14534 2208 14536 2233
rect 14502 2199 14536 2208
rect 14570 2208 14572 2233
rect 14570 2205 14604 2208
rect 14638 2205 14653 2239
rect 14570 2199 14653 2205
rect 14502 2198 14653 2199
rect 14462 2190 14653 2198
rect 14390 2176 14653 2190
rect 14356 2171 14653 2176
rect 14356 2169 14604 2171
rect 14390 2163 14500 2169
rect 14534 2164 14572 2169
rect 14390 2152 14468 2163
rect 14390 2118 14428 2152
rect 14462 2129 14468 2152
rect 14534 2135 14536 2164
rect 14502 2130 14536 2135
rect 14570 2135 14572 2164
rect 14638 2137 14653 2171
rect 14606 2135 14653 2137
rect 14570 2130 14653 2135
rect 14502 2129 14653 2130
rect 14462 2118 14653 2129
rect 14390 2108 14653 2118
rect 14356 2103 14653 2108
rect 14356 2096 14604 2103
rect 14390 2094 14500 2096
rect 14534 2095 14572 2096
rect 14390 2080 14468 2094
rect 14390 2046 14428 2080
rect 14462 2060 14468 2080
rect 14534 2062 14536 2095
rect 14502 2061 14536 2062
rect 14570 2062 14572 2095
rect 14638 2069 14653 2103
rect 14606 2062 14653 2069
rect 14570 2061 14653 2062
rect 14502 2060 14653 2061
rect 14462 2046 14653 2060
rect 14390 2040 14653 2046
rect 14356 2035 14653 2040
rect 14356 2026 14604 2035
rect 14356 2025 14536 2026
rect 14356 2023 14468 2025
rect 14502 2023 14536 2025
rect 14390 2008 14468 2023
rect 14390 1974 14428 2008
rect 14462 1991 14468 2008
rect 14534 1992 14536 2023
rect 14570 2023 14604 2026
rect 14570 1992 14572 2023
rect 14638 2001 14653 2035
rect 14462 1989 14500 1991
rect 14534 1989 14572 1992
rect 14606 1989 14653 2001
rect 14462 1974 14653 1989
rect 14390 1972 14653 1974
rect 14356 1967 14653 1972
rect 14356 1957 14604 1967
rect 14356 1956 14536 1957
rect 14356 1950 14468 1956
rect 14502 1950 14536 1956
rect 14390 1936 14468 1950
rect 14390 1904 14428 1936
rect 14356 1902 14428 1904
rect 14462 1922 14468 1936
rect 14534 1923 14536 1950
rect 14570 1950 14604 1957
rect 14570 1923 14572 1950
rect 14638 1933 14653 1967
rect 14462 1916 14500 1922
rect 14534 1916 14572 1923
rect 14606 1916 14653 1933
rect 14462 1902 14653 1916
rect 14356 1899 14653 1902
rect 14356 1888 14604 1899
rect 14356 1887 14536 1888
rect 14356 1877 14468 1887
rect 14502 1877 14536 1887
rect 14390 1864 14468 1877
rect 14390 1836 14428 1864
rect 14356 1830 14428 1836
rect 14462 1853 14468 1864
rect 14534 1854 14536 1877
rect 14570 1877 14604 1888
rect 14570 1854 14572 1877
rect 14638 1865 14653 1899
rect 14462 1843 14500 1853
rect 14534 1843 14572 1854
rect 14606 1843 14653 1865
rect 14462 1831 14653 1843
rect 14462 1830 14604 1831
rect 14356 1819 14604 1830
rect 14356 1818 14536 1819
rect 14356 1804 14468 1818
rect 14502 1804 14536 1818
rect 14390 1792 14468 1804
rect 14390 1768 14428 1792
rect 14356 1758 14428 1768
rect 14462 1784 14468 1792
rect 14534 1785 14536 1804
rect 14570 1804 14604 1819
rect 14570 1785 14572 1804
rect 14638 1797 14653 1831
rect 14462 1770 14500 1784
rect 14534 1770 14572 1785
rect 14606 1770 14653 1797
rect 14462 1763 14653 1770
rect 14462 1758 14604 1763
rect 14356 1750 14604 1758
rect 14356 1749 14536 1750
rect 14356 1734 14468 1749
rect 14390 1720 14468 1734
rect 14502 1731 14536 1749
rect 14390 1697 14428 1720
rect 14356 1686 14428 1697
rect 14462 1715 14468 1720
rect 14534 1716 14536 1731
rect 14570 1731 14604 1750
rect 14570 1716 14572 1731
rect 14638 1729 14653 1763
rect 14462 1697 14500 1715
rect 14534 1697 14572 1716
rect 14606 1697 14653 1729
rect 14462 1695 14653 1697
rect 14462 1686 14604 1695
rect 14356 1681 14604 1686
rect 14356 1680 14536 1681
rect 14356 1666 14468 1680
rect 14390 1648 14468 1666
rect 14502 1658 14536 1680
rect 14390 1623 14428 1648
rect 14356 1614 14428 1623
rect 14462 1646 14468 1648
rect 14534 1647 14536 1658
rect 14570 1661 14604 1681
rect 14638 1661 14653 1695
rect 14570 1658 14653 1661
rect 14570 1647 14572 1658
rect 14462 1624 14500 1646
rect 14534 1624 14572 1647
rect 14606 1627 14653 1658
rect 14462 1614 14604 1624
rect 14356 1612 14604 1614
rect 14356 1611 14536 1612
rect 14356 1598 14468 1611
rect 14390 1577 14468 1598
rect 14502 1585 14536 1611
rect 14534 1578 14536 1585
rect 14570 1593 14604 1612
rect 14638 1593 14653 1627
rect 14570 1585 14653 1593
rect 14570 1578 14572 1585
rect 14390 1576 14500 1577
rect 14390 1549 14428 1576
rect 14356 1542 14428 1549
rect 14462 1551 14500 1576
rect 14534 1551 14572 1578
rect 14606 1559 14653 1585
rect 14462 1543 14604 1551
rect 14462 1542 14536 1543
rect 14356 1509 14468 1542
rect 14502 1512 14536 1542
rect 14390 1508 14468 1509
rect 14534 1509 14536 1512
rect 14570 1525 14604 1543
rect 14638 1525 14653 1559
rect 14570 1512 14653 1525
rect 14570 1509 14572 1512
rect 14390 1504 14500 1508
rect 14390 1475 14428 1504
rect 14356 1470 14428 1475
rect 14462 1478 14500 1504
rect 14534 1478 14572 1509
rect 14606 1491 14653 1512
rect 14462 1474 14604 1478
rect 14462 1473 14536 1474
rect 14462 1470 14468 1473
rect 14356 1439 14468 1470
rect 14502 1440 14536 1473
rect 14570 1457 14604 1474
rect 14638 1457 14653 1491
rect 14570 1440 14653 1457
rect 14502 1439 14653 1440
rect 14356 1435 14500 1439
rect 14390 1432 14500 1435
rect 14390 1401 14428 1432
rect 14356 1398 14428 1401
rect 14462 1405 14500 1432
rect 14534 1405 14572 1439
rect 14606 1423 14653 1439
rect 14462 1404 14536 1405
rect 14462 1398 14468 1404
rect 14356 1370 14468 1398
rect 14502 1371 14536 1404
rect 14570 1389 14604 1405
rect 14638 1389 14653 1423
rect 14570 1371 14653 1389
rect 14502 1370 14653 1371
rect 14356 1366 14653 1370
rect 14356 1361 14500 1366
rect 14390 1360 14500 1361
rect 14390 1327 14428 1360
rect 14356 1326 14428 1327
rect 14462 1335 14500 1360
rect 14534 1336 14572 1366
rect 14606 1355 14653 1366
rect 14462 1326 14468 1335
rect 14534 1332 14536 1336
rect 14356 1301 14468 1326
rect 14502 1302 14536 1332
rect 14570 1332 14572 1336
rect 14570 1321 14604 1332
rect 14638 1321 14653 1355
rect 14570 1302 14653 1321
rect 14502 1301 14653 1302
rect 14356 1293 14653 1301
rect 14356 1288 14500 1293
rect 14356 1287 14428 1288
rect 14390 1254 14428 1287
rect 14462 1266 14500 1288
rect 14534 1267 14572 1293
rect 14606 1287 14653 1293
rect 14462 1254 14468 1266
rect 14534 1259 14536 1267
rect 14390 1253 14468 1254
rect 14356 1232 14468 1253
rect 14502 1233 14536 1259
rect 14570 1259 14572 1267
rect 14570 1253 14604 1259
rect 14638 1253 14653 1287
rect 14570 1233 14653 1253
rect 14502 1232 14653 1233
rect 14356 1220 14653 1232
rect 14356 1216 14500 1220
rect 14356 1213 14428 1216
rect 14390 1182 14428 1213
rect 14462 1197 14500 1216
rect 14534 1198 14572 1220
rect 14606 1218 14653 1220
rect 14462 1182 14468 1197
rect 14534 1186 14536 1198
rect 14390 1179 14468 1182
rect 14356 1163 14468 1179
rect 14502 1164 14536 1186
rect 14570 1186 14572 1198
rect 14570 1184 14604 1186
rect 14638 1184 14653 1218
rect 14570 1164 14653 1184
rect 14502 1163 14653 1164
rect 14356 1149 14653 1163
rect 14356 1147 14604 1149
rect 14356 1144 14500 1147
rect 667 883 746 894
rect 667 867 780 883
rect 14356 1139 14428 1144
rect 14390 1110 14428 1139
rect 14462 1128 14500 1144
rect 14534 1129 14572 1147
rect 14462 1110 14468 1128
rect 14534 1113 14536 1129
rect 14390 1105 14468 1110
rect 14356 1094 14468 1105
rect 14502 1095 14536 1113
rect 14570 1113 14572 1129
rect 14638 1115 14653 1149
rect 14606 1113 14653 1115
rect 14570 1095 14653 1113
rect 14502 1094 14653 1095
rect 14356 1080 14653 1094
rect 14356 1074 14604 1080
rect 14356 1072 14500 1074
rect 14356 1065 14428 1072
rect 14390 1038 14428 1065
rect 14462 1059 14500 1072
rect 14534 1060 14572 1074
rect 14462 1038 14468 1059
rect 14534 1040 14536 1060
rect 14390 1031 14468 1038
rect 14356 1025 14468 1031
rect 14502 1026 14536 1040
rect 14570 1040 14572 1060
rect 14638 1046 14653 1080
rect 14606 1040 14653 1046
rect 14570 1026 14653 1040
rect 14502 1025 14653 1026
rect 14356 1011 14653 1025
rect 14356 1001 14604 1011
rect 14356 1000 14500 1001
rect 14356 991 14428 1000
rect 14390 966 14428 991
rect 14462 990 14500 1000
rect 14534 991 14572 1001
rect 14462 966 14468 990
rect 14534 967 14536 991
rect 14390 957 14468 966
rect 14356 956 14468 957
rect 14502 957 14536 967
rect 14570 967 14572 991
rect 14638 977 14653 1011
rect 14606 967 14653 977
rect 14570 957 14653 967
rect 14502 956 14653 957
rect 14356 942 14653 956
rect 14356 928 14604 942
rect 14356 917 14428 928
rect 14390 894 14428 917
rect 14462 921 14500 928
rect 14534 922 14572 928
rect 14462 894 14468 921
rect 14534 894 14536 922
rect 14390 887 14468 894
rect 14502 888 14536 894
rect 14570 894 14572 922
rect 14638 908 14653 942
rect 14606 894 14653 908
rect 14570 888 14653 894
rect 14502 887 14653 888
rect 14390 883 14653 887
rect 14356 873 14653 883
rect 14356 867 14604 873
rect 667 853 14604 867
rect 667 852 14536 853
rect 667 818 702 852
rect 736 820 771 852
rect 805 820 840 852
rect 874 820 909 852
rect 943 820 978 852
rect 1012 820 1047 852
rect 1081 820 1116 852
rect 1150 820 1185 852
rect 1219 820 1254 852
rect 1288 820 1323 852
rect 1357 820 1392 852
rect 1426 820 1461 852
rect 1495 820 1530 852
rect 1564 820 1599 852
rect 1633 820 1668 852
rect 1702 820 1737 852
rect 1771 820 1806 852
rect 1840 820 1875 852
rect 1909 820 1944 852
rect 1978 820 2013 852
rect 2047 820 2082 852
rect 2116 820 2151 852
rect 2185 820 2220 852
rect 2254 820 2289 852
rect 2323 820 2358 852
rect 2392 820 2427 852
rect 2461 820 2496 852
rect 2530 820 2565 852
rect 2599 820 2634 852
rect 2668 820 2703 852
rect 2737 820 2772 852
rect 743 818 771 820
rect 816 818 840 820
rect 889 818 909 820
rect 599 786 709 818
rect 743 786 782 818
rect 816 786 855 818
rect 889 786 928 818
rect 599 784 928 786
rect 482 750 565 769
rect 599 750 634 784
rect 668 750 703 784
rect 737 750 772 784
rect 806 750 841 784
rect 875 750 910 784
rect 14502 819 14536 852
rect 14570 839 14604 853
rect 14638 839 14653 873
rect 14570 819 14653 839
rect 14502 804 14653 819
rect 14502 784 14604 804
rect 14570 770 14604 784
rect 14638 770 14653 804
rect 14570 750 14653 770
rect 482 748 928 750
rect 482 716 709 748
rect 743 716 782 748
rect 816 716 855 748
rect 889 716 928 748
rect 482 682 516 716
rect 550 682 585 716
rect 619 682 654 716
rect 688 714 709 716
rect 757 714 782 716
rect 826 714 855 716
rect 895 714 928 716
rect 14551 735 14653 750
rect 688 682 723 714
rect 757 682 792 714
rect 826 682 861 714
rect 895 682 930 714
rect 964 682 999 714
rect 1033 682 1068 714
rect 1102 682 1137 714
rect 1171 682 1206 714
rect 1240 682 1275 714
rect 1309 682 1344 714
rect 1378 682 1413 714
rect 1447 682 1482 714
rect 1516 682 1551 714
rect 1585 682 1620 714
rect 1654 682 1689 714
rect 1723 682 1758 714
rect 1792 682 1827 714
rect 1861 682 1896 714
rect 1930 682 1965 714
rect 1999 682 2034 714
rect 2068 682 2103 714
rect 2137 682 2172 714
rect 2206 682 2241 714
rect 2275 682 2310 714
rect 2344 682 2379 714
rect 2413 682 2448 714
rect 2482 682 2517 714
rect 2551 682 2586 714
rect 2620 682 2655 714
rect 2689 682 2724 714
rect 2758 682 2793 714
rect 2827 682 2862 714
rect 2896 682 2931 714
rect 2965 682 3000 714
rect 3034 682 3069 714
rect 3103 682 3138 714
rect 3172 682 3207 714
rect 3241 682 3276 714
rect 3310 682 3345 714
rect 3379 682 3414 714
rect 3448 682 3483 714
rect 3517 682 3552 714
rect 3586 682 3621 714
rect 3655 682 3690 714
rect 3724 682 3759 714
rect 3793 682 3828 714
rect 3862 682 3897 714
rect 3931 682 3966 714
rect 4000 682 4035 714
rect 4069 682 4104 714
rect 4138 682 4173 714
rect 4207 682 4242 714
rect 4276 682 4311 714
rect 4345 682 4380 714
rect 4414 682 4449 714
rect 4483 682 4518 714
rect 4552 682 4587 714
rect 4621 682 4656 714
rect 4690 682 4725 714
rect 14551 701 14604 735
rect 14638 701 14653 735
rect 14551 682 14653 701
rect 482 667 14653 682
rect 14806 4645 14835 4679
rect 14806 4577 14835 4611
rect 14806 4509 14835 4543
rect 14806 4441 14835 4475
rect 14806 4373 14835 4407
rect 14806 4305 14835 4339
rect 14806 4237 14835 4271
rect 14806 4169 14835 4203
rect 14806 4101 14835 4135
rect 14806 4033 14835 4067
rect 14806 3965 14835 3999
rect 14806 3897 14835 3931
rect 14806 3829 14835 3863
rect 14806 3761 14835 3795
rect 14806 3693 14835 3727
rect 14806 3625 14835 3659
rect 14806 3557 14835 3591
rect 14806 3489 14835 3523
rect 14806 3421 14835 3455
rect 14806 3353 14835 3387
rect 14806 3285 14835 3319
rect 14806 3217 14835 3251
rect 14806 3149 14835 3183
rect 14806 3081 14835 3115
rect 14806 3013 14835 3047
rect 14806 2945 14835 2979
rect 14806 2877 14835 2911
rect 14806 2809 14835 2843
rect 14806 2741 14835 2775
rect 14806 2673 14835 2707
rect 14806 2605 14835 2639
rect 14806 2537 14835 2571
rect 14806 2469 14835 2503
rect 14806 2401 14835 2435
rect 14806 2333 14835 2367
rect 14806 2265 14835 2299
rect 14806 2197 14835 2231
rect 14806 2129 14835 2163
rect 14806 2061 14835 2095
rect 14806 1993 14835 2027
rect 14806 1925 14835 1959
rect 14806 1857 14835 1891
rect 14806 1789 14835 1823
rect 14806 1721 14835 1755
rect 14806 1653 14835 1687
rect 14806 1585 14835 1619
rect 14806 1517 14835 1551
rect 14806 1468 14835 1483
rect 14806 1449 14907 1468
rect 14840 1429 14906 1449
rect 14869 1415 14906 1429
rect 14806 1395 14835 1415
rect 14869 1395 14907 1415
rect 14806 1381 14907 1395
rect 14840 1356 14906 1381
rect 14869 1347 14906 1356
rect 14806 1322 14835 1347
rect 14869 1322 14907 1347
rect 14806 1313 14907 1322
rect 14840 1283 14906 1313
rect 14869 1279 14906 1283
rect 14806 1249 14835 1279
rect 14869 1249 14907 1279
rect 14806 1245 14907 1249
rect 14840 1211 14906 1245
rect 14806 1210 14907 1211
rect 14806 1177 14835 1210
rect 14869 1177 14907 1210
rect 14869 1176 14906 1177
rect 14840 1143 14906 1176
rect 14806 1137 14907 1143
rect 14806 1109 14835 1137
rect 14869 1109 14907 1137
rect 14869 1103 14906 1109
rect 14840 1075 14906 1103
rect 14806 1064 14907 1075
rect 14806 1041 14835 1064
rect 14869 1041 14907 1064
rect 14869 1030 14906 1041
rect 14840 1007 14906 1030
rect 14806 991 14907 1007
rect 14806 973 14835 991
rect 14869 973 14907 991
rect 14869 957 14906 973
rect 14840 939 14906 957
rect 14806 918 14907 939
rect 14806 905 14835 918
rect 14869 905 14907 918
rect 14869 884 14906 905
rect 14840 871 14906 884
rect 14806 845 14907 871
rect 14806 837 14835 845
rect 14869 837 14907 845
rect 14869 811 14906 837
rect 14840 803 14906 811
rect 14806 772 14907 803
rect 14806 769 14835 772
rect 14869 769 14907 772
rect 14869 738 14906 769
rect 14840 735 14906 738
rect 14806 701 14907 735
rect 14840 699 14906 701
rect 14869 667 14906 699
rect 303 607 329 641
rect 295 599 329 607
rect 231 567 329 599
rect 231 533 269 567
rect 303 533 329 567
rect 231 509 329 533
rect 14806 665 14835 667
rect 14869 665 14907 667
rect 14806 633 14907 665
rect 14840 626 14906 633
rect 14869 599 14906 626
rect 14806 592 14835 599
rect 14869 592 14907 599
rect 14806 553 14907 592
rect 14806 519 14835 553
rect 14869 519 14907 553
rect 14806 509 14907 519
rect 14847 420 14907 509
rect 14847 407 14940 420
rect 231 375 14939 407
rect 231 341 361 375
rect 395 341 434 375
rect 468 341 507 375
rect 541 341 580 375
rect 614 341 653 375
rect 687 341 726 375
rect 760 341 799 375
rect 833 341 872 375
rect 906 341 945 375
rect 979 341 1018 375
rect 1052 341 1091 375
rect 1125 341 1164 375
rect 1198 341 1237 375
rect 1271 341 1310 375
rect 1344 341 1383 375
rect 1417 341 1456 375
rect 1490 341 1529 375
rect 1563 341 1602 375
rect 1636 341 1675 375
rect 1709 341 1748 375
rect 1782 341 1821 375
rect 1855 341 1894 375
rect 1928 341 1967 375
rect 2001 341 2040 375
rect 2074 341 2113 375
rect 2147 341 2186 375
rect 2220 341 2259 375
rect 2293 341 2332 375
rect 2366 341 2405 375
rect 2439 341 2478 375
rect 2512 341 2551 375
rect 2585 341 2624 375
rect 2658 341 2697 375
rect 2731 341 2770 375
rect 2804 341 2843 375
rect 2877 341 2916 375
rect 2950 341 2989 375
rect 3023 341 3062 375
rect 3096 341 3135 375
rect 3169 341 3208 375
rect 3242 341 3281 375
rect 3315 341 3354 375
rect 3388 341 3427 375
rect 3461 341 3500 375
rect 3534 341 3573 375
rect 3607 341 3646 375
rect 3680 341 3719 375
rect 3753 341 3792 375
rect 3826 341 3865 375
rect 3899 341 3938 375
rect 3972 341 4011 375
rect 4045 341 4084 375
rect 4118 341 4157 375
rect 4191 341 4229 375
rect 4263 341 4301 375
rect 4335 341 4373 375
rect 4407 341 4445 375
rect 4479 341 4517 375
rect 4551 341 4589 375
rect 4623 341 4661 375
rect 4695 341 4733 375
rect 4767 341 4805 375
rect 4839 341 4877 375
rect 4911 341 4949 375
rect 4983 341 5021 375
rect 5055 341 5093 375
rect 5127 341 5165 375
rect 5199 341 5237 375
rect 5271 341 5309 375
rect 5343 341 5381 375
rect 5415 341 5453 375
rect 5487 341 5525 375
rect 5559 341 5597 375
rect 5631 341 5669 375
rect 5703 341 5741 375
rect 5775 341 5813 375
rect 5847 341 5885 375
rect 5919 341 5957 375
rect 5991 341 6029 375
rect 6063 341 6101 375
rect 6135 341 6173 375
rect 6207 341 6245 375
rect 6279 341 6317 375
rect 6351 341 6389 375
rect 6423 341 6461 375
rect 6495 341 6533 375
rect 6567 341 6605 375
rect 6639 341 6677 375
rect 6711 341 6749 375
rect 6783 341 6821 375
rect 6855 341 6893 375
rect 6927 341 6965 375
rect 6999 341 7037 375
rect 7071 341 7109 375
rect 7143 341 7181 375
rect 7215 341 7253 375
rect 7287 341 7325 375
rect 7359 341 7397 375
rect 7431 341 7469 375
rect 7503 341 7541 375
rect 7575 341 7613 375
rect 7647 341 7685 375
rect 7719 341 7757 375
rect 7791 341 7829 375
rect 7863 341 7901 375
rect 7935 341 7973 375
rect 8007 341 8045 375
rect 8079 341 8117 375
rect 8151 341 8189 375
rect 8223 341 8261 375
rect 8295 341 8333 375
rect 8367 341 8405 375
rect 8439 341 8477 375
rect 8511 341 8549 375
rect 8583 341 8621 375
rect 8655 341 8693 375
rect 8727 341 8765 375
rect 8799 341 8837 375
rect 8871 341 8909 375
rect 8943 341 8981 375
rect 9015 341 9053 375
rect 9087 341 9125 375
rect 9159 341 9197 375
rect 9231 341 9269 375
rect 9303 341 9341 375
rect 9375 341 9413 375
rect 9447 341 9485 375
rect 9519 341 9557 375
rect 9591 341 9629 375
rect 9663 341 9701 375
rect 9735 341 9773 375
rect 9807 341 9845 375
rect 9879 341 9917 375
rect 9951 341 9989 375
rect 10023 341 10061 375
rect 10095 341 10133 375
rect 10167 341 10205 375
rect 10239 341 10277 375
rect 10311 341 10349 375
rect 10383 341 10421 375
rect 10455 341 10493 375
rect 10527 341 10565 375
rect 10599 341 10637 375
rect 10671 341 10709 375
rect 10743 341 10781 375
rect 10815 341 10853 375
rect 10887 341 10925 375
rect 10959 341 10997 375
rect 11031 341 11069 375
rect 11103 341 11141 375
rect 11175 341 11213 375
rect 11247 341 11285 375
rect 11319 341 11357 375
rect 11391 341 11429 375
rect 11463 341 11501 375
rect 11535 341 11573 375
rect 11607 341 11645 375
rect 11679 341 11717 375
rect 11751 341 11789 375
rect 11823 341 11861 375
rect 11895 341 11933 375
rect 11967 341 12005 375
rect 12039 341 12077 375
rect 12111 341 12149 375
rect 12183 341 12221 375
rect 12255 341 12293 375
rect 12327 341 12365 375
rect 12399 341 12437 375
rect 12471 341 12509 375
rect 12543 341 12581 375
rect 12615 341 12653 375
rect 12687 341 12725 375
rect 12759 341 12797 375
rect 12831 341 12869 375
rect 12903 341 12941 375
rect 12975 341 13013 375
rect 13047 341 13085 375
rect 13119 341 13157 375
rect 13191 341 13229 375
rect 13263 341 13301 375
rect 13335 341 13373 375
rect 13407 341 13445 375
rect 13479 341 13517 375
rect 13551 341 13589 375
rect 13623 341 13661 375
rect 13695 341 13733 375
rect 13767 341 13805 375
rect 13839 341 13877 375
rect 13911 341 13949 375
rect 13983 341 14021 375
rect 14055 341 14093 375
rect 14127 341 14165 375
rect 14199 341 14237 375
rect 14271 341 14309 375
rect 14343 341 14381 375
rect 14415 341 14453 375
rect 14487 341 14525 375
rect 14559 341 14597 375
rect 14631 341 14669 375
rect 14703 341 14741 375
rect 14775 341 14939 375
rect 231 331 14939 341
rect 15 309 14939 331
rect 159 307 14939 309
<< viali >>
rect 361 5082 395 5111
rect 434 5082 468 5111
rect 507 5082 541 5111
rect 580 5082 614 5111
rect 653 5082 687 5111
rect 726 5082 760 5111
rect 799 5082 833 5111
rect 872 5082 906 5111
rect 945 5082 979 5111
rect 1018 5082 1052 5111
rect 1091 5082 1125 5111
rect 1164 5082 1198 5111
rect 1237 5082 1271 5111
rect 1310 5082 1344 5111
rect 1383 5082 1417 5111
rect 1456 5082 1490 5111
rect 1529 5082 1563 5111
rect 1602 5082 1636 5111
rect 1675 5082 1709 5111
rect 1748 5082 1782 5111
rect 1821 5082 1855 5111
rect 1894 5082 1928 5111
rect 1967 5082 2001 5111
rect 2040 5082 2074 5111
rect 2113 5082 2147 5111
rect 2186 5082 2220 5111
rect 2259 5082 2293 5111
rect 2332 5082 2366 5111
rect 2405 5082 2439 5111
rect 2478 5082 2512 5111
rect 2551 5082 2585 5111
rect 2624 5082 2658 5111
rect 2697 5082 2731 5111
rect 2770 5082 2804 5111
rect 2843 5082 2877 5111
rect 2916 5082 2950 5111
rect 2989 5082 3023 5111
rect 3062 5082 3096 5111
rect 3135 5082 3169 5111
rect 3208 5082 3242 5111
rect 3281 5082 3315 5111
rect 3354 5082 3388 5111
rect 3427 5082 3461 5111
rect 3500 5082 3534 5111
rect 3573 5082 3607 5111
rect 3646 5082 3680 5111
rect 3719 5082 3753 5111
rect 3792 5082 3826 5111
rect 3865 5082 3899 5111
rect 3938 5082 3972 5111
rect 4011 5082 4045 5111
rect 4084 5082 4118 5111
rect 4157 5082 4191 5111
rect 4229 5082 4263 5111
rect 4301 5082 4335 5111
rect 4373 5082 4407 5111
rect 4445 5082 4479 5111
rect 4517 5082 4551 5111
rect 4589 5082 4623 5111
rect 4661 5082 4695 5111
rect 4733 5082 4767 5111
rect 4805 5082 4839 5111
rect 4877 5082 4911 5111
rect 4949 5082 4983 5111
rect 5021 5082 5055 5111
rect 5093 5082 5127 5111
rect 5165 5082 5199 5111
rect 5237 5082 5271 5111
rect 5309 5082 5343 5111
rect 5381 5082 5415 5111
rect 5453 5082 5487 5111
rect 5525 5082 5559 5111
rect 5597 5082 5631 5111
rect 5669 5082 5703 5111
rect 5741 5082 5775 5111
rect 5813 5082 5847 5111
rect 5885 5082 5919 5111
rect 5957 5082 5991 5111
rect 6029 5082 6063 5111
rect 6101 5082 6135 5111
rect 6173 5082 6207 5111
rect 6245 5082 6279 5111
rect 6317 5082 6351 5111
rect 6389 5082 6423 5111
rect 6461 5082 6495 5111
rect 6533 5082 6567 5111
rect 6605 5082 6639 5111
rect 6677 5082 6711 5111
rect 6749 5082 6783 5111
rect 6821 5082 6855 5111
rect 6893 5082 6927 5111
rect 6965 5082 6999 5111
rect 7037 5082 7071 5111
rect 7109 5082 7143 5111
rect 7181 5082 7215 5111
rect 7253 5082 7287 5111
rect 7325 5082 7359 5111
rect 7397 5082 7431 5111
rect 7469 5082 7503 5111
rect 7541 5082 7575 5111
rect 7613 5082 7647 5111
rect 7685 5082 7719 5111
rect 7757 5082 7791 5111
rect 7829 5082 7863 5111
rect 7901 5082 7935 5111
rect 7973 5082 8007 5111
rect 8045 5082 8079 5111
rect 8117 5082 8151 5111
rect 8189 5082 8223 5111
rect 8261 5082 8295 5111
rect 8333 5082 8367 5111
rect 8405 5082 8439 5111
rect 8477 5082 8511 5111
rect 8549 5082 8583 5111
rect 8621 5082 8655 5111
rect 8693 5082 8727 5111
rect 8765 5082 8799 5111
rect 8837 5082 8871 5111
rect 8909 5082 8943 5111
rect 8981 5082 9015 5111
rect 9053 5082 9087 5111
rect 9125 5082 9159 5111
rect 9197 5082 9231 5111
rect 9269 5082 9303 5111
rect 9341 5082 9375 5111
rect 9413 5082 9447 5111
rect 9485 5082 9519 5111
rect 9557 5082 9591 5111
rect 9629 5082 9663 5111
rect 9701 5082 9735 5111
rect 9773 5082 9807 5111
rect 9845 5082 9879 5111
rect 9917 5082 9951 5111
rect 9989 5082 10023 5111
rect 10061 5082 10095 5111
rect 10133 5082 10167 5111
rect 10205 5082 10239 5111
rect 10277 5082 10311 5111
rect 10349 5082 10383 5111
rect 10421 5082 10455 5111
rect 10493 5082 10527 5111
rect 10565 5082 10599 5111
rect 10637 5082 10671 5111
rect 10709 5082 10743 5111
rect 10781 5082 10815 5111
rect 10853 5082 10887 5111
rect 10925 5082 10959 5111
rect 10997 5082 11031 5111
rect 11069 5082 11103 5111
rect 11141 5082 11175 5111
rect 11213 5082 11247 5111
rect 11285 5082 11319 5111
rect 11357 5082 11391 5111
rect 11429 5082 11463 5111
rect 11501 5082 11535 5111
rect 11573 5082 11607 5111
rect 11645 5082 11679 5111
rect 11717 5082 11751 5111
rect 11789 5082 11823 5111
rect 11861 5082 11895 5111
rect 11933 5082 11967 5111
rect 12005 5082 12039 5111
rect 12077 5082 12111 5111
rect 12149 5082 12183 5111
rect 12221 5082 12255 5111
rect 12293 5082 12327 5111
rect 12365 5082 12399 5111
rect 12437 5082 12471 5111
rect 12509 5082 12543 5111
rect 12581 5082 12615 5111
rect 12653 5082 12687 5111
rect 12725 5082 12759 5111
rect 12797 5082 12831 5111
rect 12869 5082 12903 5111
rect 12941 5082 12975 5111
rect 13013 5082 13047 5111
rect 13085 5082 13119 5111
rect 13157 5082 13191 5111
rect 13229 5082 13263 5111
rect 13301 5082 13335 5111
rect 13373 5082 13407 5111
rect 13445 5082 13479 5111
rect 13517 5082 13551 5111
rect 13589 5082 13623 5111
rect 13661 5082 13695 5111
rect 13733 5082 13767 5111
rect 13805 5082 13839 5111
rect 13877 5082 13911 5111
rect 13949 5082 13983 5111
rect 14021 5082 14055 5111
rect 14093 5082 14127 5111
rect 14165 5082 14199 5111
rect 14237 5082 14271 5111
rect 14309 5082 14343 5111
rect 14381 5082 14415 5111
rect 14453 5082 14487 5111
rect 14525 5082 14559 5111
rect 14597 5082 14631 5111
rect 14669 5082 14703 5111
rect 14741 5082 14775 5111
rect 361 5077 388 5082
rect 388 5077 395 5082
rect 434 5077 456 5082
rect 456 5077 468 5082
rect 507 5077 524 5082
rect 524 5077 541 5082
rect 580 5077 592 5082
rect 592 5077 614 5082
rect 653 5077 660 5082
rect 660 5077 687 5082
rect 726 5077 728 5082
rect 728 5077 760 5082
rect 799 5077 830 5082
rect 830 5077 833 5082
rect 872 5077 898 5082
rect 898 5077 906 5082
rect 945 5077 966 5082
rect 966 5077 979 5082
rect 1018 5077 1034 5082
rect 1034 5077 1052 5082
rect 1091 5077 1102 5082
rect 1102 5077 1125 5082
rect 1164 5077 1170 5082
rect 1170 5077 1198 5082
rect 1237 5077 1238 5082
rect 1238 5077 1271 5082
rect 1310 5077 1340 5082
rect 1340 5077 1344 5082
rect 1383 5077 1408 5082
rect 1408 5077 1417 5082
rect 1456 5077 1476 5082
rect 1476 5077 1490 5082
rect 1529 5077 1544 5082
rect 1544 5077 1563 5082
rect 1602 5077 1612 5082
rect 1612 5077 1636 5082
rect 1675 5077 1680 5082
rect 1680 5077 1709 5082
rect 1748 5077 1782 5082
rect 1821 5077 1850 5082
rect 1850 5077 1855 5082
rect 1894 5077 1918 5082
rect 1918 5077 1928 5082
rect 1967 5077 1986 5082
rect 1986 5077 2001 5082
rect 2040 5077 2054 5082
rect 2054 5077 2074 5082
rect 2113 5077 2122 5082
rect 2122 5077 2147 5082
rect 2186 5077 2190 5082
rect 2190 5077 2220 5082
rect 2259 5077 2292 5082
rect 2292 5077 2293 5082
rect 2332 5077 2360 5082
rect 2360 5077 2366 5082
rect 2405 5077 2428 5082
rect 2428 5077 2439 5082
rect 2478 5077 2496 5082
rect 2496 5077 2512 5082
rect 2551 5077 2564 5082
rect 2564 5077 2585 5082
rect 2624 5077 2632 5082
rect 2632 5077 2658 5082
rect 2697 5077 2700 5082
rect 2700 5077 2731 5082
rect 2770 5077 2802 5082
rect 2802 5077 2804 5082
rect 2843 5077 2870 5082
rect 2870 5077 2877 5082
rect 2916 5077 2938 5082
rect 2938 5077 2950 5082
rect 2989 5077 3006 5082
rect 3006 5077 3023 5082
rect 3062 5077 3074 5082
rect 3074 5077 3096 5082
rect 3135 5077 3142 5082
rect 3142 5077 3169 5082
rect 3208 5077 3210 5082
rect 3210 5077 3242 5082
rect 3281 5077 3312 5082
rect 3312 5077 3315 5082
rect 3354 5077 3380 5082
rect 3380 5077 3388 5082
rect 3427 5077 3448 5082
rect 3448 5077 3461 5082
rect 3500 5077 3516 5082
rect 3516 5077 3534 5082
rect 3573 5077 3584 5082
rect 3584 5077 3607 5082
rect 3646 5077 3652 5082
rect 3652 5077 3680 5082
rect 3719 5077 3720 5082
rect 3720 5077 3753 5082
rect 3792 5077 3822 5082
rect 3822 5077 3826 5082
rect 3865 5077 3890 5082
rect 3890 5077 3899 5082
rect 3938 5077 3958 5082
rect 3958 5077 3972 5082
rect 4011 5077 4026 5082
rect 4026 5077 4045 5082
rect 4084 5077 4094 5082
rect 4094 5077 4118 5082
rect 4157 5077 4162 5082
rect 4162 5077 4191 5082
rect 4229 5077 4230 5082
rect 4230 5077 4263 5082
rect 4301 5077 4332 5082
rect 4332 5077 4335 5082
rect 4373 5077 4400 5082
rect 4400 5077 4407 5082
rect 4445 5077 4468 5082
rect 4468 5077 4479 5082
rect 4517 5077 4536 5082
rect 4536 5077 4551 5082
rect 4589 5077 4604 5082
rect 4604 5077 4623 5082
rect 4661 5077 4672 5082
rect 4672 5077 4695 5082
rect 4733 5077 4740 5082
rect 4740 5077 4767 5082
rect 4805 5077 4808 5082
rect 4808 5077 4839 5082
rect 4877 5077 4910 5082
rect 4910 5077 4911 5082
rect 4949 5077 4978 5082
rect 4978 5077 4983 5082
rect 5021 5077 5046 5082
rect 5046 5077 5055 5082
rect 5093 5077 5114 5082
rect 5114 5077 5127 5082
rect 5165 5077 5182 5082
rect 5182 5077 5199 5082
rect 5237 5077 5250 5082
rect 5250 5077 5271 5082
rect 5309 5077 5318 5082
rect 5318 5077 5343 5082
rect 5381 5077 5386 5082
rect 5386 5077 5415 5082
rect 5453 5077 5454 5082
rect 5454 5077 5487 5082
rect 5525 5077 5556 5082
rect 5556 5077 5559 5082
rect 5597 5077 5624 5082
rect 5624 5077 5631 5082
rect 5669 5077 5692 5082
rect 5692 5077 5703 5082
rect 5741 5077 5760 5082
rect 5760 5077 5775 5082
rect 5813 5077 5828 5082
rect 5828 5077 5847 5082
rect 5885 5077 5896 5082
rect 5896 5077 5919 5082
rect 5957 5077 5964 5082
rect 5964 5077 5991 5082
rect 6029 5077 6032 5082
rect 6032 5077 6063 5082
rect 6101 5077 6134 5082
rect 6134 5077 6135 5082
rect 6173 5077 6202 5082
rect 6202 5077 6207 5082
rect 6245 5077 6270 5082
rect 6270 5077 6279 5082
rect 6317 5077 6338 5082
rect 6338 5077 6351 5082
rect 6389 5077 6406 5082
rect 6406 5077 6423 5082
rect 6461 5077 6474 5082
rect 6474 5077 6495 5082
rect 6533 5077 6542 5082
rect 6542 5077 6567 5082
rect 6605 5077 6610 5082
rect 6610 5077 6639 5082
rect 6677 5077 6678 5082
rect 6678 5077 6711 5082
rect 6749 5077 6780 5082
rect 6780 5077 6783 5082
rect 6821 5077 6848 5082
rect 6848 5077 6855 5082
rect 6893 5077 6916 5082
rect 6916 5077 6927 5082
rect 6965 5077 6984 5082
rect 6984 5077 6999 5082
rect 7037 5077 7052 5082
rect 7052 5077 7071 5082
rect 7109 5077 7120 5082
rect 7120 5077 7143 5082
rect 7181 5077 7188 5082
rect 7188 5077 7215 5082
rect 7253 5077 7256 5082
rect 7256 5077 7287 5082
rect 7325 5077 7358 5082
rect 7358 5077 7359 5082
rect 7397 5077 7426 5082
rect 7426 5077 7431 5082
rect 7469 5077 7494 5082
rect 7494 5077 7503 5082
rect 7541 5077 7562 5082
rect 7562 5077 7575 5082
rect 7613 5077 7630 5082
rect 7630 5077 7647 5082
rect 7685 5077 7698 5082
rect 7698 5077 7719 5082
rect 7757 5077 7766 5082
rect 7766 5077 7791 5082
rect 7829 5077 7834 5082
rect 7834 5077 7863 5082
rect 7901 5077 7902 5082
rect 7902 5077 7935 5082
rect 7973 5077 8004 5082
rect 8004 5077 8007 5082
rect 8045 5077 8072 5082
rect 8072 5077 8079 5082
rect 8117 5077 8140 5082
rect 8140 5077 8151 5082
rect 8189 5077 8208 5082
rect 8208 5077 8223 5082
rect 8261 5077 8276 5082
rect 8276 5077 8295 5082
rect 8333 5077 8344 5082
rect 8344 5077 8367 5082
rect 8405 5077 8412 5082
rect 8412 5077 8439 5082
rect 8477 5077 8480 5082
rect 8480 5077 8511 5082
rect 8549 5077 8582 5082
rect 8582 5077 8583 5082
rect 8621 5077 8650 5082
rect 8650 5077 8655 5082
rect 8693 5077 8718 5082
rect 8718 5077 8727 5082
rect 8765 5077 8786 5082
rect 8786 5077 8799 5082
rect 8837 5077 8854 5082
rect 8854 5077 8871 5082
rect 8909 5077 8922 5082
rect 8922 5077 8943 5082
rect 8981 5077 8990 5082
rect 8990 5077 9015 5082
rect 9053 5077 9058 5082
rect 9058 5077 9087 5082
rect 9125 5077 9126 5082
rect 9126 5077 9159 5082
rect 9197 5077 9228 5082
rect 9228 5077 9231 5082
rect 9269 5077 9296 5082
rect 9296 5077 9303 5082
rect 9341 5077 9364 5082
rect 9364 5077 9375 5082
rect 9413 5077 9432 5082
rect 9432 5077 9447 5082
rect 9485 5077 9500 5082
rect 9500 5077 9519 5082
rect 9557 5077 9568 5082
rect 9568 5077 9591 5082
rect 9629 5077 9636 5082
rect 9636 5077 9663 5082
rect 9701 5077 9704 5082
rect 9704 5077 9735 5082
rect 9773 5077 9806 5082
rect 9806 5077 9807 5082
rect 9845 5077 9874 5082
rect 9874 5077 9879 5082
rect 9917 5077 9942 5082
rect 9942 5077 9951 5082
rect 9989 5077 10010 5082
rect 10010 5077 10023 5082
rect 10061 5077 10078 5082
rect 10078 5077 10095 5082
rect 10133 5077 10146 5082
rect 10146 5077 10167 5082
rect 10205 5077 10214 5082
rect 10214 5077 10239 5082
rect 10277 5077 10282 5082
rect 10282 5077 10311 5082
rect 10349 5077 10350 5082
rect 10350 5077 10383 5082
rect 10421 5077 10452 5082
rect 10452 5077 10455 5082
rect 10493 5077 10520 5082
rect 10520 5077 10527 5082
rect 10565 5077 10588 5082
rect 10588 5077 10599 5082
rect 10637 5077 10656 5082
rect 10656 5077 10671 5082
rect 10709 5077 10724 5082
rect 10724 5077 10743 5082
rect 10781 5077 10792 5082
rect 10792 5077 10815 5082
rect 10853 5077 10860 5082
rect 10860 5077 10887 5082
rect 10925 5077 10928 5082
rect 10928 5077 10959 5082
rect 10997 5077 11030 5082
rect 11030 5077 11031 5082
rect 11069 5077 11098 5082
rect 11098 5077 11103 5082
rect 11141 5077 11166 5082
rect 11166 5077 11175 5082
rect 11213 5077 11234 5082
rect 11234 5077 11247 5082
rect 11285 5077 11302 5082
rect 11302 5077 11319 5082
rect 11357 5077 11370 5082
rect 11370 5077 11391 5082
rect 11429 5077 11438 5082
rect 11438 5077 11463 5082
rect 11501 5077 11506 5082
rect 11506 5077 11535 5082
rect 11573 5077 11574 5082
rect 11574 5077 11607 5082
rect 11645 5077 11676 5082
rect 11676 5077 11679 5082
rect 11717 5077 11744 5082
rect 11744 5077 11751 5082
rect 11789 5077 11812 5082
rect 11812 5077 11823 5082
rect 11861 5077 11880 5082
rect 11880 5077 11895 5082
rect 11933 5077 11948 5082
rect 11948 5077 11967 5082
rect 12005 5077 12016 5082
rect 12016 5077 12039 5082
rect 12077 5077 12084 5082
rect 12084 5077 12111 5082
rect 12149 5077 12152 5082
rect 12152 5077 12183 5082
rect 12221 5077 12254 5082
rect 12254 5077 12255 5082
rect 12293 5077 12322 5082
rect 12322 5077 12327 5082
rect 12365 5077 12390 5082
rect 12390 5077 12399 5082
rect 12437 5077 12458 5082
rect 12458 5077 12471 5082
rect 12509 5077 12526 5082
rect 12526 5077 12543 5082
rect 12581 5077 12594 5082
rect 12594 5077 12615 5082
rect 12653 5077 12662 5082
rect 12662 5077 12687 5082
rect 12725 5077 12730 5082
rect 12730 5077 12759 5082
rect 12797 5077 12798 5082
rect 12798 5077 12831 5082
rect 12869 5077 12900 5082
rect 12900 5077 12903 5082
rect 12941 5077 12968 5082
rect 12968 5077 12975 5082
rect 13013 5077 13036 5082
rect 13036 5077 13047 5082
rect 13085 5077 13104 5082
rect 13104 5077 13119 5082
rect 13157 5077 13172 5082
rect 13172 5077 13191 5082
rect 13229 5077 13240 5082
rect 13240 5077 13263 5082
rect 13301 5077 13308 5082
rect 13308 5077 13335 5082
rect 13373 5077 13376 5082
rect 13376 5077 13407 5082
rect 13445 5077 13478 5082
rect 13478 5077 13479 5082
rect 13517 5077 13546 5082
rect 13546 5077 13551 5082
rect 13589 5077 13614 5082
rect 13614 5077 13623 5082
rect 13661 5077 13682 5082
rect 13682 5077 13695 5082
rect 13733 5077 13750 5082
rect 13750 5077 13767 5082
rect 13805 5077 13818 5082
rect 13818 5077 13839 5082
rect 13877 5077 13886 5082
rect 13886 5077 13911 5082
rect 13949 5077 13954 5082
rect 13954 5077 13983 5082
rect 14021 5077 14022 5082
rect 14022 5077 14055 5082
rect 14093 5077 14124 5082
rect 14124 5077 14127 5082
rect 14165 5077 14192 5082
rect 14192 5077 14199 5082
rect 14237 5077 14260 5082
rect 14260 5077 14271 5082
rect 14309 5077 14328 5082
rect 14328 5077 14343 5082
rect 14381 5077 14396 5082
rect 14396 5077 14415 5082
rect 14453 5077 14464 5082
rect 14464 5077 14487 5082
rect 14525 5077 14532 5082
rect 14532 5077 14559 5082
rect 14597 5077 14600 5082
rect 14600 5077 14631 5082
rect 14669 5077 14702 5082
rect 14702 5077 14703 5082
rect 14741 5077 14770 5082
rect 14770 5077 14775 5082
rect 125 4849 231 5045
rect 269 5000 303 5029
rect 361 5001 395 5035
rect 434 5001 468 5035
rect 507 5001 541 5035
rect 580 5001 614 5035
rect 653 5001 687 5035
rect 726 5001 760 5035
rect 799 5001 833 5035
rect 872 5001 906 5035
rect 945 5001 979 5035
rect 1018 5001 1052 5035
rect 1091 5001 1125 5035
rect 1164 5001 1198 5035
rect 1237 5001 1271 5035
rect 1310 5001 1344 5035
rect 1383 5001 1417 5035
rect 1456 5001 1490 5035
rect 1529 5001 1563 5035
rect 1602 5001 1636 5035
rect 1675 5001 1709 5035
rect 1748 5001 1782 5035
rect 1821 5001 1855 5035
rect 1894 5001 1928 5035
rect 1967 5001 2001 5035
rect 2040 5001 2074 5035
rect 2113 5001 2147 5035
rect 2186 5001 2220 5035
rect 2259 5001 2293 5035
rect 2332 5001 2366 5035
rect 2405 5001 2439 5035
rect 2478 5001 2512 5035
rect 2551 5001 2585 5035
rect 2624 5001 2658 5035
rect 2697 5001 2731 5035
rect 2770 5001 2804 5035
rect 2843 5001 2877 5035
rect 2916 5001 2950 5035
rect 2989 5001 3023 5035
rect 3062 5001 3096 5035
rect 3135 5001 3169 5035
rect 3208 5001 3242 5035
rect 3281 5001 3315 5035
rect 3354 5001 3388 5035
rect 3427 5001 3461 5035
rect 3500 5001 3534 5035
rect 3573 5001 3607 5035
rect 3646 5001 3680 5035
rect 3719 5001 3753 5035
rect 3792 5001 3826 5035
rect 3865 5001 3899 5035
rect 3938 5001 3972 5035
rect 4011 5001 4045 5035
rect 4084 5001 4118 5035
rect 4157 5001 4191 5035
rect 4229 5001 4263 5035
rect 4301 5001 4335 5035
rect 4373 5001 4407 5035
rect 4445 5001 4479 5035
rect 4517 5001 4551 5035
rect 4589 5001 4623 5035
rect 4661 5001 4695 5035
rect 4733 5001 4767 5035
rect 4805 5001 4839 5035
rect 4877 5001 4911 5035
rect 4949 5001 4983 5035
rect 5021 5001 5055 5035
rect 5093 5001 5127 5035
rect 5165 5001 5199 5035
rect 5237 5001 5271 5035
rect 5309 5001 5343 5035
rect 5381 5001 5415 5035
rect 5453 5001 5487 5035
rect 5525 5001 5559 5035
rect 5597 5001 5631 5035
rect 5669 5001 5703 5035
rect 5741 5001 5775 5035
rect 5813 5001 5847 5035
rect 5885 5001 5919 5035
rect 5957 5001 5991 5035
rect 6029 5001 6063 5035
rect 6101 5001 6135 5035
rect 6173 5001 6207 5035
rect 6245 5001 6279 5035
rect 6317 5001 6351 5035
rect 6389 5001 6423 5035
rect 6461 5001 6495 5035
rect 6533 5001 6567 5035
rect 6605 5001 6639 5035
rect 6677 5001 6711 5035
rect 6749 5001 6783 5035
rect 6821 5001 6855 5035
rect 6893 5001 6927 5035
rect 6965 5001 6999 5035
rect 7037 5001 7071 5035
rect 7109 5001 7143 5035
rect 7181 5001 7215 5035
rect 7253 5001 7287 5035
rect 7325 5001 7359 5035
rect 7397 5001 7431 5035
rect 7469 5001 7503 5035
rect 7541 5001 7575 5035
rect 7613 5001 7647 5035
rect 7685 5001 7719 5035
rect 7757 5001 7791 5035
rect 7829 5001 7863 5035
rect 7901 5001 7935 5035
rect 7973 5001 8007 5035
rect 8045 5001 8079 5035
rect 8117 5001 8151 5035
rect 8189 5001 8223 5035
rect 8261 5001 8295 5035
rect 8333 5001 8367 5035
rect 8405 5001 8439 5035
rect 8477 5001 8511 5035
rect 8549 5001 8583 5035
rect 8621 5001 8655 5035
rect 8693 5001 8727 5035
rect 8765 5001 8799 5035
rect 8837 5001 8871 5035
rect 8909 5001 8943 5035
rect 8981 5001 9015 5035
rect 9053 5001 9087 5035
rect 9125 5001 9159 5035
rect 9197 5001 9231 5035
rect 9269 5001 9303 5035
rect 9341 5001 9375 5035
rect 9413 5001 9447 5035
rect 9485 5001 9519 5035
rect 9557 5001 9591 5035
rect 9629 5001 9663 5035
rect 9701 5001 9735 5035
rect 9773 5001 9807 5035
rect 9845 5001 9879 5035
rect 9917 5001 9951 5035
rect 9989 5001 10023 5035
rect 10061 5001 10095 5035
rect 10133 5001 10167 5035
rect 10205 5001 10239 5035
rect 10277 5001 10311 5035
rect 10349 5001 10383 5035
rect 10421 5001 10455 5035
rect 10493 5001 10527 5035
rect 10565 5001 10599 5035
rect 10637 5001 10671 5035
rect 10709 5001 10743 5035
rect 10781 5001 10815 5035
rect 10853 5001 10887 5035
rect 10925 5001 10959 5035
rect 10997 5001 11031 5035
rect 11069 5001 11103 5035
rect 11141 5001 11175 5035
rect 11213 5001 11247 5035
rect 11285 5001 11319 5035
rect 11357 5001 11391 5035
rect 11429 5001 11463 5035
rect 11501 5001 11535 5035
rect 11573 5001 11607 5035
rect 11645 5001 11679 5035
rect 11717 5001 11751 5035
rect 11789 5001 11823 5035
rect 11861 5001 11895 5035
rect 11933 5001 11967 5035
rect 12005 5001 12039 5035
rect 12077 5001 12111 5035
rect 12149 5001 12183 5035
rect 12221 5001 12255 5035
rect 12293 5001 12327 5035
rect 12365 5001 12399 5035
rect 12437 5001 12471 5035
rect 12509 5001 12543 5035
rect 12581 5001 12615 5035
rect 12653 5001 12687 5035
rect 12725 5001 12759 5035
rect 12797 5001 12831 5035
rect 12869 5001 12903 5035
rect 12941 5001 12975 5035
rect 13013 5001 13047 5035
rect 13085 5001 13119 5035
rect 13157 5001 13191 5035
rect 13229 5001 13263 5035
rect 13301 5001 13335 5035
rect 13373 5001 13407 5035
rect 13445 5001 13479 5035
rect 13517 5001 13551 5035
rect 13589 5001 13623 5035
rect 13661 5001 13695 5035
rect 13733 5001 13767 5035
rect 13805 5001 13839 5035
rect 13877 5001 13911 5035
rect 13949 5001 13983 5035
rect 14021 5001 14055 5035
rect 14093 5001 14127 5035
rect 14165 5001 14199 5035
rect 14237 5001 14271 5035
rect 14309 5001 14343 5035
rect 14381 5001 14415 5035
rect 14453 5001 14487 5035
rect 14525 5001 14559 5035
rect 14597 5001 14631 5035
rect 14669 5001 14703 5035
rect 14741 5001 14775 5035
rect 14907 5030 15013 5062
rect 14835 5000 15013 5030
rect 269 4995 286 5000
rect 286 4995 303 5000
rect 14835 4966 14838 5000
rect 14838 4966 14872 5000
rect 14872 4966 14906 5000
rect 14906 4966 15013 5000
rect 269 4922 303 4956
rect 361 4925 395 4959
rect 434 4925 468 4959
rect 507 4925 541 4959
rect 580 4925 614 4959
rect 653 4925 687 4959
rect 726 4925 760 4959
rect 799 4925 833 4959
rect 872 4925 906 4959
rect 945 4925 979 4959
rect 1018 4925 1052 4959
rect 1091 4925 1125 4959
rect 1164 4925 1198 4959
rect 1237 4925 1271 4959
rect 1310 4925 1344 4959
rect 1383 4925 1417 4959
rect 1456 4925 1490 4959
rect 1529 4925 1563 4959
rect 1602 4925 1636 4959
rect 1675 4925 1709 4959
rect 1748 4925 1782 4959
rect 1821 4925 1855 4959
rect 1894 4925 1928 4959
rect 1967 4925 2001 4959
rect 2040 4925 2074 4959
rect 2113 4925 2147 4959
rect 2186 4925 2220 4959
rect 2259 4925 2293 4959
rect 2332 4925 2366 4959
rect 2405 4925 2439 4959
rect 2478 4925 2512 4959
rect 2551 4925 2585 4959
rect 2624 4925 2658 4959
rect 2697 4925 2731 4959
rect 2770 4925 2804 4959
rect 2843 4925 2877 4959
rect 2916 4925 2950 4959
rect 2989 4925 3023 4959
rect 3062 4925 3096 4959
rect 3135 4925 3169 4959
rect 3208 4925 3242 4959
rect 3281 4925 3315 4959
rect 3354 4925 3388 4959
rect 3427 4925 3461 4959
rect 3500 4925 3534 4959
rect 3573 4925 3607 4959
rect 3646 4925 3680 4959
rect 3719 4925 3753 4959
rect 3792 4925 3826 4959
rect 3865 4925 3899 4959
rect 3938 4925 3972 4959
rect 4011 4925 4045 4959
rect 4084 4925 4118 4959
rect 4157 4925 4191 4959
rect 4229 4925 4263 4959
rect 4301 4925 4335 4959
rect 4373 4925 4407 4959
rect 4445 4925 4479 4959
rect 4517 4925 4551 4959
rect 4589 4925 4623 4959
rect 4661 4925 4695 4959
rect 4733 4925 4767 4959
rect 4805 4925 4839 4959
rect 4877 4925 4911 4959
rect 4949 4925 4983 4959
rect 5021 4925 5055 4959
rect 5093 4925 5127 4959
rect 5165 4925 5199 4959
rect 5237 4925 5271 4959
rect 5309 4925 5343 4959
rect 5381 4925 5415 4959
rect 5453 4925 5487 4959
rect 5525 4925 5559 4959
rect 5597 4925 5631 4959
rect 5669 4925 5703 4959
rect 5741 4925 5775 4959
rect 5813 4925 5847 4959
rect 5885 4925 5919 4959
rect 5957 4925 5991 4959
rect 6029 4925 6063 4959
rect 6101 4925 6135 4959
rect 6173 4925 6207 4959
rect 6245 4925 6279 4959
rect 6317 4925 6351 4959
rect 6389 4925 6423 4959
rect 6461 4925 6495 4959
rect 6533 4925 6567 4959
rect 6605 4925 6639 4959
rect 6677 4925 6711 4959
rect 6749 4925 6783 4959
rect 6821 4925 6855 4959
rect 6893 4925 6927 4959
rect 6965 4925 6999 4959
rect 7037 4925 7071 4959
rect 7109 4925 7143 4959
rect 7181 4925 7215 4959
rect 7253 4925 7287 4959
rect 7325 4925 7359 4959
rect 7397 4925 7431 4959
rect 7469 4925 7503 4959
rect 7541 4925 7575 4959
rect 7613 4925 7647 4959
rect 7685 4925 7719 4959
rect 7757 4925 7791 4959
rect 7829 4925 7863 4959
rect 7901 4925 7935 4959
rect 7973 4925 8007 4959
rect 8045 4925 8079 4959
rect 8117 4925 8151 4959
rect 8189 4925 8223 4959
rect 8261 4925 8295 4959
rect 8333 4925 8367 4959
rect 8405 4925 8439 4959
rect 8477 4925 8511 4959
rect 8549 4925 8583 4959
rect 8621 4925 8655 4959
rect 8693 4925 8727 4959
rect 8765 4925 8799 4959
rect 8837 4925 8871 4959
rect 8909 4925 8943 4959
rect 8981 4925 9015 4959
rect 9053 4925 9087 4959
rect 9125 4925 9159 4959
rect 9197 4925 9231 4959
rect 9269 4925 9303 4959
rect 9341 4925 9375 4959
rect 9413 4925 9447 4959
rect 9485 4925 9519 4959
rect 9557 4925 9591 4959
rect 9629 4925 9663 4959
rect 9701 4925 9735 4959
rect 9773 4925 9807 4959
rect 9845 4925 9879 4959
rect 9917 4925 9951 4959
rect 9989 4925 10023 4959
rect 10061 4925 10095 4959
rect 10133 4925 10167 4959
rect 10205 4925 10239 4959
rect 10277 4925 10311 4959
rect 10349 4925 10383 4959
rect 10421 4925 10455 4959
rect 10493 4925 10527 4959
rect 10565 4925 10599 4959
rect 10637 4925 10671 4959
rect 10709 4925 10743 4959
rect 10781 4925 10815 4959
rect 10853 4925 10887 4959
rect 10925 4925 10959 4959
rect 10997 4925 11031 4959
rect 11069 4925 11103 4959
rect 11141 4925 11175 4959
rect 11213 4925 11247 4959
rect 11285 4925 11319 4959
rect 11357 4925 11391 4959
rect 11429 4925 11463 4959
rect 11501 4925 11535 4959
rect 11573 4925 11607 4959
rect 11645 4925 11679 4959
rect 11717 4925 11751 4959
rect 11789 4925 11823 4959
rect 11861 4925 11895 4959
rect 11933 4925 11967 4959
rect 12005 4925 12039 4959
rect 12077 4925 12111 4959
rect 12149 4925 12183 4959
rect 12221 4925 12255 4959
rect 12293 4925 12327 4959
rect 12365 4925 12399 4959
rect 12437 4925 12471 4959
rect 12509 4925 12543 4959
rect 12581 4925 12615 4959
rect 12653 4925 12687 4959
rect 12725 4925 12759 4959
rect 12797 4925 12831 4959
rect 12869 4925 12903 4959
rect 12941 4925 12975 4959
rect 13013 4925 13047 4959
rect 13085 4925 13119 4959
rect 13157 4925 13191 4959
rect 13229 4925 13263 4959
rect 13301 4925 13335 4959
rect 13373 4925 13407 4959
rect 13445 4925 13479 4959
rect 13517 4925 13551 4959
rect 13589 4925 13623 4959
rect 13661 4925 13695 4959
rect 13733 4925 13767 4959
rect 13805 4925 13839 4959
rect 13877 4925 13911 4959
rect 13949 4925 13983 4959
rect 14021 4925 14055 4959
rect 14093 4925 14127 4959
rect 14165 4925 14199 4959
rect 14237 4925 14271 4959
rect 14309 4925 14343 4959
rect 14381 4925 14415 4959
rect 14453 4925 14487 4959
rect 14525 4925 14559 4959
rect 14597 4925 14631 4959
rect 14669 4925 14703 4959
rect 14741 4925 14775 4959
rect 14835 4918 15013 4966
rect 14835 4884 14838 4918
rect 14838 4884 14872 4918
rect 14872 4884 14906 4918
rect 14906 4884 15013 4918
rect 269 4849 303 4883
rect 125 599 193 4849
rect 193 599 231 4849
rect 269 4776 295 4810
rect 295 4776 303 4810
rect 269 4703 295 4737
rect 295 4703 303 4737
rect 269 4630 295 4664
rect 295 4630 303 4664
rect 14835 4849 15013 4884
rect 14835 4815 14840 4849
rect 14840 4815 14906 4849
rect 14906 4815 14940 4849
rect 14940 4815 15013 4849
rect 14835 4781 15013 4815
rect 14835 4747 14840 4781
rect 14840 4747 14906 4781
rect 14906 4747 14940 4781
rect 14940 4747 15013 4781
rect 14835 4713 15013 4747
rect 14835 4679 14840 4713
rect 14840 4679 14906 4713
rect 14906 4679 14940 4713
rect 14940 4679 15013 4713
rect 269 4557 295 4591
rect 295 4557 303 4591
rect 269 4484 295 4518
rect 295 4484 303 4518
rect 269 4411 295 4445
rect 295 4411 303 4445
rect 269 4338 295 4372
rect 295 4338 303 4372
rect 269 4265 295 4299
rect 295 4265 303 4299
rect 269 4192 295 4226
rect 295 4192 303 4226
rect 269 4119 295 4153
rect 295 4119 303 4153
rect 269 4046 295 4080
rect 295 4046 303 4080
rect 269 3973 295 4007
rect 295 3973 303 4007
rect 269 3900 295 3934
rect 295 3900 303 3934
rect 269 3827 295 3861
rect 295 3827 303 3861
rect 269 3754 295 3788
rect 295 3754 303 3788
rect 269 3681 295 3715
rect 295 3681 303 3715
rect 269 3608 295 3642
rect 295 3608 303 3642
rect 269 3535 295 3569
rect 295 3535 303 3569
rect 269 3462 295 3496
rect 295 3462 303 3496
rect 269 3389 295 3423
rect 295 3389 303 3423
rect 269 3316 295 3350
rect 295 3316 303 3350
rect 269 3243 295 3277
rect 295 3243 303 3277
rect 269 3170 295 3204
rect 295 3170 303 3204
rect 269 3097 295 3131
rect 295 3097 303 3131
rect 269 3024 295 3058
rect 295 3024 303 3058
rect 269 2951 295 2985
rect 295 2951 303 2985
rect 269 2878 295 2912
rect 295 2878 303 2912
rect 269 2805 295 2839
rect 295 2805 303 2839
rect 269 2732 295 2766
rect 295 2732 303 2766
rect 269 2659 295 2693
rect 295 2659 303 2693
rect 269 2586 295 2620
rect 295 2586 303 2620
rect 269 2513 295 2547
rect 295 2513 303 2547
rect 269 2440 295 2474
rect 295 2440 303 2474
rect 269 2367 295 2401
rect 295 2367 303 2401
rect 269 2294 295 2328
rect 295 2294 303 2328
rect 269 2221 295 2255
rect 295 2221 303 2255
rect 269 2148 295 2182
rect 295 2148 303 2182
rect 269 2075 295 2109
rect 295 2075 303 2109
rect 269 2002 295 2036
rect 295 2002 303 2036
rect 269 1929 295 1963
rect 295 1929 303 1963
rect 269 1856 295 1890
rect 295 1856 303 1890
rect 269 1783 295 1817
rect 295 1783 303 1817
rect 269 1710 295 1744
rect 295 1710 303 1744
rect 269 1637 295 1671
rect 295 1637 303 1671
rect 269 1564 295 1598
rect 295 1564 303 1598
rect 269 1491 295 1525
rect 295 1491 303 1525
rect 269 1418 295 1452
rect 295 1418 303 1452
rect 269 1345 295 1379
rect 295 1345 303 1379
rect 269 1272 295 1306
rect 295 1272 303 1306
rect 269 1199 295 1233
rect 295 1199 303 1233
rect 269 1125 295 1159
rect 295 1125 303 1159
rect 269 1051 295 1085
rect 295 1051 303 1085
rect 269 977 295 1011
rect 295 977 303 1011
rect 269 903 295 937
rect 295 903 303 937
rect 269 829 295 863
rect 295 829 303 863
rect 269 755 295 789
rect 295 755 303 789
rect 269 681 295 715
rect 295 681 303 715
rect 709 4570 10410 4606
rect 10410 4604 10445 4606
rect 10445 4604 10479 4606
rect 10479 4604 10514 4606
rect 10514 4604 10548 4606
rect 10548 4604 10583 4606
rect 10583 4604 10617 4606
rect 10617 4604 10652 4606
rect 10652 4604 10686 4606
rect 10686 4604 10721 4606
rect 10721 4604 10755 4606
rect 10755 4604 10790 4606
rect 10790 4604 10824 4606
rect 10824 4604 10859 4606
rect 10859 4604 10893 4606
rect 10893 4604 10928 4606
rect 10928 4604 10962 4606
rect 10962 4604 10997 4606
rect 10997 4604 11031 4606
rect 11031 4604 11066 4606
rect 11066 4604 11100 4606
rect 11100 4604 11135 4606
rect 11135 4604 11169 4606
rect 11169 4604 11204 4606
rect 11204 4604 11238 4606
rect 11238 4604 11273 4606
rect 11273 4604 11307 4606
rect 11307 4604 11342 4606
rect 11342 4604 11376 4606
rect 11376 4604 11411 4606
rect 11411 4604 11445 4606
rect 11445 4604 11480 4606
rect 11480 4604 11514 4606
rect 11514 4604 11549 4606
rect 11549 4604 11583 4606
rect 11583 4604 11618 4606
rect 11618 4604 11652 4606
rect 11652 4604 11687 4606
rect 11687 4604 11721 4606
rect 11721 4604 11756 4606
rect 11756 4604 11790 4606
rect 11790 4604 11825 4606
rect 11825 4604 11859 4606
rect 11859 4604 11894 4606
rect 11894 4604 11928 4606
rect 11928 4604 11963 4606
rect 11963 4604 11997 4606
rect 11997 4604 12032 4606
rect 12032 4604 12066 4606
rect 12066 4604 12101 4606
rect 12101 4604 12135 4606
rect 12135 4604 12170 4606
rect 12170 4604 12204 4606
rect 12204 4604 12239 4606
rect 12239 4604 12273 4606
rect 12273 4604 12308 4606
rect 12308 4604 12342 4606
rect 12342 4604 12377 4606
rect 12377 4604 12411 4606
rect 12411 4604 12446 4606
rect 12446 4604 12480 4606
rect 12480 4604 12515 4606
rect 12515 4604 12549 4606
rect 12549 4604 12584 4606
rect 12584 4604 12618 4606
rect 12618 4604 12653 4606
rect 12653 4604 12687 4606
rect 12687 4604 12722 4606
rect 12722 4604 12756 4606
rect 12756 4604 12791 4606
rect 12791 4604 12825 4606
rect 12825 4604 12860 4606
rect 12860 4604 12894 4606
rect 12894 4604 12929 4606
rect 12929 4604 12963 4606
rect 12963 4604 12998 4606
rect 12998 4604 13032 4606
rect 13032 4604 13067 4606
rect 13067 4604 13101 4606
rect 13101 4604 13136 4606
rect 13136 4604 13170 4606
rect 13170 4604 13205 4606
rect 13205 4604 13239 4606
rect 13239 4604 13274 4606
rect 13274 4604 13308 4606
rect 13308 4604 13343 4606
rect 13343 4604 13377 4606
rect 13377 4604 13412 4606
rect 13412 4604 13446 4606
rect 13446 4604 13481 4606
rect 13481 4604 13515 4606
rect 13515 4604 13550 4606
rect 13550 4604 13584 4606
rect 13584 4604 13619 4606
rect 13619 4604 13653 4606
rect 13653 4604 13688 4606
rect 13688 4604 13722 4606
rect 13722 4604 13757 4606
rect 13757 4604 13791 4606
rect 13791 4604 13826 4606
rect 13826 4604 13860 4606
rect 13860 4604 13895 4606
rect 13895 4604 13929 4606
rect 13929 4604 13964 4606
rect 13964 4604 13998 4606
rect 13998 4604 14033 4606
rect 14033 4604 14067 4606
rect 14067 4604 14102 4606
rect 14102 4604 14136 4606
rect 14136 4604 14171 4606
rect 14171 4604 14205 4606
rect 14205 4604 14207 4606
rect 14246 4604 14274 4606
rect 14274 4604 14280 4606
rect 14319 4604 14343 4606
rect 14343 4604 14353 4606
rect 14392 4604 14412 4606
rect 14412 4604 14426 4606
rect 10410 4570 14207 4604
rect 14246 4572 14280 4604
rect 14319 4572 14353 4604
rect 14392 4572 14426 4604
rect 709 4500 12363 4570
rect 12363 4536 12397 4570
rect 12397 4536 12431 4570
rect 12431 4536 12466 4570
rect 12466 4536 12500 4570
rect 12500 4536 12535 4570
rect 12535 4536 12569 4570
rect 12569 4536 12604 4570
rect 12604 4536 12638 4570
rect 12638 4536 12673 4570
rect 12673 4536 12707 4570
rect 12707 4536 12742 4570
rect 12742 4536 12776 4570
rect 12776 4536 12811 4570
rect 12811 4536 12845 4570
rect 12845 4536 12880 4570
rect 12880 4536 12914 4570
rect 12914 4536 12949 4570
rect 12949 4536 12983 4570
rect 12983 4536 13018 4570
rect 13018 4536 13052 4570
rect 13052 4536 13087 4570
rect 13087 4536 13121 4570
rect 13121 4536 13156 4570
rect 13156 4536 13190 4570
rect 13190 4536 13225 4570
rect 13225 4536 13259 4570
rect 13259 4536 13294 4570
rect 13294 4536 13328 4570
rect 13328 4536 13363 4570
rect 13363 4536 13397 4570
rect 13397 4536 13432 4570
rect 13432 4536 13466 4570
rect 13466 4536 13501 4570
rect 13501 4536 13535 4570
rect 13535 4536 13570 4570
rect 13570 4536 13604 4570
rect 13604 4536 13639 4570
rect 13639 4536 13673 4570
rect 13673 4536 13708 4570
rect 13708 4536 13742 4570
rect 13742 4536 13777 4570
rect 13777 4536 13811 4570
rect 13811 4536 13846 4570
rect 13846 4536 13880 4570
rect 13880 4536 13915 4570
rect 13915 4536 13949 4570
rect 13949 4536 13984 4570
rect 13984 4536 14018 4570
rect 14018 4536 14053 4570
rect 14053 4536 14087 4570
rect 14087 4536 14122 4570
rect 14122 4536 14156 4570
rect 14156 4536 14191 4570
rect 14191 4536 14207 4570
rect 12363 4502 14207 4536
rect 14246 4502 14280 4534
rect 14319 4502 14353 4534
rect 14392 4502 14426 4534
rect 12363 4500 12398 4502
rect 12398 4500 12432 4502
rect 12432 4500 12467 4502
rect 12467 4500 12501 4502
rect 12501 4500 12536 4502
rect 12536 4500 12570 4502
rect 12570 4500 12605 4502
rect 12605 4500 12639 4502
rect 12639 4500 12674 4502
rect 12674 4500 12708 4502
rect 12708 4500 12743 4502
rect 12743 4500 12777 4502
rect 12777 4500 12812 4502
rect 12812 4500 12846 4502
rect 12846 4500 12881 4502
rect 12881 4500 12915 4502
rect 12915 4500 12950 4502
rect 12950 4500 12984 4502
rect 12984 4500 13019 4502
rect 13019 4500 13053 4502
rect 13053 4500 13088 4502
rect 13088 4500 13122 4502
rect 13122 4500 13157 4502
rect 13157 4500 13191 4502
rect 13191 4500 13226 4502
rect 13226 4500 13260 4502
rect 13260 4500 13295 4502
rect 13295 4500 13329 4502
rect 13329 4500 13364 4502
rect 13364 4500 13398 4502
rect 13398 4500 13433 4502
rect 13433 4500 13467 4502
rect 13467 4500 13502 4502
rect 13502 4500 13536 4502
rect 13536 4500 13571 4502
rect 13571 4500 13605 4502
rect 13605 4500 13640 4502
rect 13640 4500 13674 4502
rect 13674 4500 13709 4502
rect 13709 4500 13743 4502
rect 13743 4500 13778 4502
rect 13778 4500 13812 4502
rect 13812 4500 13847 4502
rect 13847 4500 13881 4502
rect 13881 4500 13916 4502
rect 13916 4500 13950 4502
rect 13950 4500 13985 4502
rect 13985 4500 14019 4502
rect 14019 4500 14054 4502
rect 14054 4500 14088 4502
rect 14088 4500 14123 4502
rect 14123 4500 14157 4502
rect 14157 4500 14192 4502
rect 14192 4500 14207 4502
rect 14246 4500 14261 4502
rect 14261 4500 14280 4502
rect 14319 4500 14330 4502
rect 14330 4500 14353 4502
rect 14392 4500 14399 4502
rect 14399 4500 14426 4502
rect 674 4445 708 4456
rect 529 4409 563 4426
rect 529 4392 531 4409
rect 531 4392 563 4409
rect 601 4395 633 4426
rect 633 4395 635 4426
rect 601 4392 635 4395
rect 529 4339 563 4351
rect 529 4317 531 4339
rect 531 4317 563 4339
rect 601 4322 633 4351
rect 633 4322 635 4351
rect 601 4317 635 4322
rect 529 4269 563 4276
rect 529 4242 531 4269
rect 531 4242 563 4269
rect 601 4249 633 4276
rect 633 4249 635 4276
rect 601 4242 635 4249
rect 529 4199 563 4201
rect 529 4167 531 4199
rect 531 4167 563 4199
rect 601 4177 633 4201
rect 633 4177 635 4201
rect 601 4167 635 4177
rect 529 4095 531 4126
rect 531 4095 563 4126
rect 601 4105 633 4126
rect 633 4105 635 4126
rect 529 4092 563 4095
rect 601 4092 635 4105
rect 674 4082 780 4445
rect 14356 4398 14390 4432
rect 14428 4426 14462 4456
rect 14356 4325 14390 4359
rect 529 4025 531 4052
rect 531 4025 563 4052
rect 601 4033 633 4052
rect 633 4033 635 4052
rect 674 4048 745 4082
rect 745 4048 779 4082
rect 779 4048 780 4082
rect 529 4018 563 4025
rect 601 4018 635 4033
rect 674 4014 780 4048
rect 529 3955 531 3978
rect 531 3955 563 3978
rect 601 3961 633 3978
rect 633 3961 635 3978
rect 674 3980 745 4014
rect 745 3980 779 4014
rect 779 3980 780 4014
rect 529 3944 563 3955
rect 601 3944 635 3961
rect 674 3946 780 3980
rect 529 3886 531 3904
rect 531 3886 563 3904
rect 601 3889 633 3904
rect 633 3889 635 3904
rect 674 3912 745 3946
rect 745 3912 779 3946
rect 779 3912 780 3946
rect 529 3870 563 3886
rect 601 3870 635 3889
rect 674 3878 780 3912
rect 674 3844 745 3878
rect 745 3844 779 3878
rect 779 3844 780 3878
rect 674 3810 780 3844
rect 529 3760 563 3794
rect 601 3760 635 3794
rect 674 3776 745 3810
rect 745 3776 779 3810
rect 779 3776 780 3810
rect 529 3715 531 3720
rect 531 3715 563 3720
rect 601 3715 633 3720
rect 633 3715 635 3720
rect 674 3742 780 3776
rect 529 3686 563 3715
rect 601 3686 635 3715
rect 674 3708 745 3742
rect 745 3708 779 3742
rect 779 3708 780 3742
rect 674 3674 780 3708
rect 529 3612 563 3646
rect 601 3612 635 3646
rect 674 3640 745 3674
rect 745 3640 779 3674
rect 779 3640 780 3674
rect 674 3606 780 3640
rect 674 3572 745 3606
rect 745 3572 779 3606
rect 779 3572 780 3606
rect 529 3542 563 3572
rect 601 3542 635 3572
rect 529 3538 531 3542
rect 531 3538 563 3542
rect 601 3538 633 3542
rect 633 3538 635 3542
rect 674 3538 780 3572
rect 674 3504 745 3538
rect 745 3504 779 3538
rect 779 3504 780 3538
rect 529 3473 563 3498
rect 601 3473 635 3498
rect 529 3464 531 3473
rect 531 3464 563 3473
rect 601 3464 633 3473
rect 633 3464 635 3473
rect 674 3470 780 3504
rect 674 3436 745 3470
rect 745 3436 779 3470
rect 779 3436 780 3470
rect 529 3404 563 3424
rect 601 3404 635 3424
rect 529 3390 531 3404
rect 531 3390 563 3404
rect 601 3390 633 3404
rect 633 3390 635 3404
rect 674 3402 780 3436
rect 674 3368 745 3402
rect 745 3368 779 3402
rect 779 3368 780 3402
rect 529 3335 563 3350
rect 601 3335 635 3350
rect 529 3316 531 3335
rect 531 3316 563 3335
rect 601 3316 633 3335
rect 633 3316 635 3335
rect 674 3334 780 3368
rect 674 3300 745 3334
rect 745 3300 779 3334
rect 779 3300 780 3334
rect 529 3266 563 3276
rect 601 3266 635 3276
rect 674 3266 780 3300
rect 529 3242 531 3266
rect 531 3242 563 3266
rect 601 3242 633 3266
rect 633 3242 635 3266
rect 674 3232 745 3266
rect 745 3232 779 3266
rect 779 3232 780 3266
rect 529 3197 563 3202
rect 601 3197 635 3202
rect 674 3198 780 3232
rect 529 3168 531 3197
rect 531 3168 563 3197
rect 601 3168 633 3197
rect 633 3168 635 3197
rect 674 3164 745 3198
rect 745 3164 779 3198
rect 779 3164 780 3198
rect 529 3094 531 3128
rect 531 3094 563 3128
rect 601 3094 633 3128
rect 633 3094 635 3128
rect 529 3025 531 3054
rect 531 3025 563 3054
rect 601 3025 633 3054
rect 633 3025 635 3054
rect 529 3020 563 3025
rect 601 3020 635 3025
rect 529 2956 531 2980
rect 531 2956 563 2980
rect 601 2956 633 2980
rect 633 2956 635 2980
rect 529 2946 563 2956
rect 601 2946 635 2956
rect 529 2887 531 2906
rect 531 2887 563 2906
rect 601 2887 633 2906
rect 633 2887 635 2906
rect 529 2872 563 2887
rect 601 2872 635 2887
rect 529 2818 531 2832
rect 531 2818 563 2832
rect 601 2818 633 2832
rect 633 2818 635 2832
rect 529 2798 563 2818
rect 601 2798 635 2818
rect 529 2749 531 2758
rect 531 2749 563 2758
rect 601 2749 633 2758
rect 633 2749 635 2758
rect 529 2724 563 2749
rect 601 2724 635 2749
rect 529 2680 531 2684
rect 531 2680 563 2684
rect 601 2680 633 2684
rect 633 2680 635 2684
rect 529 2650 563 2680
rect 601 2650 635 2680
rect 529 2576 563 2610
rect 601 2576 635 2610
rect 529 2507 563 2536
rect 601 2507 635 2536
rect 529 2502 531 2507
rect 531 2502 563 2507
rect 601 2502 633 2507
rect 633 2502 635 2507
rect 674 2482 780 3164
rect 529 2438 563 2462
rect 601 2438 635 2462
rect 674 2448 745 2482
rect 745 2448 779 2482
rect 779 2448 780 2482
rect 529 2428 531 2438
rect 531 2428 563 2438
rect 601 2428 633 2438
rect 633 2428 635 2438
rect 674 2414 780 2448
rect 529 2369 563 2389
rect 601 2369 635 2389
rect 674 2380 745 2414
rect 745 2380 779 2414
rect 779 2380 780 2414
rect 529 2355 531 2369
rect 531 2355 563 2369
rect 601 2355 633 2369
rect 633 2355 635 2369
rect 674 2346 780 2380
rect 529 2300 563 2316
rect 601 2300 635 2316
rect 674 2312 745 2346
rect 745 2312 779 2346
rect 779 2312 780 2346
rect 529 2282 531 2300
rect 531 2282 563 2300
rect 601 2282 633 2300
rect 633 2282 635 2300
rect 674 2278 780 2312
rect 674 2244 745 2278
rect 745 2244 779 2278
rect 779 2244 780 2278
rect 529 2231 563 2243
rect 601 2231 635 2243
rect 529 2209 531 2231
rect 531 2209 563 2231
rect 601 2209 633 2231
rect 633 2209 635 2231
rect 674 2210 780 2244
rect 674 2176 745 2210
rect 745 2176 779 2210
rect 779 2176 780 2210
rect 529 2163 563 2170
rect 529 2136 531 2163
rect 531 2136 563 2163
rect 601 2162 635 2170
rect 601 2136 633 2162
rect 633 2136 635 2162
rect 674 2142 780 2176
rect 674 2108 745 2142
rect 745 2108 779 2142
rect 779 2108 780 2142
rect 529 2095 563 2097
rect 529 2063 531 2095
rect 531 2063 563 2095
rect 601 2093 635 2097
rect 601 2063 633 2093
rect 633 2063 635 2093
rect 674 2074 780 2108
rect 674 2040 745 2074
rect 745 2040 779 2074
rect 779 2040 780 2074
rect 529 1993 531 2024
rect 531 1993 563 2024
rect 529 1990 563 1993
rect 601 1990 633 2024
rect 633 1990 635 2024
rect 674 2006 780 2040
rect 674 1972 745 2006
rect 745 1972 779 2006
rect 779 1972 780 2006
rect 529 1925 531 1951
rect 531 1925 563 1951
rect 529 1917 563 1925
rect 601 1921 633 1951
rect 633 1921 635 1951
rect 674 1938 780 1972
rect 601 1917 635 1921
rect 674 1904 745 1938
rect 745 1904 779 1938
rect 779 1904 780 1938
rect 529 1857 531 1878
rect 531 1857 563 1878
rect 529 1844 563 1857
rect 601 1852 633 1878
rect 633 1852 635 1878
rect 674 1870 780 1904
rect 601 1844 635 1852
rect 674 1836 745 1870
rect 745 1836 779 1870
rect 779 1836 780 1870
rect 529 1789 531 1805
rect 531 1789 563 1805
rect 529 1771 563 1789
rect 601 1783 633 1805
rect 633 1783 635 1805
rect 674 1802 780 1836
rect 601 1771 635 1783
rect 674 1768 745 1802
rect 745 1768 779 1802
rect 779 1768 780 1802
rect 529 1721 531 1732
rect 531 1721 563 1732
rect 529 1698 563 1721
rect 601 1714 633 1732
rect 633 1714 635 1732
rect 674 1734 780 1768
rect 601 1698 635 1714
rect 674 1700 745 1734
rect 745 1700 779 1734
rect 779 1700 780 1734
rect 529 1653 531 1659
rect 531 1653 563 1659
rect 529 1625 563 1653
rect 601 1645 633 1659
rect 633 1645 635 1659
rect 674 1666 780 1700
rect 601 1625 635 1645
rect 674 1632 745 1666
rect 745 1632 779 1666
rect 779 1632 780 1666
rect 529 1585 531 1586
rect 531 1585 563 1586
rect 529 1552 563 1585
rect 601 1576 633 1586
rect 633 1576 635 1586
rect 674 1598 780 1632
rect 601 1552 635 1576
rect 674 1564 745 1598
rect 745 1564 779 1598
rect 779 1564 780 1598
rect 529 1483 563 1513
rect 601 1507 633 1513
rect 633 1507 635 1513
rect 529 1479 531 1483
rect 531 1479 563 1483
rect 601 1479 635 1507
rect 529 1415 563 1440
rect 601 1438 633 1440
rect 633 1438 635 1440
rect 529 1406 531 1415
rect 531 1406 563 1415
rect 601 1406 635 1438
rect 529 1347 563 1367
rect 529 1333 531 1347
rect 531 1333 563 1347
rect 601 1334 635 1367
rect 601 1333 633 1334
rect 633 1333 635 1334
rect 529 1279 563 1294
rect 529 1260 531 1279
rect 531 1260 563 1279
rect 601 1265 635 1294
rect 601 1260 633 1265
rect 633 1260 635 1265
rect 529 1211 563 1221
rect 529 1187 531 1211
rect 531 1187 563 1211
rect 601 1196 635 1221
rect 601 1187 633 1196
rect 633 1187 635 1196
rect 529 1143 563 1148
rect 529 1114 531 1143
rect 531 1114 563 1143
rect 601 1127 635 1148
rect 601 1114 633 1127
rect 633 1114 635 1127
rect 529 1041 531 1075
rect 531 1041 563 1075
rect 601 1058 635 1075
rect 601 1041 633 1058
rect 633 1041 635 1058
rect 529 973 531 1002
rect 531 973 563 1002
rect 601 989 635 1002
rect 529 968 563 973
rect 601 968 633 989
rect 633 968 635 989
rect 529 920 531 929
rect 531 920 563 929
rect 601 920 635 929
rect 529 895 563 920
rect 601 895 635 920
rect 674 894 780 1564
rect 1067 4064 1101 4098
rect 1139 4064 1173 4098
rect 1211 4064 1245 4098
rect 1067 3991 1101 4025
rect 1139 3991 1173 4025
rect 1211 3991 1245 4025
rect 1067 3918 1101 3952
rect 1139 3918 1173 3952
rect 1211 3918 1245 3952
rect 1067 3845 1101 3879
rect 1139 3845 1173 3879
rect 1211 3845 1245 3879
rect 1067 3772 1101 3806
rect 1139 3772 1173 3806
rect 1211 3772 1245 3806
rect 1067 3699 1101 3733
rect 1139 3699 1173 3733
rect 1211 3699 1245 3733
rect 1067 3626 1101 3660
rect 1139 3626 1173 3660
rect 1211 3626 1245 3660
rect 1067 3553 1101 3587
rect 1139 3553 1173 3587
rect 1211 3553 1245 3587
rect 1067 3480 1101 3514
rect 1139 3480 1173 3514
rect 1211 3480 1245 3514
rect 1067 3407 1101 3441
rect 1139 3407 1173 3441
rect 1211 3407 1245 3441
rect 1067 3334 1101 3368
rect 1139 3334 1173 3368
rect 1211 3334 1245 3368
rect 1067 3261 1101 3295
rect 1139 3261 1173 3295
rect 1211 3261 1245 3295
rect 1067 3188 1101 3222
rect 1139 3188 1173 3222
rect 1211 3188 1245 3222
rect 1067 3115 1101 3149
rect 1139 3115 1173 3149
rect 1211 3115 1245 3149
rect 1067 3042 1101 3076
rect 1139 3042 1173 3076
rect 1211 3042 1245 3076
rect 1067 2969 1101 3003
rect 1139 2969 1173 3003
rect 1211 2969 1245 3003
rect 1067 2896 1101 2930
rect 1139 2896 1173 2930
rect 1211 2896 1245 2930
rect 1067 2823 1101 2857
rect 1139 2823 1173 2857
rect 1211 2823 1245 2857
rect 1067 2750 1101 2784
rect 1139 2750 1173 2784
rect 1211 2750 1245 2784
rect 1067 2677 1101 2711
rect 1139 2677 1173 2711
rect 1211 2677 1245 2711
rect 1067 2604 1101 2638
rect 1139 2604 1173 2638
rect 1211 2604 1245 2638
rect 1067 2531 1101 2565
rect 1139 2531 1173 2565
rect 1211 2531 1245 2565
rect 1067 2458 1101 2492
rect 1139 2458 1173 2492
rect 1211 2458 1245 2492
rect 1067 2385 1101 2419
rect 1139 2385 1173 2419
rect 1211 2385 1245 2419
rect 1067 2312 1101 2346
rect 1139 2312 1173 2346
rect 1211 2312 1245 2346
rect 1067 2239 1101 2273
rect 1139 2239 1173 2273
rect 1211 2239 1245 2273
rect 1067 2166 1101 2200
rect 1139 2166 1173 2200
rect 1211 2166 1245 2200
rect 1067 2092 1101 2126
rect 1139 2092 1173 2126
rect 1211 2092 1245 2126
rect 1067 2018 1101 2052
rect 1139 2018 1173 2052
rect 1211 2018 1245 2052
rect 1067 1944 1101 1978
rect 1139 1944 1173 1978
rect 1211 1944 1245 1978
rect 1067 1870 1101 1904
rect 1139 1870 1173 1904
rect 1211 1870 1245 1904
rect 1067 1796 1101 1830
rect 1139 1796 1173 1830
rect 1211 1796 1245 1830
rect 1067 1722 1101 1756
rect 1139 1722 1173 1756
rect 1211 1722 1245 1756
rect 1067 1648 1101 1682
rect 1139 1648 1173 1682
rect 1211 1648 1245 1682
rect 1067 1574 1101 1608
rect 1139 1574 1173 1608
rect 1211 1574 1245 1608
rect 924 1216 958 1250
rect 924 1144 958 1178
rect 1635 4092 1669 4118
rect 1563 4082 1741 4092
rect 1563 4048 1567 4082
rect 1567 4048 1635 4082
rect 1635 4048 1669 4082
rect 1669 4048 1737 4082
rect 1737 4048 1741 4082
rect 1563 4014 1741 4048
rect 1563 3980 1567 4014
rect 1567 3980 1635 4014
rect 1635 3980 1669 4014
rect 1669 3980 1737 4014
rect 1737 3980 1741 4014
rect 1563 3946 1741 3980
rect 1563 3912 1567 3946
rect 1567 3912 1635 3946
rect 1635 3912 1669 3946
rect 1669 3912 1737 3946
rect 1737 3912 1741 3946
rect 1563 3878 1741 3912
rect 1563 3844 1567 3878
rect 1567 3844 1635 3878
rect 1635 3844 1669 3878
rect 1669 3844 1737 3878
rect 1737 3844 1741 3878
rect 1563 3810 1741 3844
rect 1563 3776 1567 3810
rect 1567 3776 1635 3810
rect 1635 3776 1669 3810
rect 1669 3776 1737 3810
rect 1737 3776 1741 3810
rect 1563 3742 1741 3776
rect 1563 3708 1567 3742
rect 1567 3708 1635 3742
rect 1635 3708 1669 3742
rect 1669 3708 1737 3742
rect 1737 3708 1741 3742
rect 1563 3674 1741 3708
rect 1563 3640 1567 3674
rect 1567 3640 1635 3674
rect 1635 3640 1669 3674
rect 1669 3640 1737 3674
rect 1737 3640 1741 3674
rect 1563 3606 1741 3640
rect 1563 3572 1567 3606
rect 1567 3572 1635 3606
rect 1635 3572 1669 3606
rect 1669 3572 1737 3606
rect 1737 3572 1741 3606
rect 1563 3538 1741 3572
rect 1563 3504 1567 3538
rect 1567 3504 1635 3538
rect 1635 3504 1669 3538
rect 1669 3504 1737 3538
rect 1737 3504 1741 3538
rect 1563 3470 1741 3504
rect 1563 3436 1567 3470
rect 1567 3436 1635 3470
rect 1635 3436 1669 3470
rect 1669 3436 1737 3470
rect 1737 3436 1741 3470
rect 1563 3402 1741 3436
rect 1563 3368 1567 3402
rect 1567 3368 1635 3402
rect 1635 3368 1669 3402
rect 1669 3368 1737 3402
rect 1737 3368 1741 3402
rect 1563 3334 1741 3368
rect 1563 3300 1567 3334
rect 1567 3300 1635 3334
rect 1635 3300 1669 3334
rect 1669 3300 1737 3334
rect 1737 3300 1741 3334
rect 1563 3266 1741 3300
rect 1563 3232 1567 3266
rect 1567 3232 1635 3266
rect 1635 3232 1669 3266
rect 1669 3232 1737 3266
rect 1737 3232 1741 3266
rect 1563 3198 1741 3232
rect 1563 3194 1567 3198
rect 1567 3194 1635 3198
rect 1635 3194 1669 3198
rect 1669 3194 1737 3198
rect 1737 3194 1741 3198
rect 1635 3164 1669 3182
rect 1635 3148 1669 3164
rect 1563 3074 1597 3108
rect 1635 3074 1669 3108
rect 1707 3074 1741 3108
rect 1563 2994 1597 3028
rect 1635 2994 1669 3028
rect 1707 2994 1741 3028
rect 1563 2914 1597 2948
rect 1635 2914 1669 2948
rect 1707 2914 1741 2948
rect 1563 2834 1597 2868
rect 1635 2834 1669 2868
rect 1707 2834 1741 2868
rect 1563 2754 1597 2788
rect 1635 2754 1669 2788
rect 1707 2754 1741 2788
rect 1563 2674 1597 2708
rect 1635 2674 1669 2708
rect 1707 2674 1741 2708
rect 1563 2594 1597 2628
rect 1635 2594 1669 2628
rect 1707 2594 1741 2628
rect 1635 2540 1669 2556
rect 1635 2522 1669 2540
rect 1563 2506 1567 2518
rect 1567 2506 1635 2518
rect 1635 2506 1669 2518
rect 1669 2506 1737 2518
rect 1737 2506 1741 2518
rect 1563 2472 1741 2506
rect 1563 2438 1567 2472
rect 1567 2438 1635 2472
rect 1635 2438 1669 2472
rect 1669 2438 1737 2472
rect 1737 2438 1741 2472
rect 1563 2404 1741 2438
rect 1563 2370 1567 2404
rect 1567 2370 1635 2404
rect 1635 2370 1669 2404
rect 1669 2370 1737 2404
rect 1737 2370 1741 2404
rect 1563 2336 1741 2370
rect 1563 2302 1567 2336
rect 1567 2302 1635 2336
rect 1635 2302 1669 2336
rect 1669 2302 1737 2336
rect 1737 2302 1741 2336
rect 1563 2268 1741 2302
rect 1563 2234 1567 2268
rect 1567 2234 1635 2268
rect 1635 2234 1669 2268
rect 1669 2234 1737 2268
rect 1737 2234 1741 2268
rect 1563 2200 1741 2234
rect 1563 2166 1567 2200
rect 1567 2166 1635 2200
rect 1635 2166 1669 2200
rect 1669 2166 1737 2200
rect 1737 2166 1741 2200
rect 1563 2132 1741 2166
rect 1563 2098 1567 2132
rect 1567 2098 1635 2132
rect 1635 2098 1669 2132
rect 1669 2098 1737 2132
rect 1737 2098 1741 2132
rect 1563 2064 1741 2098
rect 1563 2030 1567 2064
rect 1567 2030 1635 2064
rect 1635 2030 1669 2064
rect 1669 2030 1737 2064
rect 1737 2030 1741 2064
rect 1563 1996 1741 2030
rect 1563 1962 1567 1996
rect 1567 1962 1635 1996
rect 1635 1962 1669 1996
rect 1669 1962 1737 1996
rect 1737 1962 1741 1996
rect 1563 1928 1741 1962
rect 1563 1894 1567 1928
rect 1567 1894 1635 1928
rect 1635 1894 1669 1928
rect 1669 1894 1737 1928
rect 1737 1894 1741 1928
rect 1563 1860 1741 1894
rect 1563 1826 1567 1860
rect 1567 1826 1635 1860
rect 1635 1826 1669 1860
rect 1669 1826 1737 1860
rect 1737 1826 1741 1860
rect 1563 1792 1741 1826
rect 1563 1758 1567 1792
rect 1567 1758 1635 1792
rect 1635 1758 1669 1792
rect 1669 1758 1737 1792
rect 1737 1758 1741 1792
rect 1563 1724 1741 1758
rect 1563 1690 1567 1724
rect 1567 1690 1635 1724
rect 1635 1690 1669 1724
rect 1669 1690 1737 1724
rect 1737 1690 1741 1724
rect 1563 1656 1741 1690
rect 1563 1622 1567 1656
rect 1567 1622 1635 1656
rect 1635 1622 1669 1656
rect 1669 1622 1737 1656
rect 1737 1622 1741 1656
rect 1563 1620 1741 1622
rect 1635 1586 1669 1620
rect 1318 1144 1424 1250
rect 2059 4064 2093 4098
rect 2131 4064 2165 4098
rect 2203 4064 2237 4098
rect 2059 3991 2093 4025
rect 2131 3991 2165 4025
rect 2203 3991 2237 4025
rect 2059 3918 2093 3952
rect 2131 3918 2165 3952
rect 2203 3918 2237 3952
rect 2059 3845 2093 3879
rect 2131 3845 2165 3879
rect 2203 3845 2237 3879
rect 2059 3772 2093 3806
rect 2131 3772 2165 3806
rect 2203 3772 2237 3806
rect 2059 3699 2093 3733
rect 2131 3699 2165 3733
rect 2203 3699 2237 3733
rect 2059 3626 2093 3660
rect 2131 3626 2165 3660
rect 2203 3626 2237 3660
rect 2059 3553 2093 3587
rect 2131 3553 2165 3587
rect 2203 3553 2237 3587
rect 2059 3480 2093 3514
rect 2131 3480 2165 3514
rect 2203 3480 2237 3514
rect 2059 3407 2093 3441
rect 2131 3407 2165 3441
rect 2203 3407 2237 3441
rect 2059 3334 2093 3368
rect 2131 3334 2165 3368
rect 2203 3334 2237 3368
rect 2059 3261 2093 3295
rect 2131 3261 2165 3295
rect 2203 3261 2237 3295
rect 2059 3188 2093 3222
rect 2131 3188 2165 3222
rect 2203 3188 2237 3222
rect 2059 3115 2093 3149
rect 2131 3115 2165 3149
rect 2203 3115 2237 3149
rect 2059 3042 2093 3076
rect 2131 3042 2165 3076
rect 2203 3042 2237 3076
rect 2059 2969 2093 3003
rect 2131 2969 2165 3003
rect 2203 2969 2237 3003
rect 2059 2896 2093 2930
rect 2131 2896 2165 2930
rect 2203 2896 2237 2930
rect 2059 2823 2093 2857
rect 2131 2823 2165 2857
rect 2203 2823 2237 2857
rect 2059 2750 2093 2784
rect 2131 2750 2165 2784
rect 2203 2750 2237 2784
rect 2059 2677 2093 2711
rect 2131 2677 2165 2711
rect 2203 2677 2237 2711
rect 2059 2604 2093 2638
rect 2131 2604 2165 2638
rect 2203 2604 2237 2638
rect 2059 2531 2093 2565
rect 2131 2531 2165 2565
rect 2203 2531 2237 2565
rect 2059 2458 2093 2492
rect 2131 2458 2165 2492
rect 2203 2458 2237 2492
rect 2059 2385 2093 2419
rect 2131 2385 2165 2419
rect 2203 2385 2237 2419
rect 2059 2312 2093 2346
rect 2131 2312 2165 2346
rect 2203 2312 2237 2346
rect 2059 2239 2093 2273
rect 2131 2239 2165 2273
rect 2203 2239 2237 2273
rect 2059 2166 2093 2200
rect 2131 2166 2165 2200
rect 2203 2166 2237 2200
rect 2059 2092 2093 2126
rect 2131 2092 2165 2126
rect 2203 2092 2237 2126
rect 2059 2018 2093 2052
rect 2131 2018 2165 2052
rect 2203 2018 2237 2052
rect 2059 1944 2093 1978
rect 2131 1944 2165 1978
rect 2203 1944 2237 1978
rect 2059 1870 2093 1904
rect 2131 1870 2165 1904
rect 2203 1870 2237 1904
rect 2059 1796 2093 1830
rect 2131 1796 2165 1830
rect 2203 1796 2237 1830
rect 2059 1722 2093 1756
rect 2131 1722 2165 1756
rect 2203 1722 2237 1756
rect 2059 1648 2093 1682
rect 2131 1648 2165 1682
rect 2203 1648 2237 1682
rect 2059 1574 2093 1608
rect 2131 1574 2165 1608
rect 2203 1574 2237 1608
rect 1880 1144 1986 1250
rect 2627 4092 2661 4118
rect 2555 4082 2733 4092
rect 2555 4048 2559 4082
rect 2559 4048 2627 4082
rect 2627 4048 2661 4082
rect 2661 4048 2729 4082
rect 2729 4048 2733 4082
rect 2555 4014 2733 4048
rect 2555 3980 2559 4014
rect 2559 3980 2627 4014
rect 2627 3980 2661 4014
rect 2661 3980 2729 4014
rect 2729 3980 2733 4014
rect 2555 3946 2733 3980
rect 2555 3912 2559 3946
rect 2559 3912 2627 3946
rect 2627 3912 2661 3946
rect 2661 3912 2729 3946
rect 2729 3912 2733 3946
rect 2555 3878 2733 3912
rect 2555 3844 2559 3878
rect 2559 3844 2627 3878
rect 2627 3844 2661 3878
rect 2661 3844 2729 3878
rect 2729 3844 2733 3878
rect 2555 3810 2733 3844
rect 2555 3776 2559 3810
rect 2559 3776 2627 3810
rect 2627 3776 2661 3810
rect 2661 3776 2729 3810
rect 2729 3776 2733 3810
rect 2555 3742 2733 3776
rect 2555 3708 2559 3742
rect 2559 3708 2627 3742
rect 2627 3708 2661 3742
rect 2661 3708 2729 3742
rect 2729 3708 2733 3742
rect 2555 3674 2733 3708
rect 2555 3640 2559 3674
rect 2559 3640 2627 3674
rect 2627 3640 2661 3674
rect 2661 3640 2729 3674
rect 2729 3640 2733 3674
rect 2555 3606 2733 3640
rect 2555 3572 2559 3606
rect 2559 3572 2627 3606
rect 2627 3572 2661 3606
rect 2661 3572 2729 3606
rect 2729 3572 2733 3606
rect 2555 3538 2733 3572
rect 2555 3504 2559 3538
rect 2559 3504 2627 3538
rect 2627 3504 2661 3538
rect 2661 3504 2729 3538
rect 2729 3504 2733 3538
rect 2555 3470 2733 3504
rect 2555 3436 2559 3470
rect 2559 3436 2627 3470
rect 2627 3436 2661 3470
rect 2661 3436 2729 3470
rect 2729 3436 2733 3470
rect 2555 3402 2733 3436
rect 2555 3368 2559 3402
rect 2559 3368 2627 3402
rect 2627 3368 2661 3402
rect 2661 3368 2729 3402
rect 2729 3368 2733 3402
rect 2555 3334 2733 3368
rect 2555 3300 2559 3334
rect 2559 3300 2627 3334
rect 2627 3300 2661 3334
rect 2661 3300 2729 3334
rect 2729 3300 2733 3334
rect 2555 3266 2733 3300
rect 2555 3232 2559 3266
rect 2559 3232 2627 3266
rect 2627 3232 2661 3266
rect 2661 3232 2729 3266
rect 2729 3232 2733 3266
rect 2555 3198 2733 3232
rect 2555 3194 2559 3198
rect 2559 3194 2627 3198
rect 2627 3194 2661 3198
rect 2661 3194 2729 3198
rect 2729 3194 2733 3198
rect 2627 3164 2661 3182
rect 2627 3148 2661 3164
rect 2555 3074 2589 3108
rect 2627 3074 2661 3108
rect 2699 3074 2733 3108
rect 2555 2994 2589 3028
rect 2627 2994 2661 3028
rect 2699 2994 2733 3028
rect 2555 2914 2589 2948
rect 2627 2914 2661 2948
rect 2699 2914 2733 2948
rect 2555 2834 2589 2868
rect 2627 2834 2661 2868
rect 2699 2834 2733 2868
rect 2555 2754 2589 2788
rect 2627 2754 2661 2788
rect 2699 2754 2733 2788
rect 2555 2674 2589 2708
rect 2627 2674 2661 2708
rect 2699 2674 2733 2708
rect 2555 2594 2589 2628
rect 2627 2594 2661 2628
rect 2699 2594 2733 2628
rect 2627 2540 2661 2556
rect 2627 2522 2661 2540
rect 2555 2506 2559 2518
rect 2559 2506 2627 2518
rect 2627 2506 2661 2518
rect 2661 2506 2729 2518
rect 2729 2506 2733 2518
rect 2555 2472 2733 2506
rect 2555 2438 2559 2472
rect 2559 2438 2627 2472
rect 2627 2438 2661 2472
rect 2661 2438 2729 2472
rect 2729 2438 2733 2472
rect 2555 2404 2733 2438
rect 2555 2370 2559 2404
rect 2559 2370 2627 2404
rect 2627 2370 2661 2404
rect 2661 2370 2729 2404
rect 2729 2370 2733 2404
rect 2555 2336 2733 2370
rect 2555 2302 2559 2336
rect 2559 2302 2627 2336
rect 2627 2302 2661 2336
rect 2661 2302 2729 2336
rect 2729 2302 2733 2336
rect 2555 2268 2733 2302
rect 2555 2234 2559 2268
rect 2559 2234 2627 2268
rect 2627 2234 2661 2268
rect 2661 2234 2729 2268
rect 2729 2234 2733 2268
rect 2555 2200 2733 2234
rect 2555 2166 2559 2200
rect 2559 2166 2627 2200
rect 2627 2166 2661 2200
rect 2661 2166 2729 2200
rect 2729 2166 2733 2200
rect 2555 2132 2733 2166
rect 2555 2098 2559 2132
rect 2559 2098 2627 2132
rect 2627 2098 2661 2132
rect 2661 2098 2729 2132
rect 2729 2098 2733 2132
rect 2555 2064 2733 2098
rect 2555 2030 2559 2064
rect 2559 2030 2627 2064
rect 2627 2030 2661 2064
rect 2661 2030 2729 2064
rect 2729 2030 2733 2064
rect 2555 1996 2733 2030
rect 2555 1962 2559 1996
rect 2559 1962 2627 1996
rect 2627 1962 2661 1996
rect 2661 1962 2729 1996
rect 2729 1962 2733 1996
rect 2555 1928 2733 1962
rect 2555 1894 2559 1928
rect 2559 1894 2627 1928
rect 2627 1894 2661 1928
rect 2661 1894 2729 1928
rect 2729 1894 2733 1928
rect 2555 1860 2733 1894
rect 2555 1826 2559 1860
rect 2559 1826 2627 1860
rect 2627 1826 2661 1860
rect 2661 1826 2729 1860
rect 2729 1826 2733 1860
rect 2555 1792 2733 1826
rect 2555 1758 2559 1792
rect 2559 1758 2627 1792
rect 2627 1758 2661 1792
rect 2661 1758 2729 1792
rect 2729 1758 2733 1792
rect 2555 1724 2733 1758
rect 2555 1690 2559 1724
rect 2559 1690 2627 1724
rect 2627 1690 2661 1724
rect 2661 1690 2729 1724
rect 2729 1690 2733 1724
rect 2555 1656 2733 1690
rect 2555 1622 2559 1656
rect 2559 1622 2627 1656
rect 2627 1622 2661 1656
rect 2661 1622 2729 1656
rect 2729 1622 2733 1656
rect 2555 1620 2733 1622
rect 2627 1586 2661 1620
rect 2310 1144 2416 1250
rect 3051 4064 3085 4098
rect 3123 4064 3157 4098
rect 3195 4064 3229 4098
rect 3051 3991 3085 4025
rect 3123 3991 3157 4025
rect 3195 3991 3229 4025
rect 3051 3918 3085 3952
rect 3123 3918 3157 3952
rect 3195 3918 3229 3952
rect 3051 3845 3085 3879
rect 3123 3845 3157 3879
rect 3195 3845 3229 3879
rect 3051 3772 3085 3806
rect 3123 3772 3157 3806
rect 3195 3772 3229 3806
rect 3051 3699 3085 3733
rect 3123 3699 3157 3733
rect 3195 3699 3229 3733
rect 3051 3626 3085 3660
rect 3123 3626 3157 3660
rect 3195 3626 3229 3660
rect 3051 3553 3085 3587
rect 3123 3553 3157 3587
rect 3195 3553 3229 3587
rect 3051 3480 3085 3514
rect 3123 3480 3157 3514
rect 3195 3480 3229 3514
rect 3051 3407 3085 3441
rect 3123 3407 3157 3441
rect 3195 3407 3229 3441
rect 3051 3334 3085 3368
rect 3123 3334 3157 3368
rect 3195 3334 3229 3368
rect 3051 3261 3085 3295
rect 3123 3261 3157 3295
rect 3195 3261 3229 3295
rect 3051 3188 3085 3222
rect 3123 3188 3157 3222
rect 3195 3188 3229 3222
rect 3051 3115 3085 3149
rect 3123 3115 3157 3149
rect 3195 3115 3229 3149
rect 3051 3042 3085 3076
rect 3123 3042 3157 3076
rect 3195 3042 3229 3076
rect 3051 2969 3085 3003
rect 3123 2969 3157 3003
rect 3195 2969 3229 3003
rect 3051 2896 3085 2930
rect 3123 2896 3157 2930
rect 3195 2896 3229 2930
rect 3051 2823 3085 2857
rect 3123 2823 3157 2857
rect 3195 2823 3229 2857
rect 3051 2750 3085 2784
rect 3123 2750 3157 2784
rect 3195 2750 3229 2784
rect 3051 2677 3085 2711
rect 3123 2677 3157 2711
rect 3195 2677 3229 2711
rect 3051 2604 3085 2638
rect 3123 2604 3157 2638
rect 3195 2604 3229 2638
rect 3051 2531 3085 2565
rect 3123 2531 3157 2565
rect 3195 2531 3229 2565
rect 3051 2458 3085 2492
rect 3123 2458 3157 2492
rect 3195 2458 3229 2492
rect 3051 2385 3085 2419
rect 3123 2385 3157 2419
rect 3195 2385 3229 2419
rect 3051 2312 3085 2346
rect 3123 2312 3157 2346
rect 3195 2312 3229 2346
rect 3051 2239 3085 2273
rect 3123 2239 3157 2273
rect 3195 2239 3229 2273
rect 3051 2166 3085 2200
rect 3123 2166 3157 2200
rect 3195 2166 3229 2200
rect 3051 2092 3085 2126
rect 3123 2092 3157 2126
rect 3195 2092 3229 2126
rect 3051 2018 3085 2052
rect 3123 2018 3157 2052
rect 3195 2018 3229 2052
rect 3051 1944 3085 1978
rect 3123 1944 3157 1978
rect 3195 1944 3229 1978
rect 3051 1870 3085 1904
rect 3123 1870 3157 1904
rect 3195 1870 3229 1904
rect 3051 1796 3085 1830
rect 3123 1796 3157 1830
rect 3195 1796 3229 1830
rect 3051 1722 3085 1756
rect 3123 1722 3157 1756
rect 3195 1722 3229 1756
rect 3051 1648 3085 1682
rect 3123 1648 3157 1682
rect 3195 1648 3229 1682
rect 3051 1574 3085 1608
rect 3123 1574 3157 1608
rect 3195 1574 3229 1608
rect 2872 1144 2978 1250
rect 3619 4092 3653 4118
rect 3547 4082 3725 4092
rect 3547 4048 3551 4082
rect 3551 4048 3619 4082
rect 3619 4048 3653 4082
rect 3653 4048 3721 4082
rect 3721 4048 3725 4082
rect 3547 4014 3725 4048
rect 3547 3980 3551 4014
rect 3551 3980 3619 4014
rect 3619 3980 3653 4014
rect 3653 3980 3721 4014
rect 3721 3980 3725 4014
rect 3547 3946 3725 3980
rect 3547 3912 3551 3946
rect 3551 3912 3619 3946
rect 3619 3912 3653 3946
rect 3653 3912 3721 3946
rect 3721 3912 3725 3946
rect 3547 3878 3725 3912
rect 3547 3844 3551 3878
rect 3551 3844 3619 3878
rect 3619 3844 3653 3878
rect 3653 3844 3721 3878
rect 3721 3844 3725 3878
rect 3547 3810 3725 3844
rect 3547 3776 3551 3810
rect 3551 3776 3619 3810
rect 3619 3776 3653 3810
rect 3653 3776 3721 3810
rect 3721 3776 3725 3810
rect 3547 3742 3725 3776
rect 3547 3708 3551 3742
rect 3551 3708 3619 3742
rect 3619 3708 3653 3742
rect 3653 3708 3721 3742
rect 3721 3708 3725 3742
rect 3547 3674 3725 3708
rect 3547 3640 3551 3674
rect 3551 3640 3619 3674
rect 3619 3640 3653 3674
rect 3653 3640 3721 3674
rect 3721 3640 3725 3674
rect 3547 3606 3725 3640
rect 3547 3572 3551 3606
rect 3551 3572 3619 3606
rect 3619 3572 3653 3606
rect 3653 3572 3721 3606
rect 3721 3572 3725 3606
rect 3547 3538 3725 3572
rect 3547 3504 3551 3538
rect 3551 3504 3619 3538
rect 3619 3504 3653 3538
rect 3653 3504 3721 3538
rect 3721 3504 3725 3538
rect 3547 3470 3725 3504
rect 3547 3436 3551 3470
rect 3551 3436 3619 3470
rect 3619 3436 3653 3470
rect 3653 3436 3721 3470
rect 3721 3436 3725 3470
rect 3547 3402 3725 3436
rect 3547 3368 3551 3402
rect 3551 3368 3619 3402
rect 3619 3368 3653 3402
rect 3653 3368 3721 3402
rect 3721 3368 3725 3402
rect 3547 3334 3725 3368
rect 3547 3300 3551 3334
rect 3551 3300 3619 3334
rect 3619 3300 3653 3334
rect 3653 3300 3721 3334
rect 3721 3300 3725 3334
rect 3547 3266 3725 3300
rect 3547 3232 3551 3266
rect 3551 3232 3619 3266
rect 3619 3232 3653 3266
rect 3653 3232 3721 3266
rect 3721 3232 3725 3266
rect 3547 3198 3725 3232
rect 3547 3194 3551 3198
rect 3551 3194 3619 3198
rect 3619 3194 3653 3198
rect 3653 3194 3721 3198
rect 3721 3194 3725 3198
rect 3619 3164 3653 3182
rect 3619 3148 3653 3164
rect 3547 3074 3581 3108
rect 3619 3074 3653 3108
rect 3691 3074 3725 3108
rect 3547 2994 3581 3028
rect 3619 2994 3653 3028
rect 3691 2994 3725 3028
rect 3547 2914 3581 2948
rect 3619 2914 3653 2948
rect 3691 2914 3725 2948
rect 3547 2834 3581 2868
rect 3619 2834 3653 2868
rect 3691 2834 3725 2868
rect 3547 2754 3581 2788
rect 3619 2754 3653 2788
rect 3691 2754 3725 2788
rect 3547 2674 3581 2708
rect 3619 2674 3653 2708
rect 3691 2674 3725 2708
rect 3547 2594 3581 2628
rect 3619 2594 3653 2628
rect 3691 2594 3725 2628
rect 3619 2540 3653 2556
rect 3619 2522 3653 2540
rect 3547 2506 3551 2518
rect 3551 2506 3619 2518
rect 3619 2506 3653 2518
rect 3653 2506 3721 2518
rect 3721 2506 3725 2518
rect 3547 2472 3725 2506
rect 3547 2438 3551 2472
rect 3551 2438 3619 2472
rect 3619 2438 3653 2472
rect 3653 2438 3721 2472
rect 3721 2438 3725 2472
rect 3547 2404 3725 2438
rect 3547 2370 3551 2404
rect 3551 2370 3619 2404
rect 3619 2370 3653 2404
rect 3653 2370 3721 2404
rect 3721 2370 3725 2404
rect 3547 2336 3725 2370
rect 3547 2302 3551 2336
rect 3551 2302 3619 2336
rect 3619 2302 3653 2336
rect 3653 2302 3721 2336
rect 3721 2302 3725 2336
rect 3547 2268 3725 2302
rect 3547 2234 3551 2268
rect 3551 2234 3619 2268
rect 3619 2234 3653 2268
rect 3653 2234 3721 2268
rect 3721 2234 3725 2268
rect 3547 2200 3725 2234
rect 3547 2166 3551 2200
rect 3551 2166 3619 2200
rect 3619 2166 3653 2200
rect 3653 2166 3721 2200
rect 3721 2166 3725 2200
rect 3547 2132 3725 2166
rect 3547 2098 3551 2132
rect 3551 2098 3619 2132
rect 3619 2098 3653 2132
rect 3653 2098 3721 2132
rect 3721 2098 3725 2132
rect 3547 2064 3725 2098
rect 3547 2030 3551 2064
rect 3551 2030 3619 2064
rect 3619 2030 3653 2064
rect 3653 2030 3721 2064
rect 3721 2030 3725 2064
rect 3547 1996 3725 2030
rect 3547 1962 3551 1996
rect 3551 1962 3619 1996
rect 3619 1962 3653 1996
rect 3653 1962 3721 1996
rect 3721 1962 3725 1996
rect 3547 1928 3725 1962
rect 3547 1894 3551 1928
rect 3551 1894 3619 1928
rect 3619 1894 3653 1928
rect 3653 1894 3721 1928
rect 3721 1894 3725 1928
rect 3547 1860 3725 1894
rect 3547 1826 3551 1860
rect 3551 1826 3619 1860
rect 3619 1826 3653 1860
rect 3653 1826 3721 1860
rect 3721 1826 3725 1860
rect 3547 1792 3725 1826
rect 3547 1758 3551 1792
rect 3551 1758 3619 1792
rect 3619 1758 3653 1792
rect 3653 1758 3721 1792
rect 3721 1758 3725 1792
rect 3547 1724 3725 1758
rect 3547 1690 3551 1724
rect 3551 1690 3619 1724
rect 3619 1690 3653 1724
rect 3653 1690 3721 1724
rect 3721 1690 3725 1724
rect 3547 1656 3725 1690
rect 3547 1622 3551 1656
rect 3551 1622 3619 1656
rect 3619 1622 3653 1656
rect 3653 1622 3721 1656
rect 3721 1622 3725 1656
rect 3547 1620 3725 1622
rect 3619 1586 3653 1620
rect 3302 1144 3408 1250
rect 4043 4064 4077 4098
rect 4115 4064 4149 4098
rect 4187 4064 4221 4098
rect 4043 3991 4077 4025
rect 4115 3991 4149 4025
rect 4187 3991 4221 4025
rect 4043 3918 4077 3952
rect 4115 3918 4149 3952
rect 4187 3918 4221 3952
rect 4043 3845 4077 3879
rect 4115 3845 4149 3879
rect 4187 3845 4221 3879
rect 4043 3772 4077 3806
rect 4115 3772 4149 3806
rect 4187 3772 4221 3806
rect 4043 3699 4077 3733
rect 4115 3699 4149 3733
rect 4187 3699 4221 3733
rect 4043 3626 4077 3660
rect 4115 3626 4149 3660
rect 4187 3626 4221 3660
rect 4043 3553 4077 3587
rect 4115 3553 4149 3587
rect 4187 3553 4221 3587
rect 4043 3480 4077 3514
rect 4115 3480 4149 3514
rect 4187 3480 4221 3514
rect 4043 3407 4077 3441
rect 4115 3407 4149 3441
rect 4187 3407 4221 3441
rect 4043 3334 4077 3368
rect 4115 3334 4149 3368
rect 4187 3334 4221 3368
rect 4043 3261 4077 3295
rect 4115 3261 4149 3295
rect 4187 3261 4221 3295
rect 4043 3188 4077 3222
rect 4115 3188 4149 3222
rect 4187 3188 4221 3222
rect 4043 3115 4077 3149
rect 4115 3115 4149 3149
rect 4187 3115 4221 3149
rect 4043 3042 4077 3076
rect 4115 3042 4149 3076
rect 4187 3042 4221 3076
rect 4043 2969 4077 3003
rect 4115 2969 4149 3003
rect 4187 2969 4221 3003
rect 4043 2896 4077 2930
rect 4115 2896 4149 2930
rect 4187 2896 4221 2930
rect 4043 2823 4077 2857
rect 4115 2823 4149 2857
rect 4187 2823 4221 2857
rect 4043 2750 4077 2784
rect 4115 2750 4149 2784
rect 4187 2750 4221 2784
rect 4043 2677 4077 2711
rect 4115 2677 4149 2711
rect 4187 2677 4221 2711
rect 4043 2604 4077 2638
rect 4115 2604 4149 2638
rect 4187 2604 4221 2638
rect 4043 2531 4077 2565
rect 4115 2531 4149 2565
rect 4187 2531 4221 2565
rect 4043 2458 4077 2492
rect 4115 2458 4149 2492
rect 4187 2458 4221 2492
rect 4043 2385 4077 2419
rect 4115 2385 4149 2419
rect 4187 2385 4221 2419
rect 4043 2312 4077 2346
rect 4115 2312 4149 2346
rect 4187 2312 4221 2346
rect 4043 2239 4077 2273
rect 4115 2239 4149 2273
rect 4187 2239 4221 2273
rect 4043 2166 4077 2200
rect 4115 2166 4149 2200
rect 4187 2166 4221 2200
rect 4043 2092 4077 2126
rect 4115 2092 4149 2126
rect 4187 2092 4221 2126
rect 4043 2018 4077 2052
rect 4115 2018 4149 2052
rect 4187 2018 4221 2052
rect 4043 1944 4077 1978
rect 4115 1944 4149 1978
rect 4187 1944 4221 1978
rect 4043 1870 4077 1904
rect 4115 1870 4149 1904
rect 4187 1870 4221 1904
rect 4043 1796 4077 1830
rect 4115 1796 4149 1830
rect 4187 1796 4221 1830
rect 4043 1722 4077 1756
rect 4115 1722 4149 1756
rect 4187 1722 4221 1756
rect 4043 1648 4077 1682
rect 4115 1648 4149 1682
rect 4187 1648 4221 1682
rect 4043 1574 4077 1608
rect 4115 1574 4149 1608
rect 4187 1574 4221 1608
rect 3864 1144 3970 1250
rect 4611 4092 4645 4118
rect 4539 4082 4717 4092
rect 4539 4048 4543 4082
rect 4543 4048 4611 4082
rect 4611 4048 4645 4082
rect 4645 4048 4713 4082
rect 4713 4048 4717 4082
rect 4539 4014 4717 4048
rect 4539 3980 4543 4014
rect 4543 3980 4611 4014
rect 4611 3980 4645 4014
rect 4645 3980 4713 4014
rect 4713 3980 4717 4014
rect 4539 3946 4717 3980
rect 4539 3912 4543 3946
rect 4543 3912 4611 3946
rect 4611 3912 4645 3946
rect 4645 3912 4713 3946
rect 4713 3912 4717 3946
rect 4539 3878 4717 3912
rect 4539 3844 4543 3878
rect 4543 3844 4611 3878
rect 4611 3844 4645 3878
rect 4645 3844 4713 3878
rect 4713 3844 4717 3878
rect 4539 3810 4717 3844
rect 4539 3776 4543 3810
rect 4543 3776 4611 3810
rect 4611 3776 4645 3810
rect 4645 3776 4713 3810
rect 4713 3776 4717 3810
rect 4539 3742 4717 3776
rect 4539 3708 4543 3742
rect 4543 3708 4611 3742
rect 4611 3708 4645 3742
rect 4645 3708 4713 3742
rect 4713 3708 4717 3742
rect 4539 3674 4717 3708
rect 4539 3640 4543 3674
rect 4543 3640 4611 3674
rect 4611 3640 4645 3674
rect 4645 3640 4713 3674
rect 4713 3640 4717 3674
rect 4539 3606 4717 3640
rect 4539 3572 4543 3606
rect 4543 3572 4611 3606
rect 4611 3572 4645 3606
rect 4645 3572 4713 3606
rect 4713 3572 4717 3606
rect 4539 3538 4717 3572
rect 4539 3504 4543 3538
rect 4543 3504 4611 3538
rect 4611 3504 4645 3538
rect 4645 3504 4713 3538
rect 4713 3504 4717 3538
rect 4539 3470 4717 3504
rect 4539 3436 4543 3470
rect 4543 3436 4611 3470
rect 4611 3436 4645 3470
rect 4645 3436 4713 3470
rect 4713 3436 4717 3470
rect 4539 3402 4717 3436
rect 4539 3368 4543 3402
rect 4543 3368 4611 3402
rect 4611 3368 4645 3402
rect 4645 3368 4713 3402
rect 4713 3368 4717 3402
rect 4539 3334 4717 3368
rect 4539 3300 4543 3334
rect 4543 3300 4611 3334
rect 4611 3300 4645 3334
rect 4645 3300 4713 3334
rect 4713 3300 4717 3334
rect 4539 3266 4717 3300
rect 4539 3232 4543 3266
rect 4543 3232 4611 3266
rect 4611 3232 4645 3266
rect 4645 3232 4713 3266
rect 4713 3232 4717 3266
rect 4539 3198 4717 3232
rect 4539 3194 4543 3198
rect 4543 3194 4611 3198
rect 4611 3194 4645 3198
rect 4645 3194 4713 3198
rect 4713 3194 4717 3198
rect 4611 3164 4645 3182
rect 4611 3148 4645 3164
rect 4539 3074 4573 3108
rect 4611 3074 4645 3108
rect 4683 3074 4717 3108
rect 4539 2994 4573 3028
rect 4611 2994 4645 3028
rect 4683 2994 4717 3028
rect 4539 2914 4573 2948
rect 4611 2914 4645 2948
rect 4683 2914 4717 2948
rect 4539 2834 4573 2868
rect 4611 2834 4645 2868
rect 4683 2834 4717 2868
rect 4539 2754 4573 2788
rect 4611 2754 4645 2788
rect 4683 2754 4717 2788
rect 4539 2674 4573 2708
rect 4611 2674 4645 2708
rect 4683 2674 4717 2708
rect 4539 2594 4573 2628
rect 4611 2594 4645 2628
rect 4683 2594 4717 2628
rect 4611 2540 4645 2556
rect 4611 2522 4645 2540
rect 4539 2506 4543 2518
rect 4543 2506 4611 2518
rect 4611 2506 4645 2518
rect 4645 2506 4713 2518
rect 4713 2506 4717 2518
rect 4539 2472 4717 2506
rect 4539 2438 4543 2472
rect 4543 2438 4611 2472
rect 4611 2438 4645 2472
rect 4645 2438 4713 2472
rect 4713 2438 4717 2472
rect 4539 2404 4717 2438
rect 4539 2370 4543 2404
rect 4543 2370 4611 2404
rect 4611 2370 4645 2404
rect 4645 2370 4713 2404
rect 4713 2370 4717 2404
rect 4539 2336 4717 2370
rect 4539 2302 4543 2336
rect 4543 2302 4611 2336
rect 4611 2302 4645 2336
rect 4645 2302 4713 2336
rect 4713 2302 4717 2336
rect 4539 2268 4717 2302
rect 4539 2234 4543 2268
rect 4543 2234 4611 2268
rect 4611 2234 4645 2268
rect 4645 2234 4713 2268
rect 4713 2234 4717 2268
rect 4539 2200 4717 2234
rect 4539 2166 4543 2200
rect 4543 2166 4611 2200
rect 4611 2166 4645 2200
rect 4645 2166 4713 2200
rect 4713 2166 4717 2200
rect 4539 2132 4717 2166
rect 4539 2098 4543 2132
rect 4543 2098 4611 2132
rect 4611 2098 4645 2132
rect 4645 2098 4713 2132
rect 4713 2098 4717 2132
rect 4539 2064 4717 2098
rect 4539 2030 4543 2064
rect 4543 2030 4611 2064
rect 4611 2030 4645 2064
rect 4645 2030 4713 2064
rect 4713 2030 4717 2064
rect 4539 1996 4717 2030
rect 4539 1962 4543 1996
rect 4543 1962 4611 1996
rect 4611 1962 4645 1996
rect 4645 1962 4713 1996
rect 4713 1962 4717 1996
rect 4539 1928 4717 1962
rect 4539 1894 4543 1928
rect 4543 1894 4611 1928
rect 4611 1894 4645 1928
rect 4645 1894 4713 1928
rect 4713 1894 4717 1928
rect 4539 1860 4717 1894
rect 4539 1826 4543 1860
rect 4543 1826 4611 1860
rect 4611 1826 4645 1860
rect 4645 1826 4713 1860
rect 4713 1826 4717 1860
rect 4539 1792 4717 1826
rect 4539 1758 4543 1792
rect 4543 1758 4611 1792
rect 4611 1758 4645 1792
rect 4645 1758 4713 1792
rect 4713 1758 4717 1792
rect 4539 1724 4717 1758
rect 4539 1690 4543 1724
rect 4543 1690 4611 1724
rect 4611 1690 4645 1724
rect 4645 1690 4713 1724
rect 4713 1690 4717 1724
rect 4539 1656 4717 1690
rect 4539 1622 4543 1656
rect 4543 1622 4611 1656
rect 4611 1622 4645 1656
rect 4645 1622 4713 1656
rect 4713 1622 4717 1656
rect 4539 1620 4717 1622
rect 4611 1586 4645 1620
rect 4294 1144 4400 1250
rect 5035 4064 5069 4098
rect 5107 4064 5141 4098
rect 5179 4064 5213 4098
rect 5035 3991 5069 4025
rect 5107 3991 5141 4025
rect 5179 3991 5213 4025
rect 5035 3918 5069 3952
rect 5107 3918 5141 3952
rect 5179 3918 5213 3952
rect 5035 3845 5069 3879
rect 5107 3845 5141 3879
rect 5179 3845 5213 3879
rect 5035 3772 5069 3806
rect 5107 3772 5141 3806
rect 5179 3772 5213 3806
rect 5035 3699 5069 3733
rect 5107 3699 5141 3733
rect 5179 3699 5213 3733
rect 5035 3626 5069 3660
rect 5107 3626 5141 3660
rect 5179 3626 5213 3660
rect 5035 3553 5069 3587
rect 5107 3553 5141 3587
rect 5179 3553 5213 3587
rect 5035 3480 5069 3514
rect 5107 3480 5141 3514
rect 5179 3480 5213 3514
rect 5035 3407 5069 3441
rect 5107 3407 5141 3441
rect 5179 3407 5213 3441
rect 5035 3334 5069 3368
rect 5107 3334 5141 3368
rect 5179 3334 5213 3368
rect 5035 3261 5069 3295
rect 5107 3261 5141 3295
rect 5179 3261 5213 3295
rect 5035 3188 5069 3222
rect 5107 3188 5141 3222
rect 5179 3188 5213 3222
rect 5035 3115 5069 3149
rect 5107 3115 5141 3149
rect 5179 3115 5213 3149
rect 5035 3042 5069 3076
rect 5107 3042 5141 3076
rect 5179 3042 5213 3076
rect 5035 2969 5069 3003
rect 5107 2969 5141 3003
rect 5179 2969 5213 3003
rect 5035 2896 5069 2930
rect 5107 2896 5141 2930
rect 5179 2896 5213 2930
rect 5035 2823 5069 2857
rect 5107 2823 5141 2857
rect 5179 2823 5213 2857
rect 5035 2750 5069 2784
rect 5107 2750 5141 2784
rect 5179 2750 5213 2784
rect 5035 2677 5069 2711
rect 5107 2677 5141 2711
rect 5179 2677 5213 2711
rect 5035 2604 5069 2638
rect 5107 2604 5141 2638
rect 5179 2604 5213 2638
rect 5035 2531 5069 2565
rect 5107 2531 5141 2565
rect 5179 2531 5213 2565
rect 5035 2458 5069 2492
rect 5107 2458 5141 2492
rect 5179 2458 5213 2492
rect 5035 2385 5069 2419
rect 5107 2385 5141 2419
rect 5179 2385 5213 2419
rect 5035 2312 5069 2346
rect 5107 2312 5141 2346
rect 5179 2312 5213 2346
rect 5035 2239 5069 2273
rect 5107 2239 5141 2273
rect 5179 2239 5213 2273
rect 5035 2166 5069 2200
rect 5107 2166 5141 2200
rect 5179 2166 5213 2200
rect 5035 2092 5069 2126
rect 5107 2092 5141 2126
rect 5179 2092 5213 2126
rect 5035 2018 5069 2052
rect 5107 2018 5141 2052
rect 5179 2018 5213 2052
rect 5035 1944 5069 1978
rect 5107 1944 5141 1978
rect 5179 1944 5213 1978
rect 5035 1870 5069 1904
rect 5107 1870 5141 1904
rect 5179 1870 5213 1904
rect 5035 1796 5069 1830
rect 5107 1796 5141 1830
rect 5179 1796 5213 1830
rect 5035 1722 5069 1756
rect 5107 1722 5141 1756
rect 5179 1722 5213 1756
rect 5035 1648 5069 1682
rect 5107 1648 5141 1682
rect 5179 1648 5213 1682
rect 5035 1574 5069 1608
rect 5107 1574 5141 1608
rect 5179 1574 5213 1608
rect 4856 1144 4962 1250
rect 5603 4092 5637 4118
rect 5531 4082 5709 4092
rect 5531 4048 5535 4082
rect 5535 4048 5603 4082
rect 5603 4048 5637 4082
rect 5637 4048 5705 4082
rect 5705 4048 5709 4082
rect 5531 4014 5709 4048
rect 5531 3980 5535 4014
rect 5535 3980 5603 4014
rect 5603 3980 5637 4014
rect 5637 3980 5705 4014
rect 5705 3980 5709 4014
rect 5531 3946 5709 3980
rect 5531 3912 5535 3946
rect 5535 3912 5603 3946
rect 5603 3912 5637 3946
rect 5637 3912 5705 3946
rect 5705 3912 5709 3946
rect 5531 3878 5709 3912
rect 5531 3844 5535 3878
rect 5535 3844 5603 3878
rect 5603 3844 5637 3878
rect 5637 3844 5705 3878
rect 5705 3844 5709 3878
rect 5531 3810 5709 3844
rect 5531 3776 5535 3810
rect 5535 3776 5603 3810
rect 5603 3776 5637 3810
rect 5637 3776 5705 3810
rect 5705 3776 5709 3810
rect 5531 3742 5709 3776
rect 5531 3708 5535 3742
rect 5535 3708 5603 3742
rect 5603 3708 5637 3742
rect 5637 3708 5705 3742
rect 5705 3708 5709 3742
rect 5531 3674 5709 3708
rect 5531 3640 5535 3674
rect 5535 3640 5603 3674
rect 5603 3640 5637 3674
rect 5637 3640 5705 3674
rect 5705 3640 5709 3674
rect 5531 3606 5709 3640
rect 5531 3572 5535 3606
rect 5535 3572 5603 3606
rect 5603 3572 5637 3606
rect 5637 3572 5705 3606
rect 5705 3572 5709 3606
rect 5531 3538 5709 3572
rect 5531 3504 5535 3538
rect 5535 3504 5603 3538
rect 5603 3504 5637 3538
rect 5637 3504 5705 3538
rect 5705 3504 5709 3538
rect 5531 3470 5709 3504
rect 5531 3436 5535 3470
rect 5535 3436 5603 3470
rect 5603 3436 5637 3470
rect 5637 3436 5705 3470
rect 5705 3436 5709 3470
rect 5531 3402 5709 3436
rect 5531 3368 5535 3402
rect 5535 3368 5603 3402
rect 5603 3368 5637 3402
rect 5637 3368 5705 3402
rect 5705 3368 5709 3402
rect 5531 3334 5709 3368
rect 5531 3300 5535 3334
rect 5535 3300 5603 3334
rect 5603 3300 5637 3334
rect 5637 3300 5705 3334
rect 5705 3300 5709 3334
rect 5531 3266 5709 3300
rect 5531 3232 5535 3266
rect 5535 3232 5603 3266
rect 5603 3232 5637 3266
rect 5637 3232 5705 3266
rect 5705 3232 5709 3266
rect 5531 3198 5709 3232
rect 5531 3194 5535 3198
rect 5535 3194 5603 3198
rect 5603 3194 5637 3198
rect 5637 3194 5705 3198
rect 5705 3194 5709 3198
rect 5603 3164 5637 3182
rect 5603 3148 5637 3164
rect 5531 3074 5565 3108
rect 5603 3074 5637 3108
rect 5675 3074 5709 3108
rect 5531 2994 5565 3028
rect 5603 2994 5637 3028
rect 5675 2994 5709 3028
rect 5531 2914 5565 2948
rect 5603 2914 5637 2948
rect 5675 2914 5709 2948
rect 5531 2834 5565 2868
rect 5603 2834 5637 2868
rect 5675 2834 5709 2868
rect 5531 2754 5565 2788
rect 5603 2754 5637 2788
rect 5675 2754 5709 2788
rect 5531 2674 5565 2708
rect 5603 2674 5637 2708
rect 5675 2674 5709 2708
rect 5531 2594 5565 2628
rect 5603 2594 5637 2628
rect 5675 2594 5709 2628
rect 5603 2540 5637 2556
rect 5603 2522 5637 2540
rect 5531 2506 5535 2518
rect 5535 2506 5603 2518
rect 5603 2506 5637 2518
rect 5637 2506 5705 2518
rect 5705 2506 5709 2518
rect 5531 2472 5709 2506
rect 5531 2438 5535 2472
rect 5535 2438 5603 2472
rect 5603 2438 5637 2472
rect 5637 2438 5705 2472
rect 5705 2438 5709 2472
rect 5531 2404 5709 2438
rect 5531 2370 5535 2404
rect 5535 2370 5603 2404
rect 5603 2370 5637 2404
rect 5637 2370 5705 2404
rect 5705 2370 5709 2404
rect 5531 2336 5709 2370
rect 5531 2302 5535 2336
rect 5535 2302 5603 2336
rect 5603 2302 5637 2336
rect 5637 2302 5705 2336
rect 5705 2302 5709 2336
rect 5531 2268 5709 2302
rect 5531 2234 5535 2268
rect 5535 2234 5603 2268
rect 5603 2234 5637 2268
rect 5637 2234 5705 2268
rect 5705 2234 5709 2268
rect 5531 2200 5709 2234
rect 5531 2166 5535 2200
rect 5535 2166 5603 2200
rect 5603 2166 5637 2200
rect 5637 2166 5705 2200
rect 5705 2166 5709 2200
rect 5531 2132 5709 2166
rect 5531 2098 5535 2132
rect 5535 2098 5603 2132
rect 5603 2098 5637 2132
rect 5637 2098 5705 2132
rect 5705 2098 5709 2132
rect 5531 2064 5709 2098
rect 5531 2030 5535 2064
rect 5535 2030 5603 2064
rect 5603 2030 5637 2064
rect 5637 2030 5705 2064
rect 5705 2030 5709 2064
rect 5531 1996 5709 2030
rect 5531 1962 5535 1996
rect 5535 1962 5603 1996
rect 5603 1962 5637 1996
rect 5637 1962 5705 1996
rect 5705 1962 5709 1996
rect 5531 1928 5709 1962
rect 5531 1894 5535 1928
rect 5535 1894 5603 1928
rect 5603 1894 5637 1928
rect 5637 1894 5705 1928
rect 5705 1894 5709 1928
rect 5531 1860 5709 1894
rect 5531 1826 5535 1860
rect 5535 1826 5603 1860
rect 5603 1826 5637 1860
rect 5637 1826 5705 1860
rect 5705 1826 5709 1860
rect 5531 1792 5709 1826
rect 5531 1758 5535 1792
rect 5535 1758 5603 1792
rect 5603 1758 5637 1792
rect 5637 1758 5705 1792
rect 5705 1758 5709 1792
rect 5531 1724 5709 1758
rect 5531 1690 5535 1724
rect 5535 1690 5603 1724
rect 5603 1690 5637 1724
rect 5637 1690 5705 1724
rect 5705 1690 5709 1724
rect 5531 1656 5709 1690
rect 5531 1622 5535 1656
rect 5535 1622 5603 1656
rect 5603 1622 5637 1656
rect 5637 1622 5705 1656
rect 5705 1622 5709 1656
rect 5531 1620 5709 1622
rect 5603 1586 5637 1620
rect 5286 1144 5392 1250
rect 6027 4064 6061 4098
rect 6099 4064 6133 4098
rect 6171 4064 6205 4098
rect 6027 3991 6061 4025
rect 6099 3991 6133 4025
rect 6171 3991 6205 4025
rect 6027 3918 6061 3952
rect 6099 3918 6133 3952
rect 6171 3918 6205 3952
rect 6027 3845 6061 3879
rect 6099 3845 6133 3879
rect 6171 3845 6205 3879
rect 6027 3772 6061 3806
rect 6099 3772 6133 3806
rect 6171 3772 6205 3806
rect 6027 3699 6061 3733
rect 6099 3699 6133 3733
rect 6171 3699 6205 3733
rect 6027 3626 6061 3660
rect 6099 3626 6133 3660
rect 6171 3626 6205 3660
rect 6027 3553 6061 3587
rect 6099 3553 6133 3587
rect 6171 3553 6205 3587
rect 6027 3480 6061 3514
rect 6099 3480 6133 3514
rect 6171 3480 6205 3514
rect 6027 3407 6061 3441
rect 6099 3407 6133 3441
rect 6171 3407 6205 3441
rect 6027 3334 6061 3368
rect 6099 3334 6133 3368
rect 6171 3334 6205 3368
rect 6027 3261 6061 3295
rect 6099 3261 6133 3295
rect 6171 3261 6205 3295
rect 6027 3188 6061 3222
rect 6099 3188 6133 3222
rect 6171 3188 6205 3222
rect 6027 3115 6061 3149
rect 6099 3115 6133 3149
rect 6171 3115 6205 3149
rect 6027 3042 6061 3076
rect 6099 3042 6133 3076
rect 6171 3042 6205 3076
rect 6027 2969 6061 3003
rect 6099 2969 6133 3003
rect 6171 2969 6205 3003
rect 6027 2896 6061 2930
rect 6099 2896 6133 2930
rect 6171 2896 6205 2930
rect 6027 2823 6061 2857
rect 6099 2823 6133 2857
rect 6171 2823 6205 2857
rect 6027 2750 6061 2784
rect 6099 2750 6133 2784
rect 6171 2750 6205 2784
rect 6027 2677 6061 2711
rect 6099 2677 6133 2711
rect 6171 2677 6205 2711
rect 6027 2604 6061 2638
rect 6099 2604 6133 2638
rect 6171 2604 6205 2638
rect 6027 2531 6061 2565
rect 6099 2531 6133 2565
rect 6171 2531 6205 2565
rect 6027 2458 6061 2492
rect 6099 2458 6133 2492
rect 6171 2458 6205 2492
rect 6027 2385 6061 2419
rect 6099 2385 6133 2419
rect 6171 2385 6205 2419
rect 6027 2312 6061 2346
rect 6099 2312 6133 2346
rect 6171 2312 6205 2346
rect 6027 2239 6061 2273
rect 6099 2239 6133 2273
rect 6171 2239 6205 2273
rect 6027 2166 6061 2200
rect 6099 2166 6133 2200
rect 6171 2166 6205 2200
rect 6027 2092 6061 2126
rect 6099 2092 6133 2126
rect 6171 2092 6205 2126
rect 6027 2018 6061 2052
rect 6099 2018 6133 2052
rect 6171 2018 6205 2052
rect 6027 1944 6061 1978
rect 6099 1944 6133 1978
rect 6171 1944 6205 1978
rect 6027 1870 6061 1904
rect 6099 1870 6133 1904
rect 6171 1870 6205 1904
rect 6027 1796 6061 1830
rect 6099 1796 6133 1830
rect 6171 1796 6205 1830
rect 6027 1722 6061 1756
rect 6099 1722 6133 1756
rect 6171 1722 6205 1756
rect 6027 1648 6061 1682
rect 6099 1648 6133 1682
rect 6171 1648 6205 1682
rect 6027 1574 6061 1608
rect 6099 1574 6133 1608
rect 6171 1574 6205 1608
rect 5848 1144 5954 1250
rect 6595 4092 6629 4118
rect 6523 4082 6701 4092
rect 6523 4048 6527 4082
rect 6527 4048 6595 4082
rect 6595 4048 6629 4082
rect 6629 4048 6697 4082
rect 6697 4048 6701 4082
rect 6523 4014 6701 4048
rect 6523 3980 6527 4014
rect 6527 3980 6595 4014
rect 6595 3980 6629 4014
rect 6629 3980 6697 4014
rect 6697 3980 6701 4014
rect 6523 3946 6701 3980
rect 6523 3912 6527 3946
rect 6527 3912 6595 3946
rect 6595 3912 6629 3946
rect 6629 3912 6697 3946
rect 6697 3912 6701 3946
rect 6523 3878 6701 3912
rect 6523 3844 6527 3878
rect 6527 3844 6595 3878
rect 6595 3844 6629 3878
rect 6629 3844 6697 3878
rect 6697 3844 6701 3878
rect 6523 3810 6701 3844
rect 6523 3776 6527 3810
rect 6527 3776 6595 3810
rect 6595 3776 6629 3810
rect 6629 3776 6697 3810
rect 6697 3776 6701 3810
rect 6523 3742 6701 3776
rect 6523 3708 6527 3742
rect 6527 3708 6595 3742
rect 6595 3708 6629 3742
rect 6629 3708 6697 3742
rect 6697 3708 6701 3742
rect 6523 3674 6701 3708
rect 6523 3640 6527 3674
rect 6527 3640 6595 3674
rect 6595 3640 6629 3674
rect 6629 3640 6697 3674
rect 6697 3640 6701 3674
rect 6523 3606 6701 3640
rect 6523 3572 6527 3606
rect 6527 3572 6595 3606
rect 6595 3572 6629 3606
rect 6629 3572 6697 3606
rect 6697 3572 6701 3606
rect 6523 3538 6701 3572
rect 6523 3504 6527 3538
rect 6527 3504 6595 3538
rect 6595 3504 6629 3538
rect 6629 3504 6697 3538
rect 6697 3504 6701 3538
rect 6523 3470 6701 3504
rect 6523 3436 6527 3470
rect 6527 3436 6595 3470
rect 6595 3436 6629 3470
rect 6629 3436 6697 3470
rect 6697 3436 6701 3470
rect 6523 3402 6701 3436
rect 6523 3368 6527 3402
rect 6527 3368 6595 3402
rect 6595 3368 6629 3402
rect 6629 3368 6697 3402
rect 6697 3368 6701 3402
rect 6523 3334 6701 3368
rect 6523 3300 6527 3334
rect 6527 3300 6595 3334
rect 6595 3300 6629 3334
rect 6629 3300 6697 3334
rect 6697 3300 6701 3334
rect 6523 3266 6701 3300
rect 6523 3232 6527 3266
rect 6527 3232 6595 3266
rect 6595 3232 6629 3266
rect 6629 3232 6697 3266
rect 6697 3232 6701 3266
rect 6523 3198 6701 3232
rect 6523 3194 6527 3198
rect 6527 3194 6595 3198
rect 6595 3194 6629 3198
rect 6629 3194 6697 3198
rect 6697 3194 6701 3198
rect 6595 3164 6629 3182
rect 6595 3148 6629 3164
rect 6523 3074 6557 3108
rect 6595 3074 6629 3108
rect 6667 3074 6701 3108
rect 6523 2994 6557 3028
rect 6595 2994 6629 3028
rect 6667 2994 6701 3028
rect 6523 2914 6557 2948
rect 6595 2914 6629 2948
rect 6667 2914 6701 2948
rect 6523 2834 6557 2868
rect 6595 2834 6629 2868
rect 6667 2834 6701 2868
rect 6523 2754 6557 2788
rect 6595 2754 6629 2788
rect 6667 2754 6701 2788
rect 6523 2674 6557 2708
rect 6595 2674 6629 2708
rect 6667 2674 6701 2708
rect 6523 2594 6557 2628
rect 6595 2594 6629 2628
rect 6667 2594 6701 2628
rect 6595 2540 6629 2556
rect 6595 2522 6629 2540
rect 6523 2506 6527 2518
rect 6527 2506 6595 2518
rect 6595 2506 6629 2518
rect 6629 2506 6697 2518
rect 6697 2506 6701 2518
rect 6523 2472 6701 2506
rect 6523 2438 6527 2472
rect 6527 2438 6595 2472
rect 6595 2438 6629 2472
rect 6629 2438 6697 2472
rect 6697 2438 6701 2472
rect 6523 2404 6701 2438
rect 6523 2370 6527 2404
rect 6527 2370 6595 2404
rect 6595 2370 6629 2404
rect 6629 2370 6697 2404
rect 6697 2370 6701 2404
rect 6523 2336 6701 2370
rect 6523 2302 6527 2336
rect 6527 2302 6595 2336
rect 6595 2302 6629 2336
rect 6629 2302 6697 2336
rect 6697 2302 6701 2336
rect 6523 2268 6701 2302
rect 6523 2234 6527 2268
rect 6527 2234 6595 2268
rect 6595 2234 6629 2268
rect 6629 2234 6697 2268
rect 6697 2234 6701 2268
rect 6523 2200 6701 2234
rect 6523 2166 6527 2200
rect 6527 2166 6595 2200
rect 6595 2166 6629 2200
rect 6629 2166 6697 2200
rect 6697 2166 6701 2200
rect 6523 2132 6701 2166
rect 6523 2098 6527 2132
rect 6527 2098 6595 2132
rect 6595 2098 6629 2132
rect 6629 2098 6697 2132
rect 6697 2098 6701 2132
rect 6523 2064 6701 2098
rect 6523 2030 6527 2064
rect 6527 2030 6595 2064
rect 6595 2030 6629 2064
rect 6629 2030 6697 2064
rect 6697 2030 6701 2064
rect 6523 1996 6701 2030
rect 6523 1962 6527 1996
rect 6527 1962 6595 1996
rect 6595 1962 6629 1996
rect 6629 1962 6697 1996
rect 6697 1962 6701 1996
rect 6523 1928 6701 1962
rect 6523 1894 6527 1928
rect 6527 1894 6595 1928
rect 6595 1894 6629 1928
rect 6629 1894 6697 1928
rect 6697 1894 6701 1928
rect 6523 1860 6701 1894
rect 6523 1826 6527 1860
rect 6527 1826 6595 1860
rect 6595 1826 6629 1860
rect 6629 1826 6697 1860
rect 6697 1826 6701 1860
rect 6523 1792 6701 1826
rect 6523 1758 6527 1792
rect 6527 1758 6595 1792
rect 6595 1758 6629 1792
rect 6629 1758 6697 1792
rect 6697 1758 6701 1792
rect 6523 1724 6701 1758
rect 6523 1690 6527 1724
rect 6527 1690 6595 1724
rect 6595 1690 6629 1724
rect 6629 1690 6697 1724
rect 6697 1690 6701 1724
rect 6523 1656 6701 1690
rect 6523 1622 6527 1656
rect 6527 1622 6595 1656
rect 6595 1622 6629 1656
rect 6629 1622 6697 1656
rect 6697 1622 6701 1656
rect 6523 1620 6701 1622
rect 6595 1586 6629 1620
rect 6278 1144 6384 1250
rect 7019 4064 7053 4098
rect 7091 4064 7125 4098
rect 7163 4064 7197 4098
rect 7019 3991 7053 4025
rect 7091 3991 7125 4025
rect 7163 3991 7197 4025
rect 7019 3918 7053 3952
rect 7091 3918 7125 3952
rect 7163 3918 7197 3952
rect 7019 3845 7053 3879
rect 7091 3845 7125 3879
rect 7163 3845 7197 3879
rect 7019 3772 7053 3806
rect 7091 3772 7125 3806
rect 7163 3772 7197 3806
rect 7019 3699 7053 3733
rect 7091 3699 7125 3733
rect 7163 3699 7197 3733
rect 7019 3626 7053 3660
rect 7091 3626 7125 3660
rect 7163 3626 7197 3660
rect 7019 3553 7053 3587
rect 7091 3553 7125 3587
rect 7163 3553 7197 3587
rect 7019 3480 7053 3514
rect 7091 3480 7125 3514
rect 7163 3480 7197 3514
rect 7019 3407 7053 3441
rect 7091 3407 7125 3441
rect 7163 3407 7197 3441
rect 7019 3334 7053 3368
rect 7091 3334 7125 3368
rect 7163 3334 7197 3368
rect 7019 3261 7053 3295
rect 7091 3261 7125 3295
rect 7163 3261 7197 3295
rect 7019 3188 7053 3222
rect 7091 3188 7125 3222
rect 7163 3188 7197 3222
rect 7019 3115 7053 3149
rect 7091 3115 7125 3149
rect 7163 3115 7197 3149
rect 7019 3042 7053 3076
rect 7091 3042 7125 3076
rect 7163 3042 7197 3076
rect 7019 2969 7053 3003
rect 7091 2969 7125 3003
rect 7163 2969 7197 3003
rect 7019 2896 7053 2930
rect 7091 2896 7125 2930
rect 7163 2896 7197 2930
rect 7019 2823 7053 2857
rect 7091 2823 7125 2857
rect 7163 2823 7197 2857
rect 7019 2750 7053 2784
rect 7091 2750 7125 2784
rect 7163 2750 7197 2784
rect 7019 2677 7053 2711
rect 7091 2677 7125 2711
rect 7163 2677 7197 2711
rect 7019 2604 7053 2638
rect 7091 2604 7125 2638
rect 7163 2604 7197 2638
rect 7019 2531 7053 2565
rect 7091 2531 7125 2565
rect 7163 2531 7197 2565
rect 7019 2458 7053 2492
rect 7091 2458 7125 2492
rect 7163 2458 7197 2492
rect 7019 2385 7053 2419
rect 7091 2385 7125 2419
rect 7163 2385 7197 2419
rect 7019 2312 7053 2346
rect 7091 2312 7125 2346
rect 7163 2312 7197 2346
rect 7019 2239 7053 2273
rect 7091 2239 7125 2273
rect 7163 2239 7197 2273
rect 7019 2166 7053 2200
rect 7091 2166 7125 2200
rect 7163 2166 7197 2200
rect 7019 2092 7053 2126
rect 7091 2092 7125 2126
rect 7163 2092 7197 2126
rect 7019 2018 7053 2052
rect 7091 2018 7125 2052
rect 7163 2018 7197 2052
rect 7019 1944 7053 1978
rect 7091 1944 7125 1978
rect 7163 1944 7197 1978
rect 7019 1870 7053 1904
rect 7091 1870 7125 1904
rect 7163 1870 7197 1904
rect 7019 1796 7053 1830
rect 7091 1796 7125 1830
rect 7163 1796 7197 1830
rect 7019 1722 7053 1756
rect 7091 1722 7125 1756
rect 7163 1722 7197 1756
rect 7019 1648 7053 1682
rect 7091 1648 7125 1682
rect 7163 1648 7197 1682
rect 7019 1574 7053 1608
rect 7091 1574 7125 1608
rect 7163 1574 7197 1608
rect 6840 1144 6946 1250
rect 7587 4092 7621 4118
rect 7515 4082 7693 4092
rect 7515 4048 7519 4082
rect 7519 4048 7587 4082
rect 7587 4048 7621 4082
rect 7621 4048 7689 4082
rect 7689 4048 7693 4082
rect 7515 4014 7693 4048
rect 7515 3980 7519 4014
rect 7519 3980 7587 4014
rect 7587 3980 7621 4014
rect 7621 3980 7689 4014
rect 7689 3980 7693 4014
rect 7515 3946 7693 3980
rect 7515 3912 7519 3946
rect 7519 3912 7587 3946
rect 7587 3912 7621 3946
rect 7621 3912 7689 3946
rect 7689 3912 7693 3946
rect 7515 3878 7693 3912
rect 7515 3844 7519 3878
rect 7519 3844 7587 3878
rect 7587 3844 7621 3878
rect 7621 3844 7689 3878
rect 7689 3844 7693 3878
rect 7515 3810 7693 3844
rect 7515 3776 7519 3810
rect 7519 3776 7587 3810
rect 7587 3776 7621 3810
rect 7621 3776 7689 3810
rect 7689 3776 7693 3810
rect 7515 3742 7693 3776
rect 7515 3708 7519 3742
rect 7519 3708 7587 3742
rect 7587 3708 7621 3742
rect 7621 3708 7689 3742
rect 7689 3708 7693 3742
rect 7515 3674 7693 3708
rect 7515 3640 7519 3674
rect 7519 3640 7587 3674
rect 7587 3640 7621 3674
rect 7621 3640 7689 3674
rect 7689 3640 7693 3674
rect 7515 3606 7693 3640
rect 7515 3572 7519 3606
rect 7519 3572 7587 3606
rect 7587 3572 7621 3606
rect 7621 3572 7689 3606
rect 7689 3572 7693 3606
rect 7515 3538 7693 3572
rect 7515 3504 7519 3538
rect 7519 3504 7587 3538
rect 7587 3504 7621 3538
rect 7621 3504 7689 3538
rect 7689 3504 7693 3538
rect 7515 3470 7693 3504
rect 7515 3436 7519 3470
rect 7519 3436 7587 3470
rect 7587 3436 7621 3470
rect 7621 3436 7689 3470
rect 7689 3436 7693 3470
rect 7515 3402 7693 3436
rect 7515 3368 7519 3402
rect 7519 3368 7587 3402
rect 7587 3368 7621 3402
rect 7621 3368 7689 3402
rect 7689 3368 7693 3402
rect 7515 3334 7693 3368
rect 7515 3300 7519 3334
rect 7519 3300 7587 3334
rect 7587 3300 7621 3334
rect 7621 3300 7689 3334
rect 7689 3300 7693 3334
rect 7515 3266 7693 3300
rect 7515 3232 7519 3266
rect 7519 3232 7587 3266
rect 7587 3232 7621 3266
rect 7621 3232 7689 3266
rect 7689 3232 7693 3266
rect 7515 3198 7693 3232
rect 7515 3194 7519 3198
rect 7519 3194 7587 3198
rect 7587 3194 7621 3198
rect 7621 3194 7689 3198
rect 7689 3194 7693 3198
rect 7587 3164 7621 3182
rect 7587 3148 7621 3164
rect 7515 3074 7549 3108
rect 7587 3074 7621 3108
rect 7659 3074 7693 3108
rect 7515 2994 7549 3028
rect 7587 2994 7621 3028
rect 7659 2994 7693 3028
rect 7515 2914 7549 2948
rect 7587 2914 7621 2948
rect 7659 2914 7693 2948
rect 7515 2834 7549 2868
rect 7587 2834 7621 2868
rect 7659 2834 7693 2868
rect 7515 2754 7549 2788
rect 7587 2754 7621 2788
rect 7659 2754 7693 2788
rect 7515 2674 7549 2708
rect 7587 2674 7621 2708
rect 7659 2674 7693 2708
rect 7515 2594 7549 2628
rect 7587 2594 7621 2628
rect 7659 2594 7693 2628
rect 7587 2540 7621 2556
rect 7587 2522 7621 2540
rect 7515 2506 7519 2518
rect 7519 2506 7587 2518
rect 7587 2506 7621 2518
rect 7621 2506 7689 2518
rect 7689 2506 7693 2518
rect 7515 2472 7693 2506
rect 7515 2438 7519 2472
rect 7519 2438 7587 2472
rect 7587 2438 7621 2472
rect 7621 2438 7689 2472
rect 7689 2438 7693 2472
rect 7515 2404 7693 2438
rect 7515 2370 7519 2404
rect 7519 2370 7587 2404
rect 7587 2370 7621 2404
rect 7621 2370 7689 2404
rect 7689 2370 7693 2404
rect 7515 2336 7693 2370
rect 7515 2302 7519 2336
rect 7519 2302 7587 2336
rect 7587 2302 7621 2336
rect 7621 2302 7689 2336
rect 7689 2302 7693 2336
rect 7515 2268 7693 2302
rect 7515 2234 7519 2268
rect 7519 2234 7587 2268
rect 7587 2234 7621 2268
rect 7621 2234 7689 2268
rect 7689 2234 7693 2268
rect 7515 2200 7693 2234
rect 7515 2166 7519 2200
rect 7519 2166 7587 2200
rect 7587 2166 7621 2200
rect 7621 2166 7689 2200
rect 7689 2166 7693 2200
rect 7515 2132 7693 2166
rect 7515 2098 7519 2132
rect 7519 2098 7587 2132
rect 7587 2098 7621 2132
rect 7621 2098 7689 2132
rect 7689 2098 7693 2132
rect 7515 2064 7693 2098
rect 7515 2030 7519 2064
rect 7519 2030 7587 2064
rect 7587 2030 7621 2064
rect 7621 2030 7689 2064
rect 7689 2030 7693 2064
rect 7515 1996 7693 2030
rect 7515 1962 7519 1996
rect 7519 1962 7587 1996
rect 7587 1962 7621 1996
rect 7621 1962 7689 1996
rect 7689 1962 7693 1996
rect 7515 1928 7693 1962
rect 7515 1894 7519 1928
rect 7519 1894 7587 1928
rect 7587 1894 7621 1928
rect 7621 1894 7689 1928
rect 7689 1894 7693 1928
rect 7515 1860 7693 1894
rect 7515 1826 7519 1860
rect 7519 1826 7587 1860
rect 7587 1826 7621 1860
rect 7621 1826 7689 1860
rect 7689 1826 7693 1860
rect 7515 1792 7693 1826
rect 7515 1758 7519 1792
rect 7519 1758 7587 1792
rect 7587 1758 7621 1792
rect 7621 1758 7689 1792
rect 7689 1758 7693 1792
rect 7515 1724 7693 1758
rect 7515 1690 7519 1724
rect 7519 1690 7587 1724
rect 7587 1690 7621 1724
rect 7621 1690 7689 1724
rect 7689 1690 7693 1724
rect 7515 1656 7693 1690
rect 7515 1622 7519 1656
rect 7519 1622 7587 1656
rect 7587 1622 7621 1656
rect 7621 1622 7689 1656
rect 7689 1622 7693 1656
rect 7515 1620 7693 1622
rect 7587 1586 7621 1620
rect 7270 1144 7376 1250
rect 8011 4064 8045 4098
rect 8083 4064 8117 4098
rect 8155 4064 8189 4098
rect 8011 3991 8045 4025
rect 8083 3991 8117 4025
rect 8155 3991 8189 4025
rect 8011 3918 8045 3952
rect 8083 3918 8117 3952
rect 8155 3918 8189 3952
rect 8011 3845 8045 3879
rect 8083 3845 8117 3879
rect 8155 3845 8189 3879
rect 8011 3772 8045 3806
rect 8083 3772 8117 3806
rect 8155 3772 8189 3806
rect 8011 3699 8045 3733
rect 8083 3699 8117 3733
rect 8155 3699 8189 3733
rect 8011 3626 8045 3660
rect 8083 3626 8117 3660
rect 8155 3626 8189 3660
rect 8011 3553 8045 3587
rect 8083 3553 8117 3587
rect 8155 3553 8189 3587
rect 8011 3480 8045 3514
rect 8083 3480 8117 3514
rect 8155 3480 8189 3514
rect 8011 3407 8045 3441
rect 8083 3407 8117 3441
rect 8155 3407 8189 3441
rect 8011 3334 8045 3368
rect 8083 3334 8117 3368
rect 8155 3334 8189 3368
rect 8011 3261 8045 3295
rect 8083 3261 8117 3295
rect 8155 3261 8189 3295
rect 8011 3188 8045 3222
rect 8083 3188 8117 3222
rect 8155 3188 8189 3222
rect 8011 3115 8045 3149
rect 8083 3115 8117 3149
rect 8155 3115 8189 3149
rect 8011 3042 8045 3076
rect 8083 3042 8117 3076
rect 8155 3042 8189 3076
rect 8011 2969 8045 3003
rect 8083 2969 8117 3003
rect 8155 2969 8189 3003
rect 8011 2896 8045 2930
rect 8083 2896 8117 2930
rect 8155 2896 8189 2930
rect 8011 2823 8045 2857
rect 8083 2823 8117 2857
rect 8155 2823 8189 2857
rect 8011 2750 8045 2784
rect 8083 2750 8117 2784
rect 8155 2750 8189 2784
rect 8011 2677 8045 2711
rect 8083 2677 8117 2711
rect 8155 2677 8189 2711
rect 8011 2604 8045 2638
rect 8083 2604 8117 2638
rect 8155 2604 8189 2638
rect 8011 2531 8045 2565
rect 8083 2531 8117 2565
rect 8155 2531 8189 2565
rect 8011 2458 8045 2492
rect 8083 2458 8117 2492
rect 8155 2458 8189 2492
rect 8011 2385 8045 2419
rect 8083 2385 8117 2419
rect 8155 2385 8189 2419
rect 8011 2312 8045 2346
rect 8083 2312 8117 2346
rect 8155 2312 8189 2346
rect 8011 2239 8045 2273
rect 8083 2239 8117 2273
rect 8155 2239 8189 2273
rect 8011 2166 8045 2200
rect 8083 2166 8117 2200
rect 8155 2166 8189 2200
rect 8011 2092 8045 2126
rect 8083 2092 8117 2126
rect 8155 2092 8189 2126
rect 8011 2018 8045 2052
rect 8083 2018 8117 2052
rect 8155 2018 8189 2052
rect 8011 1944 8045 1978
rect 8083 1944 8117 1978
rect 8155 1944 8189 1978
rect 8011 1870 8045 1904
rect 8083 1870 8117 1904
rect 8155 1870 8189 1904
rect 8011 1796 8045 1830
rect 8083 1796 8117 1830
rect 8155 1796 8189 1830
rect 8011 1722 8045 1756
rect 8083 1722 8117 1756
rect 8155 1722 8189 1756
rect 8011 1648 8045 1682
rect 8083 1648 8117 1682
rect 8155 1648 8189 1682
rect 8011 1574 8045 1608
rect 8083 1574 8117 1608
rect 8155 1574 8189 1608
rect 7832 1144 7938 1250
rect 8579 4092 8613 4118
rect 8507 4082 8685 4092
rect 8507 4048 8511 4082
rect 8511 4048 8579 4082
rect 8579 4048 8613 4082
rect 8613 4048 8681 4082
rect 8681 4048 8685 4082
rect 8507 4014 8685 4048
rect 8507 3980 8511 4014
rect 8511 3980 8579 4014
rect 8579 3980 8613 4014
rect 8613 3980 8681 4014
rect 8681 3980 8685 4014
rect 8507 3946 8685 3980
rect 8507 3912 8511 3946
rect 8511 3912 8579 3946
rect 8579 3912 8613 3946
rect 8613 3912 8681 3946
rect 8681 3912 8685 3946
rect 8507 3878 8685 3912
rect 8507 3844 8511 3878
rect 8511 3844 8579 3878
rect 8579 3844 8613 3878
rect 8613 3844 8681 3878
rect 8681 3844 8685 3878
rect 8507 3810 8685 3844
rect 8507 3776 8511 3810
rect 8511 3776 8579 3810
rect 8579 3776 8613 3810
rect 8613 3776 8681 3810
rect 8681 3776 8685 3810
rect 8507 3742 8685 3776
rect 8507 3708 8511 3742
rect 8511 3708 8579 3742
rect 8579 3708 8613 3742
rect 8613 3708 8681 3742
rect 8681 3708 8685 3742
rect 8507 3674 8685 3708
rect 8507 3640 8511 3674
rect 8511 3640 8579 3674
rect 8579 3640 8613 3674
rect 8613 3640 8681 3674
rect 8681 3640 8685 3674
rect 8507 3606 8685 3640
rect 8507 3572 8511 3606
rect 8511 3572 8579 3606
rect 8579 3572 8613 3606
rect 8613 3572 8681 3606
rect 8681 3572 8685 3606
rect 8507 3538 8685 3572
rect 8507 3504 8511 3538
rect 8511 3504 8579 3538
rect 8579 3504 8613 3538
rect 8613 3504 8681 3538
rect 8681 3504 8685 3538
rect 8507 3470 8685 3504
rect 8507 3436 8511 3470
rect 8511 3436 8579 3470
rect 8579 3436 8613 3470
rect 8613 3436 8681 3470
rect 8681 3436 8685 3470
rect 8507 3402 8685 3436
rect 8507 3368 8511 3402
rect 8511 3368 8579 3402
rect 8579 3368 8613 3402
rect 8613 3368 8681 3402
rect 8681 3368 8685 3402
rect 8507 3334 8685 3368
rect 8507 3300 8511 3334
rect 8511 3300 8579 3334
rect 8579 3300 8613 3334
rect 8613 3300 8681 3334
rect 8681 3300 8685 3334
rect 8507 3266 8685 3300
rect 8507 3232 8511 3266
rect 8511 3232 8579 3266
rect 8579 3232 8613 3266
rect 8613 3232 8681 3266
rect 8681 3232 8685 3266
rect 8507 3198 8685 3232
rect 8507 3194 8511 3198
rect 8511 3194 8579 3198
rect 8579 3194 8613 3198
rect 8613 3194 8681 3198
rect 8681 3194 8685 3198
rect 8579 3164 8613 3182
rect 8579 3148 8613 3164
rect 8507 3074 8541 3108
rect 8579 3074 8613 3108
rect 8651 3074 8685 3108
rect 8507 2994 8541 3028
rect 8579 2994 8613 3028
rect 8651 2994 8685 3028
rect 8507 2914 8541 2948
rect 8579 2914 8613 2948
rect 8651 2914 8685 2948
rect 8507 2834 8541 2868
rect 8579 2834 8613 2868
rect 8651 2834 8685 2868
rect 8507 2754 8541 2788
rect 8579 2754 8613 2788
rect 8651 2754 8685 2788
rect 8507 2674 8541 2708
rect 8579 2674 8613 2708
rect 8651 2674 8685 2708
rect 8507 2594 8541 2628
rect 8579 2594 8613 2628
rect 8651 2594 8685 2628
rect 8579 2540 8613 2556
rect 8579 2522 8613 2540
rect 8507 2506 8511 2518
rect 8511 2506 8579 2518
rect 8579 2506 8613 2518
rect 8613 2506 8681 2518
rect 8681 2506 8685 2518
rect 8507 2472 8685 2506
rect 8507 2438 8511 2472
rect 8511 2438 8579 2472
rect 8579 2438 8613 2472
rect 8613 2438 8681 2472
rect 8681 2438 8685 2472
rect 8507 2404 8685 2438
rect 8507 2370 8511 2404
rect 8511 2370 8579 2404
rect 8579 2370 8613 2404
rect 8613 2370 8681 2404
rect 8681 2370 8685 2404
rect 8507 2336 8685 2370
rect 8507 2302 8511 2336
rect 8511 2302 8579 2336
rect 8579 2302 8613 2336
rect 8613 2302 8681 2336
rect 8681 2302 8685 2336
rect 8507 2268 8685 2302
rect 8507 2234 8511 2268
rect 8511 2234 8579 2268
rect 8579 2234 8613 2268
rect 8613 2234 8681 2268
rect 8681 2234 8685 2268
rect 8507 2200 8685 2234
rect 8507 2166 8511 2200
rect 8511 2166 8579 2200
rect 8579 2166 8613 2200
rect 8613 2166 8681 2200
rect 8681 2166 8685 2200
rect 8507 2132 8685 2166
rect 8507 2098 8511 2132
rect 8511 2098 8579 2132
rect 8579 2098 8613 2132
rect 8613 2098 8681 2132
rect 8681 2098 8685 2132
rect 8507 2064 8685 2098
rect 8507 2030 8511 2064
rect 8511 2030 8579 2064
rect 8579 2030 8613 2064
rect 8613 2030 8681 2064
rect 8681 2030 8685 2064
rect 8507 1996 8685 2030
rect 8507 1962 8511 1996
rect 8511 1962 8579 1996
rect 8579 1962 8613 1996
rect 8613 1962 8681 1996
rect 8681 1962 8685 1996
rect 8507 1928 8685 1962
rect 8507 1894 8511 1928
rect 8511 1894 8579 1928
rect 8579 1894 8613 1928
rect 8613 1894 8681 1928
rect 8681 1894 8685 1928
rect 8507 1860 8685 1894
rect 8507 1826 8511 1860
rect 8511 1826 8579 1860
rect 8579 1826 8613 1860
rect 8613 1826 8681 1860
rect 8681 1826 8685 1860
rect 8507 1792 8685 1826
rect 8507 1758 8511 1792
rect 8511 1758 8579 1792
rect 8579 1758 8613 1792
rect 8613 1758 8681 1792
rect 8681 1758 8685 1792
rect 8507 1724 8685 1758
rect 8507 1690 8511 1724
rect 8511 1690 8579 1724
rect 8579 1690 8613 1724
rect 8613 1690 8681 1724
rect 8681 1690 8685 1724
rect 8507 1656 8685 1690
rect 8507 1622 8511 1656
rect 8511 1622 8579 1656
rect 8579 1622 8613 1656
rect 8613 1622 8681 1656
rect 8681 1622 8685 1656
rect 8507 1620 8685 1622
rect 8579 1586 8613 1620
rect 8262 1144 8368 1250
rect 9003 4064 9037 4098
rect 9075 4064 9109 4098
rect 9147 4064 9181 4098
rect 9003 3991 9037 4025
rect 9075 3991 9109 4025
rect 9147 3991 9181 4025
rect 9003 3918 9037 3952
rect 9075 3918 9109 3952
rect 9147 3918 9181 3952
rect 9003 3845 9037 3879
rect 9075 3845 9109 3879
rect 9147 3845 9181 3879
rect 9003 3772 9037 3806
rect 9075 3772 9109 3806
rect 9147 3772 9181 3806
rect 9003 3699 9037 3733
rect 9075 3699 9109 3733
rect 9147 3699 9181 3733
rect 9003 3626 9037 3660
rect 9075 3626 9109 3660
rect 9147 3626 9181 3660
rect 9003 3553 9037 3587
rect 9075 3553 9109 3587
rect 9147 3553 9181 3587
rect 9003 3480 9037 3514
rect 9075 3480 9109 3514
rect 9147 3480 9181 3514
rect 9003 3407 9037 3441
rect 9075 3407 9109 3441
rect 9147 3407 9181 3441
rect 9003 3334 9037 3368
rect 9075 3334 9109 3368
rect 9147 3334 9181 3368
rect 9003 3261 9037 3295
rect 9075 3261 9109 3295
rect 9147 3261 9181 3295
rect 9003 3188 9037 3222
rect 9075 3188 9109 3222
rect 9147 3188 9181 3222
rect 9003 3115 9037 3149
rect 9075 3115 9109 3149
rect 9147 3115 9181 3149
rect 9003 3042 9037 3076
rect 9075 3042 9109 3076
rect 9147 3042 9181 3076
rect 9003 2969 9037 3003
rect 9075 2969 9109 3003
rect 9147 2969 9181 3003
rect 9003 2896 9037 2930
rect 9075 2896 9109 2930
rect 9147 2896 9181 2930
rect 9003 2823 9037 2857
rect 9075 2823 9109 2857
rect 9147 2823 9181 2857
rect 9003 2750 9037 2784
rect 9075 2750 9109 2784
rect 9147 2750 9181 2784
rect 9003 2677 9037 2711
rect 9075 2677 9109 2711
rect 9147 2677 9181 2711
rect 9003 2604 9037 2638
rect 9075 2604 9109 2638
rect 9147 2604 9181 2638
rect 9003 2531 9037 2565
rect 9075 2531 9109 2565
rect 9147 2531 9181 2565
rect 9003 2458 9037 2492
rect 9075 2458 9109 2492
rect 9147 2458 9181 2492
rect 9003 2385 9037 2419
rect 9075 2385 9109 2419
rect 9147 2385 9181 2419
rect 9003 2312 9037 2346
rect 9075 2312 9109 2346
rect 9147 2312 9181 2346
rect 9003 2239 9037 2273
rect 9075 2239 9109 2273
rect 9147 2239 9181 2273
rect 9003 2166 9037 2200
rect 9075 2166 9109 2200
rect 9147 2166 9181 2200
rect 9003 2092 9037 2126
rect 9075 2092 9109 2126
rect 9147 2092 9181 2126
rect 9003 2018 9037 2052
rect 9075 2018 9109 2052
rect 9147 2018 9181 2052
rect 9003 1944 9037 1978
rect 9075 1944 9109 1978
rect 9147 1944 9181 1978
rect 9003 1870 9037 1904
rect 9075 1870 9109 1904
rect 9147 1870 9181 1904
rect 9003 1796 9037 1830
rect 9075 1796 9109 1830
rect 9147 1796 9181 1830
rect 9003 1722 9037 1756
rect 9075 1722 9109 1756
rect 9147 1722 9181 1756
rect 9003 1648 9037 1682
rect 9075 1648 9109 1682
rect 9147 1648 9181 1682
rect 9003 1574 9037 1608
rect 9075 1574 9109 1608
rect 9147 1574 9181 1608
rect 8824 1144 8930 1250
rect 9571 4092 9605 4118
rect 9499 4082 9677 4092
rect 9499 4048 9503 4082
rect 9503 4048 9571 4082
rect 9571 4048 9605 4082
rect 9605 4048 9673 4082
rect 9673 4048 9677 4082
rect 9499 4014 9677 4048
rect 9499 3980 9503 4014
rect 9503 3980 9571 4014
rect 9571 3980 9605 4014
rect 9605 3980 9673 4014
rect 9673 3980 9677 4014
rect 9499 3946 9677 3980
rect 9499 3912 9503 3946
rect 9503 3912 9571 3946
rect 9571 3912 9605 3946
rect 9605 3912 9673 3946
rect 9673 3912 9677 3946
rect 9499 3878 9677 3912
rect 9499 3844 9503 3878
rect 9503 3844 9571 3878
rect 9571 3844 9605 3878
rect 9605 3844 9673 3878
rect 9673 3844 9677 3878
rect 9499 3810 9677 3844
rect 9499 3776 9503 3810
rect 9503 3776 9571 3810
rect 9571 3776 9605 3810
rect 9605 3776 9673 3810
rect 9673 3776 9677 3810
rect 9499 3742 9677 3776
rect 9499 3708 9503 3742
rect 9503 3708 9571 3742
rect 9571 3708 9605 3742
rect 9605 3708 9673 3742
rect 9673 3708 9677 3742
rect 9499 3674 9677 3708
rect 9499 3640 9503 3674
rect 9503 3640 9571 3674
rect 9571 3640 9605 3674
rect 9605 3640 9673 3674
rect 9673 3640 9677 3674
rect 9499 3606 9677 3640
rect 9499 3572 9503 3606
rect 9503 3572 9571 3606
rect 9571 3572 9605 3606
rect 9605 3572 9673 3606
rect 9673 3572 9677 3606
rect 9499 3538 9677 3572
rect 9499 3504 9503 3538
rect 9503 3504 9571 3538
rect 9571 3504 9605 3538
rect 9605 3504 9673 3538
rect 9673 3504 9677 3538
rect 9499 3470 9677 3504
rect 9499 3436 9503 3470
rect 9503 3436 9571 3470
rect 9571 3436 9605 3470
rect 9605 3436 9673 3470
rect 9673 3436 9677 3470
rect 9499 3402 9677 3436
rect 9499 3368 9503 3402
rect 9503 3368 9571 3402
rect 9571 3368 9605 3402
rect 9605 3368 9673 3402
rect 9673 3368 9677 3402
rect 9499 3334 9677 3368
rect 9499 3300 9503 3334
rect 9503 3300 9571 3334
rect 9571 3300 9605 3334
rect 9605 3300 9673 3334
rect 9673 3300 9677 3334
rect 9499 3266 9677 3300
rect 9499 3232 9503 3266
rect 9503 3232 9571 3266
rect 9571 3232 9605 3266
rect 9605 3232 9673 3266
rect 9673 3232 9677 3266
rect 9499 3198 9677 3232
rect 9499 3194 9503 3198
rect 9503 3194 9571 3198
rect 9571 3194 9605 3198
rect 9605 3194 9673 3198
rect 9673 3194 9677 3198
rect 9571 3164 9605 3182
rect 9571 3148 9605 3164
rect 9499 3074 9533 3108
rect 9571 3074 9605 3108
rect 9643 3074 9677 3108
rect 9499 2994 9533 3028
rect 9571 2994 9605 3028
rect 9643 2994 9677 3028
rect 9499 2914 9533 2948
rect 9571 2914 9605 2948
rect 9643 2914 9677 2948
rect 9499 2834 9533 2868
rect 9571 2834 9605 2868
rect 9643 2834 9677 2868
rect 9499 2754 9533 2788
rect 9571 2754 9605 2788
rect 9643 2754 9677 2788
rect 9499 2674 9533 2708
rect 9571 2674 9605 2708
rect 9643 2674 9677 2708
rect 9499 2594 9533 2628
rect 9571 2594 9605 2628
rect 9643 2594 9677 2628
rect 9571 2540 9605 2556
rect 9571 2522 9605 2540
rect 9499 2506 9503 2518
rect 9503 2506 9571 2518
rect 9571 2506 9605 2518
rect 9605 2506 9673 2518
rect 9673 2506 9677 2518
rect 9499 2472 9677 2506
rect 9499 2438 9503 2472
rect 9503 2438 9571 2472
rect 9571 2438 9605 2472
rect 9605 2438 9673 2472
rect 9673 2438 9677 2472
rect 9499 2404 9677 2438
rect 9499 2370 9503 2404
rect 9503 2370 9571 2404
rect 9571 2370 9605 2404
rect 9605 2370 9673 2404
rect 9673 2370 9677 2404
rect 9499 2336 9677 2370
rect 9499 2302 9503 2336
rect 9503 2302 9571 2336
rect 9571 2302 9605 2336
rect 9605 2302 9673 2336
rect 9673 2302 9677 2336
rect 9499 2268 9677 2302
rect 9499 2234 9503 2268
rect 9503 2234 9571 2268
rect 9571 2234 9605 2268
rect 9605 2234 9673 2268
rect 9673 2234 9677 2268
rect 9499 2200 9677 2234
rect 9499 2166 9503 2200
rect 9503 2166 9571 2200
rect 9571 2166 9605 2200
rect 9605 2166 9673 2200
rect 9673 2166 9677 2200
rect 9499 2132 9677 2166
rect 9499 2098 9503 2132
rect 9503 2098 9571 2132
rect 9571 2098 9605 2132
rect 9605 2098 9673 2132
rect 9673 2098 9677 2132
rect 9499 2064 9677 2098
rect 9499 2030 9503 2064
rect 9503 2030 9571 2064
rect 9571 2030 9605 2064
rect 9605 2030 9673 2064
rect 9673 2030 9677 2064
rect 9499 1996 9677 2030
rect 9499 1962 9503 1996
rect 9503 1962 9571 1996
rect 9571 1962 9605 1996
rect 9605 1962 9673 1996
rect 9673 1962 9677 1996
rect 9499 1928 9677 1962
rect 9499 1894 9503 1928
rect 9503 1894 9571 1928
rect 9571 1894 9605 1928
rect 9605 1894 9673 1928
rect 9673 1894 9677 1928
rect 9499 1860 9677 1894
rect 9499 1826 9503 1860
rect 9503 1826 9571 1860
rect 9571 1826 9605 1860
rect 9605 1826 9673 1860
rect 9673 1826 9677 1860
rect 9499 1792 9677 1826
rect 9499 1758 9503 1792
rect 9503 1758 9571 1792
rect 9571 1758 9605 1792
rect 9605 1758 9673 1792
rect 9673 1758 9677 1792
rect 9499 1724 9677 1758
rect 9499 1690 9503 1724
rect 9503 1690 9571 1724
rect 9571 1690 9605 1724
rect 9605 1690 9673 1724
rect 9673 1690 9677 1724
rect 9499 1656 9677 1690
rect 9499 1622 9503 1656
rect 9503 1622 9571 1656
rect 9571 1622 9605 1656
rect 9605 1622 9673 1656
rect 9673 1622 9677 1656
rect 9499 1620 9677 1622
rect 9571 1586 9605 1620
rect 9254 1144 9360 1250
rect 9995 4064 10029 4098
rect 10067 4064 10101 4098
rect 10139 4064 10173 4098
rect 9995 3991 10029 4025
rect 10067 3991 10101 4025
rect 10139 3991 10173 4025
rect 9995 3918 10029 3952
rect 10067 3918 10101 3952
rect 10139 3918 10173 3952
rect 9995 3845 10029 3879
rect 10067 3845 10101 3879
rect 10139 3845 10173 3879
rect 9995 3772 10029 3806
rect 10067 3772 10101 3806
rect 10139 3772 10173 3806
rect 9995 3699 10029 3733
rect 10067 3699 10101 3733
rect 10139 3699 10173 3733
rect 9995 3626 10029 3660
rect 10067 3626 10101 3660
rect 10139 3626 10173 3660
rect 9995 3553 10029 3587
rect 10067 3553 10101 3587
rect 10139 3553 10173 3587
rect 9995 3480 10029 3514
rect 10067 3480 10101 3514
rect 10139 3480 10173 3514
rect 9995 3407 10029 3441
rect 10067 3407 10101 3441
rect 10139 3407 10173 3441
rect 9995 3334 10029 3368
rect 10067 3334 10101 3368
rect 10139 3334 10173 3368
rect 9995 3261 10029 3295
rect 10067 3261 10101 3295
rect 10139 3261 10173 3295
rect 9995 3188 10029 3222
rect 10067 3188 10101 3222
rect 10139 3188 10173 3222
rect 9995 3115 10029 3149
rect 10067 3115 10101 3149
rect 10139 3115 10173 3149
rect 9995 3042 10029 3076
rect 10067 3042 10101 3076
rect 10139 3042 10173 3076
rect 9995 2969 10029 3003
rect 10067 2969 10101 3003
rect 10139 2969 10173 3003
rect 9995 2896 10029 2930
rect 10067 2896 10101 2930
rect 10139 2896 10173 2930
rect 9995 2823 10029 2857
rect 10067 2823 10101 2857
rect 10139 2823 10173 2857
rect 9995 2750 10029 2784
rect 10067 2750 10101 2784
rect 10139 2750 10173 2784
rect 9995 2677 10029 2711
rect 10067 2677 10101 2711
rect 10139 2677 10173 2711
rect 9995 2604 10029 2638
rect 10067 2604 10101 2638
rect 10139 2604 10173 2638
rect 9995 2531 10029 2565
rect 10067 2531 10101 2565
rect 10139 2531 10173 2565
rect 9995 2458 10029 2492
rect 10067 2458 10101 2492
rect 10139 2458 10173 2492
rect 9995 2385 10029 2419
rect 10067 2385 10101 2419
rect 10139 2385 10173 2419
rect 9995 2312 10029 2346
rect 10067 2312 10101 2346
rect 10139 2312 10173 2346
rect 9995 2239 10029 2273
rect 10067 2239 10101 2273
rect 10139 2239 10173 2273
rect 9995 2166 10029 2200
rect 10067 2166 10101 2200
rect 10139 2166 10173 2200
rect 9995 2092 10029 2126
rect 10067 2092 10101 2126
rect 10139 2092 10173 2126
rect 9995 2018 10029 2052
rect 10067 2018 10101 2052
rect 10139 2018 10173 2052
rect 9995 1944 10029 1978
rect 10067 1944 10101 1978
rect 10139 1944 10173 1978
rect 9995 1870 10029 1904
rect 10067 1870 10101 1904
rect 10139 1870 10173 1904
rect 9995 1796 10029 1830
rect 10067 1796 10101 1830
rect 10139 1796 10173 1830
rect 9995 1722 10029 1756
rect 10067 1722 10101 1756
rect 10139 1722 10173 1756
rect 9995 1648 10029 1682
rect 10067 1648 10101 1682
rect 10139 1648 10173 1682
rect 9995 1574 10029 1608
rect 10067 1574 10101 1608
rect 10139 1574 10173 1608
rect 9816 1144 9922 1250
rect 10563 4092 10597 4118
rect 10491 4082 10669 4092
rect 10491 4048 10495 4082
rect 10495 4048 10563 4082
rect 10563 4048 10597 4082
rect 10597 4048 10665 4082
rect 10665 4048 10669 4082
rect 10491 4014 10669 4048
rect 10491 3980 10495 4014
rect 10495 3980 10563 4014
rect 10563 3980 10597 4014
rect 10597 3980 10665 4014
rect 10665 3980 10669 4014
rect 10491 3946 10669 3980
rect 10491 3912 10495 3946
rect 10495 3912 10563 3946
rect 10563 3912 10597 3946
rect 10597 3912 10665 3946
rect 10665 3912 10669 3946
rect 10491 3878 10669 3912
rect 10491 3844 10495 3878
rect 10495 3844 10563 3878
rect 10563 3844 10597 3878
rect 10597 3844 10665 3878
rect 10665 3844 10669 3878
rect 10491 3810 10669 3844
rect 10491 3776 10495 3810
rect 10495 3776 10563 3810
rect 10563 3776 10597 3810
rect 10597 3776 10665 3810
rect 10665 3776 10669 3810
rect 10491 3742 10669 3776
rect 10491 3708 10495 3742
rect 10495 3708 10563 3742
rect 10563 3708 10597 3742
rect 10597 3708 10665 3742
rect 10665 3708 10669 3742
rect 10491 3674 10669 3708
rect 10491 3640 10495 3674
rect 10495 3640 10563 3674
rect 10563 3640 10597 3674
rect 10597 3640 10665 3674
rect 10665 3640 10669 3674
rect 10491 3606 10669 3640
rect 10491 3572 10495 3606
rect 10495 3572 10563 3606
rect 10563 3572 10597 3606
rect 10597 3572 10665 3606
rect 10665 3572 10669 3606
rect 10491 3538 10669 3572
rect 10491 3504 10495 3538
rect 10495 3504 10563 3538
rect 10563 3504 10597 3538
rect 10597 3504 10665 3538
rect 10665 3504 10669 3538
rect 10491 3470 10669 3504
rect 10491 3436 10495 3470
rect 10495 3436 10563 3470
rect 10563 3436 10597 3470
rect 10597 3436 10665 3470
rect 10665 3436 10669 3470
rect 10491 3402 10669 3436
rect 10491 3368 10495 3402
rect 10495 3368 10563 3402
rect 10563 3368 10597 3402
rect 10597 3368 10665 3402
rect 10665 3368 10669 3402
rect 10491 3334 10669 3368
rect 10491 3300 10495 3334
rect 10495 3300 10563 3334
rect 10563 3300 10597 3334
rect 10597 3300 10665 3334
rect 10665 3300 10669 3334
rect 10491 3266 10669 3300
rect 10491 3232 10495 3266
rect 10495 3232 10563 3266
rect 10563 3232 10597 3266
rect 10597 3232 10665 3266
rect 10665 3232 10669 3266
rect 10491 3198 10669 3232
rect 10491 3194 10495 3198
rect 10495 3194 10563 3198
rect 10563 3194 10597 3198
rect 10597 3194 10665 3198
rect 10665 3194 10669 3198
rect 10563 3164 10597 3182
rect 10563 3148 10597 3164
rect 10491 3074 10525 3108
rect 10563 3074 10597 3108
rect 10635 3074 10669 3108
rect 10491 2994 10525 3028
rect 10563 2994 10597 3028
rect 10635 2994 10669 3028
rect 10491 2914 10525 2948
rect 10563 2914 10597 2948
rect 10635 2914 10669 2948
rect 10491 2834 10525 2868
rect 10563 2834 10597 2868
rect 10635 2834 10669 2868
rect 10491 2754 10525 2788
rect 10563 2754 10597 2788
rect 10635 2754 10669 2788
rect 10491 2674 10525 2708
rect 10563 2674 10597 2708
rect 10635 2674 10669 2708
rect 10491 2594 10525 2628
rect 10563 2594 10597 2628
rect 10635 2594 10669 2628
rect 10563 2540 10597 2556
rect 10563 2522 10597 2540
rect 10491 2506 10495 2518
rect 10495 2506 10563 2518
rect 10563 2506 10597 2518
rect 10597 2506 10665 2518
rect 10665 2506 10669 2518
rect 10491 2472 10669 2506
rect 10491 2438 10495 2472
rect 10495 2438 10563 2472
rect 10563 2438 10597 2472
rect 10597 2438 10665 2472
rect 10665 2438 10669 2472
rect 10491 2404 10669 2438
rect 10491 2370 10495 2404
rect 10495 2370 10563 2404
rect 10563 2370 10597 2404
rect 10597 2370 10665 2404
rect 10665 2370 10669 2404
rect 10491 2336 10669 2370
rect 10491 2302 10495 2336
rect 10495 2302 10563 2336
rect 10563 2302 10597 2336
rect 10597 2302 10665 2336
rect 10665 2302 10669 2336
rect 10491 2268 10669 2302
rect 10491 2234 10495 2268
rect 10495 2234 10563 2268
rect 10563 2234 10597 2268
rect 10597 2234 10665 2268
rect 10665 2234 10669 2268
rect 10491 2200 10669 2234
rect 10491 2166 10495 2200
rect 10495 2166 10563 2200
rect 10563 2166 10597 2200
rect 10597 2166 10665 2200
rect 10665 2166 10669 2200
rect 10491 2132 10669 2166
rect 10491 2098 10495 2132
rect 10495 2098 10563 2132
rect 10563 2098 10597 2132
rect 10597 2098 10665 2132
rect 10665 2098 10669 2132
rect 10491 2064 10669 2098
rect 10491 2030 10495 2064
rect 10495 2030 10563 2064
rect 10563 2030 10597 2064
rect 10597 2030 10665 2064
rect 10665 2030 10669 2064
rect 10491 1996 10669 2030
rect 10491 1962 10495 1996
rect 10495 1962 10563 1996
rect 10563 1962 10597 1996
rect 10597 1962 10665 1996
rect 10665 1962 10669 1996
rect 10491 1928 10669 1962
rect 10491 1894 10495 1928
rect 10495 1894 10563 1928
rect 10563 1894 10597 1928
rect 10597 1894 10665 1928
rect 10665 1894 10669 1928
rect 10491 1860 10669 1894
rect 10491 1826 10495 1860
rect 10495 1826 10563 1860
rect 10563 1826 10597 1860
rect 10597 1826 10665 1860
rect 10665 1826 10669 1860
rect 10491 1792 10669 1826
rect 10491 1758 10495 1792
rect 10495 1758 10563 1792
rect 10563 1758 10597 1792
rect 10597 1758 10665 1792
rect 10665 1758 10669 1792
rect 10491 1724 10669 1758
rect 10491 1690 10495 1724
rect 10495 1690 10563 1724
rect 10563 1690 10597 1724
rect 10597 1690 10665 1724
rect 10665 1690 10669 1724
rect 10491 1656 10669 1690
rect 10491 1622 10495 1656
rect 10495 1622 10563 1656
rect 10563 1622 10597 1656
rect 10597 1622 10665 1656
rect 10665 1622 10669 1656
rect 10491 1620 10669 1622
rect 10563 1586 10597 1620
rect 10246 1144 10352 1250
rect 10987 4064 11021 4098
rect 11059 4064 11093 4098
rect 11131 4064 11165 4098
rect 10987 3991 11021 4025
rect 11059 3991 11093 4025
rect 11131 3991 11165 4025
rect 10987 3918 11021 3952
rect 11059 3918 11093 3952
rect 11131 3918 11165 3952
rect 10987 3845 11021 3879
rect 11059 3845 11093 3879
rect 11131 3845 11165 3879
rect 10987 3772 11021 3806
rect 11059 3772 11093 3806
rect 11131 3772 11165 3806
rect 10987 3699 11021 3733
rect 11059 3699 11093 3733
rect 11131 3699 11165 3733
rect 10987 3626 11021 3660
rect 11059 3626 11093 3660
rect 11131 3626 11165 3660
rect 10987 3553 11021 3587
rect 11059 3553 11093 3587
rect 11131 3553 11165 3587
rect 10987 3480 11021 3514
rect 11059 3480 11093 3514
rect 11131 3480 11165 3514
rect 10987 3407 11021 3441
rect 11059 3407 11093 3441
rect 11131 3407 11165 3441
rect 10987 3334 11021 3368
rect 11059 3334 11093 3368
rect 11131 3334 11165 3368
rect 10987 3261 11021 3295
rect 11059 3261 11093 3295
rect 11131 3261 11165 3295
rect 10987 3188 11021 3222
rect 11059 3188 11093 3222
rect 11131 3188 11165 3222
rect 10987 3115 11021 3149
rect 11059 3115 11093 3149
rect 11131 3115 11165 3149
rect 10987 3042 11021 3076
rect 11059 3042 11093 3076
rect 11131 3042 11165 3076
rect 10987 2969 11021 3003
rect 11059 2969 11093 3003
rect 11131 2969 11165 3003
rect 10987 2896 11021 2930
rect 11059 2896 11093 2930
rect 11131 2896 11165 2930
rect 10987 2823 11021 2857
rect 11059 2823 11093 2857
rect 11131 2823 11165 2857
rect 10987 2750 11021 2784
rect 11059 2750 11093 2784
rect 11131 2750 11165 2784
rect 10987 2677 11021 2711
rect 11059 2677 11093 2711
rect 11131 2677 11165 2711
rect 10987 2604 11021 2638
rect 11059 2604 11093 2638
rect 11131 2604 11165 2638
rect 10987 2531 11021 2565
rect 11059 2531 11093 2565
rect 11131 2531 11165 2565
rect 10987 2458 11021 2492
rect 11059 2458 11093 2492
rect 11131 2458 11165 2492
rect 10987 2385 11021 2419
rect 11059 2385 11093 2419
rect 11131 2385 11165 2419
rect 10987 2312 11021 2346
rect 11059 2312 11093 2346
rect 11131 2312 11165 2346
rect 10987 2239 11021 2273
rect 11059 2239 11093 2273
rect 11131 2239 11165 2273
rect 10987 2166 11021 2200
rect 11059 2166 11093 2200
rect 11131 2166 11165 2200
rect 10987 2092 11021 2126
rect 11059 2092 11093 2126
rect 11131 2092 11165 2126
rect 10987 2018 11021 2052
rect 11059 2018 11093 2052
rect 11131 2018 11165 2052
rect 10987 1944 11021 1978
rect 11059 1944 11093 1978
rect 11131 1944 11165 1978
rect 10987 1870 11021 1904
rect 11059 1870 11093 1904
rect 11131 1870 11165 1904
rect 10987 1796 11021 1830
rect 11059 1796 11093 1830
rect 11131 1796 11165 1830
rect 10987 1722 11021 1756
rect 11059 1722 11093 1756
rect 11131 1722 11165 1756
rect 10987 1648 11021 1682
rect 11059 1648 11093 1682
rect 11131 1648 11165 1682
rect 10987 1574 11021 1608
rect 11059 1574 11093 1608
rect 11131 1574 11165 1608
rect 10808 1144 10914 1250
rect 11555 4092 11589 4118
rect 11483 4082 11661 4092
rect 11483 4048 11487 4082
rect 11487 4048 11555 4082
rect 11555 4048 11589 4082
rect 11589 4048 11657 4082
rect 11657 4048 11661 4082
rect 11483 4014 11661 4048
rect 11483 3980 11487 4014
rect 11487 3980 11555 4014
rect 11555 3980 11589 4014
rect 11589 3980 11657 4014
rect 11657 3980 11661 4014
rect 11483 3946 11661 3980
rect 11483 3912 11487 3946
rect 11487 3912 11555 3946
rect 11555 3912 11589 3946
rect 11589 3912 11657 3946
rect 11657 3912 11661 3946
rect 11483 3878 11661 3912
rect 11483 3844 11487 3878
rect 11487 3844 11555 3878
rect 11555 3844 11589 3878
rect 11589 3844 11657 3878
rect 11657 3844 11661 3878
rect 11483 3810 11661 3844
rect 11483 3776 11487 3810
rect 11487 3776 11555 3810
rect 11555 3776 11589 3810
rect 11589 3776 11657 3810
rect 11657 3776 11661 3810
rect 11483 3742 11661 3776
rect 11483 3708 11487 3742
rect 11487 3708 11555 3742
rect 11555 3708 11589 3742
rect 11589 3708 11657 3742
rect 11657 3708 11661 3742
rect 11483 3674 11661 3708
rect 11483 3640 11487 3674
rect 11487 3640 11555 3674
rect 11555 3640 11589 3674
rect 11589 3640 11657 3674
rect 11657 3640 11661 3674
rect 11483 3606 11661 3640
rect 11483 3572 11487 3606
rect 11487 3572 11555 3606
rect 11555 3572 11589 3606
rect 11589 3572 11657 3606
rect 11657 3572 11661 3606
rect 11483 3538 11661 3572
rect 11483 3504 11487 3538
rect 11487 3504 11555 3538
rect 11555 3504 11589 3538
rect 11589 3504 11657 3538
rect 11657 3504 11661 3538
rect 11483 3470 11661 3504
rect 11483 3436 11487 3470
rect 11487 3436 11555 3470
rect 11555 3436 11589 3470
rect 11589 3436 11657 3470
rect 11657 3436 11661 3470
rect 11483 3402 11661 3436
rect 11483 3368 11487 3402
rect 11487 3368 11555 3402
rect 11555 3368 11589 3402
rect 11589 3368 11657 3402
rect 11657 3368 11661 3402
rect 11483 3334 11661 3368
rect 11483 3300 11487 3334
rect 11487 3300 11555 3334
rect 11555 3300 11589 3334
rect 11589 3300 11657 3334
rect 11657 3300 11661 3334
rect 11483 3266 11661 3300
rect 11483 3232 11487 3266
rect 11487 3232 11555 3266
rect 11555 3232 11589 3266
rect 11589 3232 11657 3266
rect 11657 3232 11661 3266
rect 11483 3198 11661 3232
rect 11483 3194 11487 3198
rect 11487 3194 11555 3198
rect 11555 3194 11589 3198
rect 11589 3194 11657 3198
rect 11657 3194 11661 3198
rect 11555 3164 11589 3182
rect 11555 3148 11589 3164
rect 11483 3074 11517 3108
rect 11555 3074 11589 3108
rect 11627 3074 11661 3108
rect 11483 2994 11517 3028
rect 11555 2994 11589 3028
rect 11627 2994 11661 3028
rect 11483 2914 11517 2948
rect 11555 2914 11589 2948
rect 11627 2914 11661 2948
rect 11483 2834 11517 2868
rect 11555 2834 11589 2868
rect 11627 2834 11661 2868
rect 11483 2754 11517 2788
rect 11555 2754 11589 2788
rect 11627 2754 11661 2788
rect 11483 2674 11517 2708
rect 11555 2674 11589 2708
rect 11627 2674 11661 2708
rect 11483 2594 11517 2628
rect 11555 2594 11589 2628
rect 11627 2594 11661 2628
rect 11555 2540 11589 2556
rect 11555 2522 11589 2540
rect 11483 2506 11487 2518
rect 11487 2506 11555 2518
rect 11555 2506 11589 2518
rect 11589 2506 11657 2518
rect 11657 2506 11661 2518
rect 11483 2472 11661 2506
rect 11483 2438 11487 2472
rect 11487 2438 11555 2472
rect 11555 2438 11589 2472
rect 11589 2438 11657 2472
rect 11657 2438 11661 2472
rect 11483 2404 11661 2438
rect 11483 2370 11487 2404
rect 11487 2370 11555 2404
rect 11555 2370 11589 2404
rect 11589 2370 11657 2404
rect 11657 2370 11661 2404
rect 11483 2336 11661 2370
rect 11483 2302 11487 2336
rect 11487 2302 11555 2336
rect 11555 2302 11589 2336
rect 11589 2302 11657 2336
rect 11657 2302 11661 2336
rect 11483 2268 11661 2302
rect 11483 2234 11487 2268
rect 11487 2234 11555 2268
rect 11555 2234 11589 2268
rect 11589 2234 11657 2268
rect 11657 2234 11661 2268
rect 11483 2200 11661 2234
rect 11483 2166 11487 2200
rect 11487 2166 11555 2200
rect 11555 2166 11589 2200
rect 11589 2166 11657 2200
rect 11657 2166 11661 2200
rect 11483 2132 11661 2166
rect 11483 2098 11487 2132
rect 11487 2098 11555 2132
rect 11555 2098 11589 2132
rect 11589 2098 11657 2132
rect 11657 2098 11661 2132
rect 11483 2064 11661 2098
rect 11483 2030 11487 2064
rect 11487 2030 11555 2064
rect 11555 2030 11589 2064
rect 11589 2030 11657 2064
rect 11657 2030 11661 2064
rect 11483 1996 11661 2030
rect 11483 1962 11487 1996
rect 11487 1962 11555 1996
rect 11555 1962 11589 1996
rect 11589 1962 11657 1996
rect 11657 1962 11661 1996
rect 11483 1928 11661 1962
rect 11483 1894 11487 1928
rect 11487 1894 11555 1928
rect 11555 1894 11589 1928
rect 11589 1894 11657 1928
rect 11657 1894 11661 1928
rect 11483 1860 11661 1894
rect 11483 1826 11487 1860
rect 11487 1826 11555 1860
rect 11555 1826 11589 1860
rect 11589 1826 11657 1860
rect 11657 1826 11661 1860
rect 11483 1792 11661 1826
rect 11483 1758 11487 1792
rect 11487 1758 11555 1792
rect 11555 1758 11589 1792
rect 11589 1758 11657 1792
rect 11657 1758 11661 1792
rect 11483 1724 11661 1758
rect 11483 1690 11487 1724
rect 11487 1690 11555 1724
rect 11555 1690 11589 1724
rect 11589 1690 11657 1724
rect 11657 1690 11661 1724
rect 11483 1656 11661 1690
rect 11483 1622 11487 1656
rect 11487 1622 11555 1656
rect 11555 1622 11589 1656
rect 11589 1622 11657 1656
rect 11657 1622 11661 1656
rect 11483 1620 11661 1622
rect 11555 1586 11589 1620
rect 11238 1144 11344 1250
rect 11979 4064 12013 4098
rect 12051 4064 12085 4098
rect 12123 4064 12157 4098
rect 11979 3991 12013 4025
rect 12051 3991 12085 4025
rect 12123 3991 12157 4025
rect 11979 3918 12013 3952
rect 12051 3918 12085 3952
rect 12123 3918 12157 3952
rect 11979 3845 12013 3879
rect 12051 3845 12085 3879
rect 12123 3845 12157 3879
rect 11979 3772 12013 3806
rect 12051 3772 12085 3806
rect 12123 3772 12157 3806
rect 11979 3699 12013 3733
rect 12051 3699 12085 3733
rect 12123 3699 12157 3733
rect 11979 3626 12013 3660
rect 12051 3626 12085 3660
rect 12123 3626 12157 3660
rect 11979 3553 12013 3587
rect 12051 3553 12085 3587
rect 12123 3553 12157 3587
rect 11979 3480 12013 3514
rect 12051 3480 12085 3514
rect 12123 3480 12157 3514
rect 11979 3407 12013 3441
rect 12051 3407 12085 3441
rect 12123 3407 12157 3441
rect 11979 3334 12013 3368
rect 12051 3334 12085 3368
rect 12123 3334 12157 3368
rect 11979 3261 12013 3295
rect 12051 3261 12085 3295
rect 12123 3261 12157 3295
rect 11979 3188 12013 3222
rect 12051 3188 12085 3222
rect 12123 3188 12157 3222
rect 11979 3115 12013 3149
rect 12051 3115 12085 3149
rect 12123 3115 12157 3149
rect 11979 3042 12013 3076
rect 12051 3042 12085 3076
rect 12123 3042 12157 3076
rect 11979 2969 12013 3003
rect 12051 2969 12085 3003
rect 12123 2969 12157 3003
rect 11979 2896 12013 2930
rect 12051 2896 12085 2930
rect 12123 2896 12157 2930
rect 11979 2823 12013 2857
rect 12051 2823 12085 2857
rect 12123 2823 12157 2857
rect 11979 2750 12013 2784
rect 12051 2750 12085 2784
rect 12123 2750 12157 2784
rect 11979 2677 12013 2711
rect 12051 2677 12085 2711
rect 12123 2677 12157 2711
rect 11979 2604 12013 2638
rect 12051 2604 12085 2638
rect 12123 2604 12157 2638
rect 11979 2531 12013 2565
rect 12051 2531 12085 2565
rect 12123 2531 12157 2565
rect 11979 2458 12013 2492
rect 12051 2458 12085 2492
rect 12123 2458 12157 2492
rect 11979 2385 12013 2419
rect 12051 2385 12085 2419
rect 12123 2385 12157 2419
rect 11979 2312 12013 2346
rect 12051 2312 12085 2346
rect 12123 2312 12157 2346
rect 11979 2239 12013 2273
rect 12051 2239 12085 2273
rect 12123 2239 12157 2273
rect 11979 2166 12013 2200
rect 12051 2166 12085 2200
rect 12123 2166 12157 2200
rect 11979 2092 12013 2126
rect 12051 2092 12085 2126
rect 12123 2092 12157 2126
rect 11979 2018 12013 2052
rect 12051 2018 12085 2052
rect 12123 2018 12157 2052
rect 11979 1944 12013 1978
rect 12051 1944 12085 1978
rect 12123 1944 12157 1978
rect 11979 1870 12013 1904
rect 12051 1870 12085 1904
rect 12123 1870 12157 1904
rect 11979 1796 12013 1830
rect 12051 1796 12085 1830
rect 12123 1796 12157 1830
rect 11979 1722 12013 1756
rect 12051 1722 12085 1756
rect 12123 1722 12157 1756
rect 11979 1648 12013 1682
rect 12051 1648 12085 1682
rect 12123 1648 12157 1682
rect 11979 1574 12013 1608
rect 12051 1574 12085 1608
rect 12123 1574 12157 1608
rect 11800 1144 11906 1250
rect 12547 4092 12581 4118
rect 12475 4082 12653 4092
rect 12475 4048 12479 4082
rect 12479 4048 12547 4082
rect 12547 4048 12581 4082
rect 12581 4048 12649 4082
rect 12649 4048 12653 4082
rect 12475 4014 12653 4048
rect 12475 3980 12479 4014
rect 12479 3980 12547 4014
rect 12547 3980 12581 4014
rect 12581 3980 12649 4014
rect 12649 3980 12653 4014
rect 12475 3946 12653 3980
rect 12475 3912 12479 3946
rect 12479 3912 12547 3946
rect 12547 3912 12581 3946
rect 12581 3912 12649 3946
rect 12649 3912 12653 3946
rect 12475 3878 12653 3912
rect 12475 3844 12479 3878
rect 12479 3844 12547 3878
rect 12547 3844 12581 3878
rect 12581 3844 12649 3878
rect 12649 3844 12653 3878
rect 12475 3810 12653 3844
rect 12475 3776 12479 3810
rect 12479 3776 12547 3810
rect 12547 3776 12581 3810
rect 12581 3776 12649 3810
rect 12649 3776 12653 3810
rect 12475 3742 12653 3776
rect 12475 3708 12479 3742
rect 12479 3708 12547 3742
rect 12547 3708 12581 3742
rect 12581 3708 12649 3742
rect 12649 3708 12653 3742
rect 12475 3674 12653 3708
rect 12475 3640 12479 3674
rect 12479 3640 12547 3674
rect 12547 3640 12581 3674
rect 12581 3640 12649 3674
rect 12649 3640 12653 3674
rect 12475 3606 12653 3640
rect 12475 3572 12479 3606
rect 12479 3572 12547 3606
rect 12547 3572 12581 3606
rect 12581 3572 12649 3606
rect 12649 3572 12653 3606
rect 12475 3538 12653 3572
rect 12475 3504 12479 3538
rect 12479 3504 12547 3538
rect 12547 3504 12581 3538
rect 12581 3504 12649 3538
rect 12649 3504 12653 3538
rect 12475 3470 12653 3504
rect 12475 3436 12479 3470
rect 12479 3436 12547 3470
rect 12547 3436 12581 3470
rect 12581 3436 12649 3470
rect 12649 3436 12653 3470
rect 12475 3402 12653 3436
rect 12475 3368 12479 3402
rect 12479 3368 12547 3402
rect 12547 3368 12581 3402
rect 12581 3368 12649 3402
rect 12649 3368 12653 3402
rect 12475 3334 12653 3368
rect 12475 3300 12479 3334
rect 12479 3300 12547 3334
rect 12547 3300 12581 3334
rect 12581 3300 12649 3334
rect 12649 3300 12653 3334
rect 12475 3266 12653 3300
rect 12475 3232 12479 3266
rect 12479 3232 12547 3266
rect 12547 3232 12581 3266
rect 12581 3232 12649 3266
rect 12649 3232 12653 3266
rect 12475 3198 12653 3232
rect 12475 3194 12479 3198
rect 12479 3194 12547 3198
rect 12547 3194 12581 3198
rect 12581 3194 12649 3198
rect 12649 3194 12653 3198
rect 12547 3164 12581 3182
rect 12547 3148 12581 3164
rect 12475 3074 12509 3108
rect 12547 3074 12581 3108
rect 12619 3074 12653 3108
rect 12475 2994 12509 3028
rect 12547 2994 12581 3028
rect 12619 2994 12653 3028
rect 12475 2914 12509 2948
rect 12547 2914 12581 2948
rect 12619 2914 12653 2948
rect 12475 2834 12509 2868
rect 12547 2834 12581 2868
rect 12619 2834 12653 2868
rect 12475 2754 12509 2788
rect 12547 2754 12581 2788
rect 12619 2754 12653 2788
rect 12475 2674 12509 2708
rect 12547 2674 12581 2708
rect 12619 2674 12653 2708
rect 12475 2594 12509 2628
rect 12547 2594 12581 2628
rect 12619 2594 12653 2628
rect 12547 2540 12581 2556
rect 12547 2522 12581 2540
rect 12475 2506 12479 2518
rect 12479 2506 12547 2518
rect 12547 2506 12581 2518
rect 12581 2506 12649 2518
rect 12649 2506 12653 2518
rect 12475 2472 12653 2506
rect 12475 2438 12479 2472
rect 12479 2438 12547 2472
rect 12547 2438 12581 2472
rect 12581 2438 12649 2472
rect 12649 2438 12653 2472
rect 12475 2404 12653 2438
rect 12475 2370 12479 2404
rect 12479 2370 12547 2404
rect 12547 2370 12581 2404
rect 12581 2370 12649 2404
rect 12649 2370 12653 2404
rect 12475 2336 12653 2370
rect 12475 2302 12479 2336
rect 12479 2302 12547 2336
rect 12547 2302 12581 2336
rect 12581 2302 12649 2336
rect 12649 2302 12653 2336
rect 12475 2268 12653 2302
rect 12475 2234 12479 2268
rect 12479 2234 12547 2268
rect 12547 2234 12581 2268
rect 12581 2234 12649 2268
rect 12649 2234 12653 2268
rect 12475 2200 12653 2234
rect 12475 2166 12479 2200
rect 12479 2166 12547 2200
rect 12547 2166 12581 2200
rect 12581 2166 12649 2200
rect 12649 2166 12653 2200
rect 12475 2132 12653 2166
rect 12475 2098 12479 2132
rect 12479 2098 12547 2132
rect 12547 2098 12581 2132
rect 12581 2098 12649 2132
rect 12649 2098 12653 2132
rect 12475 2064 12653 2098
rect 12475 2030 12479 2064
rect 12479 2030 12547 2064
rect 12547 2030 12581 2064
rect 12581 2030 12649 2064
rect 12649 2030 12653 2064
rect 12475 1996 12653 2030
rect 12475 1962 12479 1996
rect 12479 1962 12547 1996
rect 12547 1962 12581 1996
rect 12581 1962 12649 1996
rect 12649 1962 12653 1996
rect 12475 1928 12653 1962
rect 12475 1894 12479 1928
rect 12479 1894 12547 1928
rect 12547 1894 12581 1928
rect 12581 1894 12649 1928
rect 12649 1894 12653 1928
rect 12475 1860 12653 1894
rect 12475 1826 12479 1860
rect 12479 1826 12547 1860
rect 12547 1826 12581 1860
rect 12581 1826 12649 1860
rect 12649 1826 12653 1860
rect 12475 1792 12653 1826
rect 12475 1758 12479 1792
rect 12479 1758 12547 1792
rect 12547 1758 12581 1792
rect 12581 1758 12649 1792
rect 12649 1758 12653 1792
rect 12475 1724 12653 1758
rect 12475 1690 12479 1724
rect 12479 1690 12547 1724
rect 12547 1690 12581 1724
rect 12581 1690 12649 1724
rect 12649 1690 12653 1724
rect 12475 1656 12653 1690
rect 12475 1622 12479 1656
rect 12479 1622 12547 1656
rect 12547 1622 12581 1656
rect 12581 1622 12649 1656
rect 12649 1622 12653 1656
rect 12475 1620 12653 1622
rect 12547 1586 12581 1620
rect 12230 1144 12336 1250
rect 12971 4064 13005 4098
rect 13043 4064 13077 4098
rect 13115 4064 13149 4098
rect 12971 3991 13005 4025
rect 13043 3991 13077 4025
rect 13115 3991 13149 4025
rect 12971 3918 13005 3952
rect 13043 3918 13077 3952
rect 13115 3918 13149 3952
rect 12971 3845 13005 3879
rect 13043 3845 13077 3879
rect 13115 3845 13149 3879
rect 12971 3772 13005 3806
rect 13043 3772 13077 3806
rect 13115 3772 13149 3806
rect 12971 3699 13005 3733
rect 13043 3699 13077 3733
rect 13115 3699 13149 3733
rect 12971 3626 13005 3660
rect 13043 3626 13077 3660
rect 13115 3626 13149 3660
rect 12971 3553 13005 3587
rect 13043 3553 13077 3587
rect 13115 3553 13149 3587
rect 12971 3480 13005 3514
rect 13043 3480 13077 3514
rect 13115 3480 13149 3514
rect 12971 3407 13005 3441
rect 13043 3407 13077 3441
rect 13115 3407 13149 3441
rect 12971 3334 13005 3368
rect 13043 3334 13077 3368
rect 13115 3334 13149 3368
rect 12971 3261 13005 3295
rect 13043 3261 13077 3295
rect 13115 3261 13149 3295
rect 12971 3188 13005 3222
rect 13043 3188 13077 3222
rect 13115 3188 13149 3222
rect 12971 3115 13005 3149
rect 13043 3115 13077 3149
rect 13115 3115 13149 3149
rect 12971 3042 13005 3076
rect 13043 3042 13077 3076
rect 13115 3042 13149 3076
rect 12971 2969 13005 3003
rect 13043 2969 13077 3003
rect 13115 2969 13149 3003
rect 12971 2896 13005 2930
rect 13043 2896 13077 2930
rect 13115 2896 13149 2930
rect 12971 2823 13005 2857
rect 13043 2823 13077 2857
rect 13115 2823 13149 2857
rect 12971 2750 13005 2784
rect 13043 2750 13077 2784
rect 13115 2750 13149 2784
rect 12971 2677 13005 2711
rect 13043 2677 13077 2711
rect 13115 2677 13149 2711
rect 12971 2604 13005 2638
rect 13043 2604 13077 2638
rect 13115 2604 13149 2638
rect 12971 2531 13005 2565
rect 13043 2531 13077 2565
rect 13115 2531 13149 2565
rect 12971 2458 13005 2492
rect 13043 2458 13077 2492
rect 13115 2458 13149 2492
rect 12971 2385 13005 2419
rect 13043 2385 13077 2419
rect 13115 2385 13149 2419
rect 12971 2312 13005 2346
rect 13043 2312 13077 2346
rect 13115 2312 13149 2346
rect 12971 2239 13005 2273
rect 13043 2239 13077 2273
rect 13115 2239 13149 2273
rect 12971 2166 13005 2200
rect 13043 2166 13077 2200
rect 13115 2166 13149 2200
rect 12971 2092 13005 2126
rect 13043 2092 13077 2126
rect 13115 2092 13149 2126
rect 12971 2018 13005 2052
rect 13043 2018 13077 2052
rect 13115 2018 13149 2052
rect 12971 1944 13005 1978
rect 13043 1944 13077 1978
rect 13115 1944 13149 1978
rect 12971 1870 13005 1904
rect 13043 1870 13077 1904
rect 13115 1870 13149 1904
rect 12971 1796 13005 1830
rect 13043 1796 13077 1830
rect 13115 1796 13149 1830
rect 12971 1722 13005 1756
rect 13043 1722 13077 1756
rect 13115 1722 13149 1756
rect 12971 1648 13005 1682
rect 13043 1648 13077 1682
rect 13115 1648 13149 1682
rect 12971 1574 13005 1608
rect 13043 1574 13077 1608
rect 13115 1574 13149 1608
rect 12792 1144 12898 1250
rect 13539 4092 13573 4118
rect 13467 4082 13645 4092
rect 13467 4048 13471 4082
rect 13471 4048 13539 4082
rect 13539 4048 13573 4082
rect 13573 4048 13641 4082
rect 13641 4048 13645 4082
rect 13467 4014 13645 4048
rect 13467 3980 13471 4014
rect 13471 3980 13539 4014
rect 13539 3980 13573 4014
rect 13573 3980 13641 4014
rect 13641 3980 13645 4014
rect 13467 3946 13645 3980
rect 13467 3912 13471 3946
rect 13471 3912 13539 3946
rect 13539 3912 13573 3946
rect 13573 3912 13641 3946
rect 13641 3912 13645 3946
rect 13467 3878 13645 3912
rect 13467 3844 13471 3878
rect 13471 3844 13539 3878
rect 13539 3844 13573 3878
rect 13573 3844 13641 3878
rect 13641 3844 13645 3878
rect 13467 3810 13645 3844
rect 13467 3776 13471 3810
rect 13471 3776 13539 3810
rect 13539 3776 13573 3810
rect 13573 3776 13641 3810
rect 13641 3776 13645 3810
rect 13467 3742 13645 3776
rect 13467 3708 13471 3742
rect 13471 3708 13539 3742
rect 13539 3708 13573 3742
rect 13573 3708 13641 3742
rect 13641 3708 13645 3742
rect 13467 3674 13645 3708
rect 13467 3640 13471 3674
rect 13471 3640 13539 3674
rect 13539 3640 13573 3674
rect 13573 3640 13641 3674
rect 13641 3640 13645 3674
rect 13467 3606 13645 3640
rect 13467 3572 13471 3606
rect 13471 3572 13539 3606
rect 13539 3572 13573 3606
rect 13573 3572 13641 3606
rect 13641 3572 13645 3606
rect 13467 3538 13645 3572
rect 13467 3504 13471 3538
rect 13471 3504 13539 3538
rect 13539 3504 13573 3538
rect 13573 3504 13641 3538
rect 13641 3504 13645 3538
rect 13467 3470 13645 3504
rect 13467 3436 13471 3470
rect 13471 3436 13539 3470
rect 13539 3436 13573 3470
rect 13573 3436 13641 3470
rect 13641 3436 13645 3470
rect 13467 3402 13645 3436
rect 13467 3368 13471 3402
rect 13471 3368 13539 3402
rect 13539 3368 13573 3402
rect 13573 3368 13641 3402
rect 13641 3368 13645 3402
rect 13467 3334 13645 3368
rect 13467 3300 13471 3334
rect 13471 3300 13539 3334
rect 13539 3300 13573 3334
rect 13573 3300 13641 3334
rect 13641 3300 13645 3334
rect 13467 3266 13645 3300
rect 13467 3232 13471 3266
rect 13471 3232 13539 3266
rect 13539 3232 13573 3266
rect 13573 3232 13641 3266
rect 13641 3232 13645 3266
rect 13467 3198 13645 3232
rect 13467 3194 13471 3198
rect 13471 3194 13539 3198
rect 13539 3194 13573 3198
rect 13573 3194 13641 3198
rect 13641 3194 13645 3198
rect 13539 3164 13573 3182
rect 13539 3148 13573 3164
rect 13467 3074 13501 3108
rect 13539 3074 13573 3108
rect 13611 3074 13645 3108
rect 13467 2994 13501 3028
rect 13539 2994 13573 3028
rect 13611 2994 13645 3028
rect 13467 2914 13501 2948
rect 13539 2914 13573 2948
rect 13611 2914 13645 2948
rect 13467 2834 13501 2868
rect 13539 2834 13573 2868
rect 13611 2834 13645 2868
rect 13467 2754 13501 2788
rect 13539 2754 13573 2788
rect 13611 2754 13645 2788
rect 13467 2674 13501 2708
rect 13539 2674 13573 2708
rect 13611 2674 13645 2708
rect 13467 2594 13501 2628
rect 13539 2594 13573 2628
rect 13611 2594 13645 2628
rect 13539 2540 13573 2556
rect 13539 2522 13573 2540
rect 13467 2506 13471 2518
rect 13471 2506 13539 2518
rect 13539 2506 13573 2518
rect 13573 2506 13641 2518
rect 13641 2506 13645 2518
rect 13467 2472 13645 2506
rect 13467 2438 13471 2472
rect 13471 2438 13539 2472
rect 13539 2438 13573 2472
rect 13573 2438 13641 2472
rect 13641 2438 13645 2472
rect 13467 2404 13645 2438
rect 13467 2370 13471 2404
rect 13471 2370 13539 2404
rect 13539 2370 13573 2404
rect 13573 2370 13641 2404
rect 13641 2370 13645 2404
rect 13467 2336 13645 2370
rect 13467 2302 13471 2336
rect 13471 2302 13539 2336
rect 13539 2302 13573 2336
rect 13573 2302 13641 2336
rect 13641 2302 13645 2336
rect 13467 2268 13645 2302
rect 13467 2234 13471 2268
rect 13471 2234 13539 2268
rect 13539 2234 13573 2268
rect 13573 2234 13641 2268
rect 13641 2234 13645 2268
rect 13467 2200 13645 2234
rect 13467 2166 13471 2200
rect 13471 2166 13539 2200
rect 13539 2166 13573 2200
rect 13573 2166 13641 2200
rect 13641 2166 13645 2200
rect 13467 2132 13645 2166
rect 13467 2098 13471 2132
rect 13471 2098 13539 2132
rect 13539 2098 13573 2132
rect 13573 2098 13641 2132
rect 13641 2098 13645 2132
rect 13467 2064 13645 2098
rect 13467 2030 13471 2064
rect 13471 2030 13539 2064
rect 13539 2030 13573 2064
rect 13573 2030 13641 2064
rect 13641 2030 13645 2064
rect 13467 1996 13645 2030
rect 13467 1962 13471 1996
rect 13471 1962 13539 1996
rect 13539 1962 13573 1996
rect 13573 1962 13641 1996
rect 13641 1962 13645 1996
rect 13467 1928 13645 1962
rect 13467 1894 13471 1928
rect 13471 1894 13539 1928
rect 13539 1894 13573 1928
rect 13573 1894 13641 1928
rect 13641 1894 13645 1928
rect 13467 1860 13645 1894
rect 13467 1826 13471 1860
rect 13471 1826 13539 1860
rect 13539 1826 13573 1860
rect 13573 1826 13641 1860
rect 13641 1826 13645 1860
rect 13467 1792 13645 1826
rect 13467 1758 13471 1792
rect 13471 1758 13539 1792
rect 13539 1758 13573 1792
rect 13573 1758 13641 1792
rect 13641 1758 13645 1792
rect 13467 1724 13645 1758
rect 13467 1690 13471 1724
rect 13471 1690 13539 1724
rect 13539 1690 13573 1724
rect 13573 1690 13641 1724
rect 13641 1690 13645 1724
rect 13467 1656 13645 1690
rect 13467 1622 13471 1656
rect 13471 1622 13539 1656
rect 13539 1622 13573 1656
rect 13573 1622 13641 1656
rect 13641 1622 13645 1656
rect 13467 1620 13645 1622
rect 13539 1586 13573 1620
rect 13222 1144 13328 1250
rect 13963 4064 13997 4098
rect 14035 4064 14069 4098
rect 13963 3990 13997 4024
rect 14035 3990 14069 4024
rect 13963 3916 13997 3950
rect 14035 3916 14069 3950
rect 13963 3842 13997 3876
rect 14035 3842 14069 3876
rect 13963 3768 13997 3802
rect 14035 3768 14069 3802
rect 13963 3694 13997 3728
rect 14035 3694 14069 3728
rect 13963 3620 13997 3654
rect 14035 3620 14069 3654
rect 13963 3546 13997 3580
rect 14035 3546 14069 3580
rect 13963 3472 13997 3506
rect 14035 3472 14069 3506
rect 13963 3398 13997 3432
rect 14035 3398 14069 3432
rect 13963 3324 13997 3358
rect 14035 3324 14069 3358
rect 13963 3250 13997 3284
rect 14035 3250 14069 3284
rect 13963 3176 13997 3210
rect 14035 3176 14069 3210
rect 13963 3102 13997 3136
rect 14035 3102 14069 3136
rect 13963 3028 13997 3062
rect 14035 3028 14069 3062
rect 13963 2954 13997 2988
rect 14035 2954 14069 2988
rect 13963 2880 13997 2914
rect 14035 2880 14069 2914
rect 13963 2806 13997 2840
rect 14035 2806 14069 2840
rect 13963 2732 13997 2766
rect 14035 2732 14069 2766
rect 13963 2658 13997 2692
rect 14035 2658 14069 2692
rect 13963 2584 13997 2618
rect 14035 2584 14069 2618
rect 13963 2510 13997 2544
rect 14035 2510 14069 2544
rect 13963 2436 13997 2470
rect 14035 2436 14069 2470
rect 13963 2362 13997 2396
rect 14035 2362 14069 2396
rect 13963 2288 13997 2322
rect 14035 2288 14069 2322
rect 13963 2214 13997 2248
rect 14035 2214 14069 2248
rect 13963 2140 13997 2174
rect 14035 2140 14069 2174
rect 13963 2066 13997 2100
rect 14035 2066 14069 2100
rect 13963 1992 13997 2026
rect 14035 1992 14069 2026
rect 13963 1918 13997 1952
rect 14035 1918 14069 1952
rect 13963 1844 13997 1878
rect 14035 1844 14069 1878
rect 13963 1770 13997 1804
rect 14035 1770 14069 1804
rect 13963 1696 13997 1730
rect 14035 1696 14069 1730
rect 13963 1622 13997 1656
rect 14035 1622 14069 1656
rect 13963 1548 13997 1582
rect 14035 1548 14069 1582
rect 13784 1144 13890 1250
rect 14142 1144 14248 1250
rect 14356 4252 14390 4286
rect 14356 4179 14390 4213
rect 14356 4106 14390 4140
rect 14356 4048 14390 4067
rect 14356 4033 14390 4048
rect 14356 3980 14390 3994
rect 14356 3960 14390 3980
rect 14428 3992 14468 4426
rect 14468 3992 14606 4426
rect 14428 3960 14536 3992
rect 14536 3960 14606 3992
rect 14356 3912 14390 3921
rect 14428 3918 14462 3952
rect 14356 3887 14390 3912
rect 14500 3888 14534 3921
rect 14572 3905 14604 3921
rect 14604 3905 14606 3921
rect 14500 3887 14502 3888
rect 14502 3887 14534 3888
rect 14356 3844 14390 3848
rect 14428 3846 14462 3880
rect 14572 3887 14606 3905
rect 14356 3814 14390 3844
rect 14500 3819 14534 3848
rect 14572 3837 14604 3848
rect 14604 3837 14606 3848
rect 14500 3814 14502 3819
rect 14502 3814 14534 3819
rect 14356 3742 14390 3775
rect 14428 3774 14462 3808
rect 14572 3814 14606 3837
rect 14500 3750 14534 3775
rect 14572 3769 14604 3775
rect 14604 3769 14606 3775
rect 14356 3741 14390 3742
rect 14500 3741 14502 3750
rect 14502 3741 14534 3750
rect 14428 3702 14462 3736
rect 14572 3741 14606 3769
rect 14356 3674 14390 3702
rect 14500 3681 14534 3702
rect 14572 3701 14604 3702
rect 14604 3701 14606 3702
rect 14356 3668 14390 3674
rect 14500 3668 14502 3681
rect 14502 3668 14534 3681
rect 14428 3630 14462 3664
rect 14572 3668 14606 3701
rect 14356 3606 14390 3629
rect 14500 3612 14534 3629
rect 14356 3595 14390 3606
rect 14500 3595 14502 3612
rect 14502 3595 14534 3612
rect 14428 3558 14462 3592
rect 14572 3599 14606 3629
rect 14572 3595 14604 3599
rect 14604 3595 14606 3599
rect 14356 3538 14390 3556
rect 14500 3543 14534 3556
rect 14356 3522 14390 3538
rect 14500 3522 14502 3543
rect 14502 3522 14534 3543
rect 14428 3486 14462 3520
rect 14572 3531 14606 3556
rect 14572 3522 14604 3531
rect 14604 3522 14606 3531
rect 14356 3470 14390 3483
rect 14500 3474 14534 3483
rect 14356 3449 14390 3470
rect 14500 3449 14502 3474
rect 14502 3449 14534 3474
rect 14428 3414 14462 3448
rect 14572 3463 14606 3483
rect 14572 3449 14604 3463
rect 14604 3449 14606 3463
rect 14356 3402 14390 3410
rect 14500 3405 14534 3410
rect 14356 3376 14390 3402
rect 14500 3376 14502 3405
rect 14502 3376 14534 3405
rect 14428 3342 14462 3376
rect 14572 3395 14606 3410
rect 14572 3376 14604 3395
rect 14604 3376 14606 3395
rect 14356 3334 14390 3337
rect 14500 3336 14534 3337
rect 14356 3303 14390 3334
rect 14428 3270 14462 3304
rect 14500 3303 14502 3336
rect 14502 3303 14534 3336
rect 14572 3327 14606 3337
rect 14572 3303 14604 3327
rect 14604 3303 14606 3327
rect 14356 3232 14390 3264
rect 14500 3233 14502 3264
rect 14502 3233 14534 3264
rect 14572 3259 14606 3264
rect 14356 3230 14390 3232
rect 14428 3198 14462 3232
rect 14500 3230 14534 3233
rect 14572 3230 14604 3259
rect 14604 3230 14606 3259
rect 14356 3164 14390 3191
rect 14500 3164 14502 3191
rect 14502 3164 14534 3191
rect 14356 3157 14390 3164
rect 14428 3126 14462 3160
rect 14500 3157 14534 3164
rect 14572 3157 14604 3191
rect 14604 3157 14606 3191
rect 14356 3084 14390 3118
rect 14500 3095 14502 3118
rect 14502 3095 14534 3118
rect 14428 3054 14462 3088
rect 14500 3084 14534 3095
rect 14572 3089 14604 3118
rect 14604 3089 14606 3118
rect 14572 3084 14606 3089
rect 14356 3011 14390 3045
rect 14500 3026 14502 3045
rect 14502 3026 14534 3045
rect 14428 2982 14462 3016
rect 14500 3011 14534 3026
rect 14572 3021 14604 3045
rect 14604 3021 14606 3045
rect 14572 3011 14606 3021
rect 14356 2938 14390 2972
rect 14500 2957 14502 2972
rect 14502 2957 14534 2972
rect 14428 2910 14462 2944
rect 14500 2938 14534 2957
rect 14572 2953 14604 2972
rect 14604 2953 14606 2972
rect 14572 2938 14606 2953
rect 14356 2865 14390 2899
rect 14500 2888 14502 2899
rect 14502 2888 14534 2899
rect 14428 2838 14462 2872
rect 14500 2865 14534 2888
rect 14572 2885 14604 2899
rect 14604 2885 14606 2899
rect 14572 2865 14606 2885
rect 14356 2792 14390 2826
rect 14500 2819 14502 2826
rect 14502 2819 14534 2826
rect 14428 2766 14462 2800
rect 14500 2792 14534 2819
rect 14572 2817 14604 2826
rect 14604 2817 14606 2826
rect 14572 2792 14606 2817
rect 14356 2719 14390 2753
rect 14500 2750 14502 2753
rect 14502 2750 14534 2753
rect 14428 2694 14462 2728
rect 14500 2719 14534 2750
rect 14572 2749 14604 2753
rect 14604 2749 14606 2753
rect 14572 2719 14606 2749
rect 14356 2646 14390 2680
rect 14428 2622 14462 2656
rect 14500 2646 14534 2680
rect 14572 2647 14606 2680
rect 14572 2646 14604 2647
rect 14604 2646 14606 2647
rect 14356 2573 14390 2607
rect 14428 2550 14462 2584
rect 14500 2577 14534 2607
rect 14572 2579 14606 2607
rect 14500 2573 14502 2577
rect 14502 2573 14534 2577
rect 14572 2573 14604 2579
rect 14604 2573 14606 2579
rect 14356 2500 14390 2534
rect 14428 2478 14462 2512
rect 14500 2508 14534 2534
rect 14572 2511 14606 2534
rect 14500 2500 14502 2508
rect 14502 2500 14534 2508
rect 14572 2500 14604 2511
rect 14604 2500 14606 2511
rect 14356 2448 14390 2461
rect 14356 2427 14390 2448
rect 14428 2406 14462 2440
rect 14500 2439 14534 2461
rect 14572 2443 14606 2461
rect 14500 2427 14502 2439
rect 14502 2427 14534 2439
rect 14572 2427 14604 2443
rect 14604 2427 14606 2443
rect 14356 2380 14390 2388
rect 14356 2354 14390 2380
rect 14500 2370 14534 2388
rect 14572 2375 14606 2388
rect 14428 2334 14462 2368
rect 14500 2354 14502 2370
rect 14502 2354 14534 2370
rect 14572 2354 14604 2375
rect 14604 2354 14606 2375
rect 14356 2312 14390 2315
rect 14356 2281 14390 2312
rect 14500 2301 14534 2315
rect 14572 2307 14606 2315
rect 14428 2262 14462 2296
rect 14500 2281 14502 2301
rect 14502 2281 14534 2301
rect 14572 2281 14604 2307
rect 14604 2281 14606 2307
rect 14356 2210 14390 2242
rect 14500 2232 14534 2242
rect 14572 2239 14606 2242
rect 14356 2208 14390 2210
rect 14428 2190 14462 2224
rect 14500 2208 14502 2232
rect 14502 2208 14534 2232
rect 14572 2208 14604 2239
rect 14604 2208 14606 2239
rect 14356 2142 14390 2169
rect 14500 2163 14534 2169
rect 14356 2135 14390 2142
rect 14428 2118 14462 2152
rect 14500 2135 14502 2163
rect 14502 2135 14534 2163
rect 14572 2137 14604 2169
rect 14604 2137 14606 2169
rect 14572 2135 14606 2137
rect 14356 2074 14390 2096
rect 14500 2094 14534 2096
rect 14356 2062 14390 2074
rect 14428 2046 14462 2080
rect 14500 2062 14502 2094
rect 14502 2062 14534 2094
rect 14572 2069 14604 2096
rect 14604 2069 14606 2096
rect 14572 2062 14606 2069
rect 14356 2006 14390 2023
rect 14356 1989 14390 2006
rect 14428 1974 14462 2008
rect 14500 1991 14502 2023
rect 14502 1991 14534 2023
rect 14572 2001 14604 2023
rect 14604 2001 14606 2023
rect 14500 1989 14534 1991
rect 14572 1989 14606 2001
rect 14356 1938 14390 1950
rect 14356 1916 14390 1938
rect 14428 1902 14462 1936
rect 14500 1922 14502 1950
rect 14502 1922 14534 1950
rect 14572 1933 14604 1950
rect 14604 1933 14606 1950
rect 14500 1916 14534 1922
rect 14572 1916 14606 1933
rect 14356 1870 14390 1877
rect 14356 1843 14390 1870
rect 14428 1830 14462 1864
rect 14500 1853 14502 1877
rect 14502 1853 14534 1877
rect 14572 1865 14604 1877
rect 14604 1865 14606 1877
rect 14500 1843 14534 1853
rect 14572 1843 14606 1865
rect 14356 1802 14390 1804
rect 14356 1770 14390 1802
rect 14428 1758 14462 1792
rect 14500 1784 14502 1804
rect 14502 1784 14534 1804
rect 14572 1797 14604 1804
rect 14604 1797 14606 1804
rect 14500 1770 14534 1784
rect 14572 1770 14606 1797
rect 14356 1700 14390 1731
rect 14356 1697 14390 1700
rect 14428 1686 14462 1720
rect 14500 1715 14502 1731
rect 14502 1715 14534 1731
rect 14572 1729 14604 1731
rect 14604 1729 14606 1731
rect 14500 1697 14534 1715
rect 14572 1697 14606 1729
rect 14356 1632 14390 1657
rect 14356 1623 14390 1632
rect 14428 1614 14462 1648
rect 14500 1646 14502 1658
rect 14502 1646 14534 1658
rect 14500 1624 14534 1646
rect 14572 1627 14606 1658
rect 14572 1624 14604 1627
rect 14604 1624 14606 1627
rect 14356 1564 14390 1583
rect 14500 1577 14502 1585
rect 14502 1577 14534 1585
rect 14356 1549 14390 1564
rect 14428 1542 14462 1576
rect 14500 1551 14534 1577
rect 14572 1559 14606 1585
rect 14572 1551 14604 1559
rect 14604 1551 14606 1559
rect 14356 1475 14390 1509
rect 14500 1508 14502 1512
rect 14502 1508 14534 1512
rect 14428 1470 14462 1504
rect 14500 1478 14534 1508
rect 14572 1491 14606 1512
rect 14572 1478 14604 1491
rect 14604 1478 14606 1491
rect 14356 1401 14390 1435
rect 14428 1398 14462 1432
rect 14500 1405 14534 1439
rect 14572 1423 14606 1439
rect 14572 1405 14604 1423
rect 14604 1405 14606 1423
rect 14356 1327 14390 1361
rect 14428 1326 14462 1360
rect 14500 1335 14534 1366
rect 14572 1355 14606 1366
rect 14500 1332 14502 1335
rect 14502 1332 14534 1335
rect 14572 1332 14604 1355
rect 14604 1332 14606 1355
rect 14356 1253 14390 1287
rect 14428 1254 14462 1288
rect 14500 1266 14534 1293
rect 14572 1287 14606 1293
rect 14500 1259 14502 1266
rect 14502 1259 14534 1266
rect 14572 1259 14604 1287
rect 14604 1259 14606 1287
rect 14356 1179 14390 1213
rect 14428 1182 14462 1216
rect 14500 1197 14534 1220
rect 14572 1218 14606 1220
rect 14500 1186 14502 1197
rect 14502 1186 14534 1197
rect 14572 1186 14604 1218
rect 14604 1186 14606 1218
rect 746 883 780 894
rect 14356 1105 14390 1139
rect 14428 1110 14462 1144
rect 14500 1128 14534 1147
rect 14500 1113 14502 1128
rect 14502 1113 14534 1128
rect 14572 1115 14604 1147
rect 14604 1115 14606 1147
rect 14572 1113 14606 1115
rect 14356 1031 14390 1065
rect 14428 1038 14462 1072
rect 14500 1059 14534 1074
rect 14500 1040 14502 1059
rect 14502 1040 14534 1059
rect 14572 1046 14604 1074
rect 14604 1046 14606 1074
rect 14572 1040 14606 1046
rect 14356 957 14390 991
rect 14428 966 14462 1000
rect 14500 990 14534 1001
rect 14500 967 14502 990
rect 14502 967 14534 990
rect 14572 977 14604 1001
rect 14604 977 14606 1001
rect 14572 967 14606 977
rect 14356 883 14390 917
rect 14428 894 14462 928
rect 14500 921 14534 928
rect 14500 894 14502 921
rect 14502 894 14534 921
rect 14572 908 14604 928
rect 14604 908 14606 928
rect 14572 894 14606 908
rect 709 818 736 820
rect 736 818 743 820
rect 782 818 805 820
rect 805 818 816 820
rect 855 818 874 820
rect 874 818 889 820
rect 928 818 943 820
rect 943 818 978 820
rect 978 818 1012 820
rect 1012 818 1047 820
rect 1047 818 1081 820
rect 1081 818 1116 820
rect 1116 818 1150 820
rect 1150 818 1185 820
rect 1185 818 1219 820
rect 1219 818 1254 820
rect 1254 818 1288 820
rect 1288 818 1323 820
rect 1323 818 1357 820
rect 1357 818 1392 820
rect 1392 818 1426 820
rect 1426 818 1461 820
rect 1461 818 1495 820
rect 1495 818 1530 820
rect 1530 818 1564 820
rect 1564 818 1599 820
rect 1599 818 1633 820
rect 1633 818 1668 820
rect 1668 818 1702 820
rect 1702 818 1737 820
rect 1737 818 1771 820
rect 1771 818 1806 820
rect 1806 818 1840 820
rect 1840 818 1875 820
rect 1875 818 1909 820
rect 1909 818 1944 820
rect 1944 818 1978 820
rect 1978 818 2013 820
rect 2013 818 2047 820
rect 2047 818 2082 820
rect 2082 818 2116 820
rect 2116 818 2151 820
rect 2151 818 2185 820
rect 2185 818 2220 820
rect 2220 818 2254 820
rect 2254 818 2289 820
rect 2289 818 2323 820
rect 2323 818 2358 820
rect 2358 818 2392 820
rect 2392 818 2427 820
rect 2427 818 2461 820
rect 2461 818 2496 820
rect 2496 818 2530 820
rect 2530 818 2565 820
rect 2565 818 2599 820
rect 2599 818 2634 820
rect 2634 818 2668 820
rect 2668 818 2703 820
rect 2703 818 2737 820
rect 2737 818 2772 820
rect 709 786 743 818
rect 782 786 816 818
rect 855 786 889 818
rect 928 784 2772 818
rect 928 750 944 784
rect 944 750 979 784
rect 979 750 1013 784
rect 1013 750 1048 784
rect 1048 750 1082 784
rect 1082 750 1117 784
rect 1117 750 1151 784
rect 1151 750 1186 784
rect 1186 750 1220 784
rect 1220 750 1255 784
rect 1255 750 1289 784
rect 1289 750 1324 784
rect 1324 750 1358 784
rect 1358 750 1393 784
rect 1393 750 1427 784
rect 1427 750 1462 784
rect 1462 750 1496 784
rect 1496 750 1531 784
rect 1531 750 1565 784
rect 1565 750 1600 784
rect 1600 750 1634 784
rect 1634 750 1669 784
rect 1669 750 1703 784
rect 1703 750 1738 784
rect 1738 750 1772 784
rect 1772 750 1807 784
rect 1807 750 1841 784
rect 1841 750 1876 784
rect 1876 750 1910 784
rect 1910 750 1945 784
rect 1945 750 1979 784
rect 1979 750 2014 784
rect 2014 750 2048 784
rect 2048 750 2083 784
rect 2083 750 2117 784
rect 2117 750 2152 784
rect 2152 750 2186 784
rect 2186 750 2221 784
rect 2221 750 2255 784
rect 2255 750 2290 784
rect 2290 750 2324 784
rect 2324 750 2359 784
rect 2359 750 2393 784
rect 2393 750 2428 784
rect 2428 750 2462 784
rect 2462 750 2497 784
rect 2497 750 2531 784
rect 2531 750 2566 784
rect 2566 750 2600 784
rect 2600 750 2635 784
rect 2635 750 2669 784
rect 2669 750 2704 784
rect 2704 750 2738 784
rect 2738 750 2772 784
rect 2772 750 14426 820
rect 709 716 743 748
rect 782 716 816 748
rect 855 716 889 748
rect 928 716 4725 750
rect 709 714 723 716
rect 723 714 743 716
rect 782 714 792 716
rect 792 714 816 716
rect 855 714 861 716
rect 861 714 889 716
rect 928 714 930 716
rect 930 714 964 716
rect 964 714 999 716
rect 999 714 1033 716
rect 1033 714 1068 716
rect 1068 714 1102 716
rect 1102 714 1137 716
rect 1137 714 1171 716
rect 1171 714 1206 716
rect 1206 714 1240 716
rect 1240 714 1275 716
rect 1275 714 1309 716
rect 1309 714 1344 716
rect 1344 714 1378 716
rect 1378 714 1413 716
rect 1413 714 1447 716
rect 1447 714 1482 716
rect 1482 714 1516 716
rect 1516 714 1551 716
rect 1551 714 1585 716
rect 1585 714 1620 716
rect 1620 714 1654 716
rect 1654 714 1689 716
rect 1689 714 1723 716
rect 1723 714 1758 716
rect 1758 714 1792 716
rect 1792 714 1827 716
rect 1827 714 1861 716
rect 1861 714 1896 716
rect 1896 714 1930 716
rect 1930 714 1965 716
rect 1965 714 1999 716
rect 1999 714 2034 716
rect 2034 714 2068 716
rect 2068 714 2103 716
rect 2103 714 2137 716
rect 2137 714 2172 716
rect 2172 714 2206 716
rect 2206 714 2241 716
rect 2241 714 2275 716
rect 2275 714 2310 716
rect 2310 714 2344 716
rect 2344 714 2379 716
rect 2379 714 2413 716
rect 2413 714 2448 716
rect 2448 714 2482 716
rect 2482 714 2517 716
rect 2517 714 2551 716
rect 2551 714 2586 716
rect 2586 714 2620 716
rect 2620 714 2655 716
rect 2655 714 2689 716
rect 2689 714 2724 716
rect 2724 714 2758 716
rect 2758 714 2793 716
rect 2793 714 2827 716
rect 2827 714 2862 716
rect 2862 714 2896 716
rect 2896 714 2931 716
rect 2931 714 2965 716
rect 2965 714 3000 716
rect 3000 714 3034 716
rect 3034 714 3069 716
rect 3069 714 3103 716
rect 3103 714 3138 716
rect 3138 714 3172 716
rect 3172 714 3207 716
rect 3207 714 3241 716
rect 3241 714 3276 716
rect 3276 714 3310 716
rect 3310 714 3345 716
rect 3345 714 3379 716
rect 3379 714 3414 716
rect 3414 714 3448 716
rect 3448 714 3483 716
rect 3483 714 3517 716
rect 3517 714 3552 716
rect 3552 714 3586 716
rect 3586 714 3621 716
rect 3621 714 3655 716
rect 3655 714 3690 716
rect 3690 714 3724 716
rect 3724 714 3759 716
rect 3759 714 3793 716
rect 3793 714 3828 716
rect 3828 714 3862 716
rect 3862 714 3897 716
rect 3897 714 3931 716
rect 3931 714 3966 716
rect 3966 714 4000 716
rect 4000 714 4035 716
rect 4035 714 4069 716
rect 4069 714 4104 716
rect 4104 714 4138 716
rect 4138 714 4173 716
rect 4173 714 4207 716
rect 4207 714 4242 716
rect 4242 714 4276 716
rect 4276 714 4311 716
rect 4311 714 4345 716
rect 4345 714 4380 716
rect 4380 714 4414 716
rect 4414 714 4449 716
rect 4449 714 4483 716
rect 4483 714 4518 716
rect 4518 714 4552 716
rect 4552 714 4587 716
rect 4587 714 4621 716
rect 4621 714 4656 716
rect 4656 714 4690 716
rect 4690 714 4725 716
rect 4725 714 14426 750
rect 14835 4645 15013 4679
rect 14835 4611 14840 4645
rect 14840 4611 14906 4645
rect 14906 4611 14940 4645
rect 14940 4611 15013 4645
rect 14835 4577 15013 4611
rect 14835 4543 14840 4577
rect 14840 4543 14906 4577
rect 14906 4543 14940 4577
rect 14940 4543 15013 4577
rect 14835 4509 15013 4543
rect 14835 4475 14840 4509
rect 14840 4475 14906 4509
rect 14906 4475 14940 4509
rect 14940 4475 15013 4509
rect 14835 4441 15013 4475
rect 14835 4407 14840 4441
rect 14840 4407 14906 4441
rect 14906 4407 14940 4441
rect 14940 4407 15013 4441
rect 14835 4373 15013 4407
rect 14835 4339 14840 4373
rect 14840 4339 14906 4373
rect 14906 4339 14940 4373
rect 14940 4339 15013 4373
rect 14835 4305 15013 4339
rect 14835 4271 14840 4305
rect 14840 4271 14906 4305
rect 14906 4271 14940 4305
rect 14940 4271 15013 4305
rect 14835 4237 15013 4271
rect 14835 4203 14840 4237
rect 14840 4203 14906 4237
rect 14906 4203 14940 4237
rect 14940 4203 15013 4237
rect 14835 4169 15013 4203
rect 14835 4135 14840 4169
rect 14840 4135 14906 4169
rect 14906 4135 14940 4169
rect 14940 4135 15013 4169
rect 14835 4101 15013 4135
rect 14835 4067 14840 4101
rect 14840 4067 14906 4101
rect 14906 4067 14940 4101
rect 14940 4067 15013 4101
rect 14835 4033 15013 4067
rect 14835 3999 14840 4033
rect 14840 3999 14906 4033
rect 14906 3999 14940 4033
rect 14940 3999 15013 4033
rect 14835 3965 15013 3999
rect 14835 3931 14840 3965
rect 14840 3931 14906 3965
rect 14906 3931 14940 3965
rect 14940 3931 15013 3965
rect 14835 3897 15013 3931
rect 14835 3863 14840 3897
rect 14840 3863 14906 3897
rect 14906 3863 14940 3897
rect 14940 3863 15013 3897
rect 14835 3829 15013 3863
rect 14835 3795 14840 3829
rect 14840 3795 14906 3829
rect 14906 3795 14940 3829
rect 14940 3795 15013 3829
rect 14835 3761 15013 3795
rect 14835 3727 14840 3761
rect 14840 3727 14906 3761
rect 14906 3727 14940 3761
rect 14940 3727 15013 3761
rect 14835 3693 15013 3727
rect 14835 3659 14840 3693
rect 14840 3659 14906 3693
rect 14906 3659 14940 3693
rect 14940 3659 15013 3693
rect 14835 3625 15013 3659
rect 14835 3591 14840 3625
rect 14840 3591 14906 3625
rect 14906 3591 14940 3625
rect 14940 3591 15013 3625
rect 14835 3557 15013 3591
rect 14835 3523 14840 3557
rect 14840 3523 14906 3557
rect 14906 3523 14940 3557
rect 14940 3523 15013 3557
rect 14835 3489 15013 3523
rect 14835 3455 14840 3489
rect 14840 3455 14906 3489
rect 14906 3455 14940 3489
rect 14940 3455 15013 3489
rect 14835 3421 15013 3455
rect 14835 3387 14840 3421
rect 14840 3387 14906 3421
rect 14906 3387 14940 3421
rect 14940 3387 15013 3421
rect 14835 3353 15013 3387
rect 14835 3319 14840 3353
rect 14840 3319 14906 3353
rect 14906 3319 14940 3353
rect 14940 3319 15013 3353
rect 14835 3285 15013 3319
rect 14835 3251 14840 3285
rect 14840 3251 14906 3285
rect 14906 3251 14940 3285
rect 14940 3251 15013 3285
rect 14835 3217 15013 3251
rect 14835 3183 14840 3217
rect 14840 3183 14906 3217
rect 14906 3183 14940 3217
rect 14940 3183 15013 3217
rect 14835 3149 15013 3183
rect 14835 3115 14840 3149
rect 14840 3115 14906 3149
rect 14906 3115 14940 3149
rect 14940 3115 15013 3149
rect 14835 3081 15013 3115
rect 14835 3047 14840 3081
rect 14840 3047 14906 3081
rect 14906 3047 14940 3081
rect 14940 3047 15013 3081
rect 14835 3013 15013 3047
rect 14835 2979 14840 3013
rect 14840 2979 14906 3013
rect 14906 2979 14940 3013
rect 14940 2979 15013 3013
rect 14835 2945 15013 2979
rect 14835 2911 14840 2945
rect 14840 2911 14906 2945
rect 14906 2911 14940 2945
rect 14940 2911 15013 2945
rect 14835 2877 15013 2911
rect 14835 2843 14840 2877
rect 14840 2843 14906 2877
rect 14906 2843 14940 2877
rect 14940 2843 15013 2877
rect 14835 2809 15013 2843
rect 14835 2775 14840 2809
rect 14840 2775 14906 2809
rect 14906 2775 14940 2809
rect 14940 2775 15013 2809
rect 14835 2741 15013 2775
rect 14835 2707 14840 2741
rect 14840 2707 14906 2741
rect 14906 2707 14940 2741
rect 14940 2707 15013 2741
rect 14835 2673 15013 2707
rect 14835 2639 14840 2673
rect 14840 2639 14906 2673
rect 14906 2639 14940 2673
rect 14940 2639 15013 2673
rect 14835 2605 15013 2639
rect 14835 2571 14840 2605
rect 14840 2571 14906 2605
rect 14906 2571 14940 2605
rect 14940 2571 15013 2605
rect 14835 2537 15013 2571
rect 14835 2503 14840 2537
rect 14840 2503 14906 2537
rect 14906 2503 14940 2537
rect 14940 2503 15013 2537
rect 14835 2469 15013 2503
rect 14835 2435 14840 2469
rect 14840 2435 14906 2469
rect 14906 2435 14940 2469
rect 14940 2435 15013 2469
rect 14835 2401 15013 2435
rect 14835 2367 14840 2401
rect 14840 2367 14906 2401
rect 14906 2367 14940 2401
rect 14940 2367 15013 2401
rect 14835 2333 15013 2367
rect 14835 2299 14840 2333
rect 14840 2299 14906 2333
rect 14906 2299 14940 2333
rect 14940 2299 15013 2333
rect 14835 2265 15013 2299
rect 14835 2231 14840 2265
rect 14840 2231 14906 2265
rect 14906 2231 14940 2265
rect 14940 2231 15013 2265
rect 14835 2197 15013 2231
rect 14835 2163 14840 2197
rect 14840 2163 14906 2197
rect 14906 2163 14940 2197
rect 14940 2163 15013 2197
rect 14835 2129 15013 2163
rect 14835 2095 14840 2129
rect 14840 2095 14906 2129
rect 14906 2095 14940 2129
rect 14940 2095 15013 2129
rect 14835 2061 15013 2095
rect 14835 2027 14840 2061
rect 14840 2027 14906 2061
rect 14906 2027 14940 2061
rect 14940 2027 15013 2061
rect 14835 1993 15013 2027
rect 14835 1959 14840 1993
rect 14840 1959 14906 1993
rect 14906 1959 14940 1993
rect 14940 1959 15013 1993
rect 14835 1925 15013 1959
rect 14835 1891 14840 1925
rect 14840 1891 14906 1925
rect 14906 1891 14940 1925
rect 14940 1891 15013 1925
rect 14835 1857 15013 1891
rect 14835 1823 14840 1857
rect 14840 1823 14906 1857
rect 14906 1823 14940 1857
rect 14940 1823 15013 1857
rect 14835 1789 15013 1823
rect 14835 1755 14840 1789
rect 14840 1755 14906 1789
rect 14906 1755 14940 1789
rect 14940 1755 15013 1789
rect 14835 1721 15013 1755
rect 14835 1687 14840 1721
rect 14840 1687 14906 1721
rect 14906 1687 14940 1721
rect 14940 1687 15013 1721
rect 14835 1653 15013 1687
rect 14835 1619 14840 1653
rect 14840 1619 14906 1653
rect 14906 1619 14940 1653
rect 14940 1619 15013 1653
rect 14835 1585 15013 1619
rect 14835 1551 14840 1585
rect 14840 1551 14906 1585
rect 14906 1551 14940 1585
rect 14940 1551 15013 1585
rect 14835 1517 15013 1551
rect 14835 1483 14840 1517
rect 14840 1483 14906 1517
rect 14906 1483 14940 1517
rect 14940 1483 15013 1517
rect 14835 1468 15013 1483
rect 14907 1449 15013 1468
rect 14835 1415 14840 1429
rect 14840 1415 14869 1429
rect 14907 1415 14940 1449
rect 14940 1415 15013 1449
rect 14835 1395 14869 1415
rect 14907 1381 15013 1415
rect 14835 1347 14840 1356
rect 14840 1347 14869 1356
rect 14907 1347 14940 1381
rect 14940 1347 15013 1381
rect 14835 1322 14869 1347
rect 14907 1313 15013 1347
rect 14835 1279 14840 1283
rect 14840 1279 14869 1283
rect 14907 1279 14940 1313
rect 14940 1279 15013 1313
rect 14835 1249 14869 1279
rect 14907 1245 15013 1279
rect 14907 1211 14940 1245
rect 14940 1211 15013 1245
rect 14835 1177 14869 1210
rect 14907 1177 15013 1211
rect 14835 1176 14840 1177
rect 14840 1176 14869 1177
rect 14907 1143 14940 1177
rect 14940 1143 15013 1177
rect 14835 1109 14869 1137
rect 14907 1109 15013 1143
rect 14835 1103 14840 1109
rect 14840 1103 14869 1109
rect 14907 1075 14940 1109
rect 14940 1075 15013 1109
rect 14835 1041 14869 1064
rect 14907 1041 15013 1075
rect 14835 1030 14840 1041
rect 14840 1030 14869 1041
rect 14907 1007 14940 1041
rect 14940 1007 15013 1041
rect 14835 973 14869 991
rect 14907 973 15013 1007
rect 14835 957 14840 973
rect 14840 957 14869 973
rect 14907 939 14940 973
rect 14940 939 15013 973
rect 14835 905 14869 918
rect 14907 905 15013 939
rect 14835 884 14840 905
rect 14840 884 14869 905
rect 14907 871 14940 905
rect 14940 871 15013 905
rect 14835 837 14869 845
rect 14907 837 15013 871
rect 14835 811 14840 837
rect 14840 811 14869 837
rect 14907 803 14940 837
rect 14940 803 15013 837
rect 14835 769 14869 772
rect 14907 769 15013 803
rect 14835 738 14840 769
rect 14840 738 14869 769
rect 14907 735 14940 769
rect 14940 735 15013 769
rect 14907 701 15013 735
rect 14835 667 14840 699
rect 14840 667 14869 699
rect 14907 667 14940 701
rect 14940 667 15013 701
rect 269 607 295 641
rect 295 607 303 641
rect 125 509 231 599
rect 269 533 303 567
rect 14835 665 14869 667
rect 14907 633 15013 667
rect 14835 599 14840 626
rect 14840 599 14869 626
rect 14907 599 14940 633
rect 14940 599 15013 633
rect 14835 592 14869 599
rect 14835 519 14869 553
rect 125 407 193 509
rect 193 407 231 509
rect 343 463 377 497
rect 419 463 453 497
rect 495 463 529 497
rect 571 463 605 497
rect 648 463 682 497
rect 14468 447 14502 481
rect 14542 447 14576 481
rect 14616 447 14650 481
rect 14689 447 14723 481
rect 14762 447 14796 481
rect 14907 420 15013 599
rect 125 331 231 407
rect 361 341 395 375
rect 434 341 468 375
rect 507 341 541 375
rect 580 341 614 375
rect 653 341 687 375
rect 726 341 760 375
rect 799 341 833 375
rect 872 341 906 375
rect 945 341 979 375
rect 1018 341 1052 375
rect 1091 341 1125 375
rect 1164 341 1198 375
rect 1237 341 1271 375
rect 1310 341 1344 375
rect 1383 341 1417 375
rect 1456 341 1490 375
rect 1529 341 1563 375
rect 1602 341 1636 375
rect 1675 341 1709 375
rect 1748 341 1782 375
rect 1821 341 1855 375
rect 1894 341 1928 375
rect 1967 341 2001 375
rect 2040 341 2074 375
rect 2113 341 2147 375
rect 2186 341 2220 375
rect 2259 341 2293 375
rect 2332 341 2366 375
rect 2405 341 2439 375
rect 2478 341 2512 375
rect 2551 341 2585 375
rect 2624 341 2658 375
rect 2697 341 2731 375
rect 2770 341 2804 375
rect 2843 341 2877 375
rect 2916 341 2950 375
rect 2989 341 3023 375
rect 3062 341 3096 375
rect 3135 341 3169 375
rect 3208 341 3242 375
rect 3281 341 3315 375
rect 3354 341 3388 375
rect 3427 341 3461 375
rect 3500 341 3534 375
rect 3573 341 3607 375
rect 3646 341 3680 375
rect 3719 341 3753 375
rect 3792 341 3826 375
rect 3865 341 3899 375
rect 3938 341 3972 375
rect 4011 341 4045 375
rect 4084 341 4118 375
rect 4157 341 4191 375
rect 4229 341 4263 375
rect 4301 341 4335 375
rect 4373 341 4407 375
rect 4445 341 4479 375
rect 4517 341 4551 375
rect 4589 341 4623 375
rect 4661 341 4695 375
rect 4733 341 4767 375
rect 4805 341 4839 375
rect 4877 341 4911 375
rect 4949 341 4983 375
rect 5021 341 5055 375
rect 5093 341 5127 375
rect 5165 341 5199 375
rect 5237 341 5271 375
rect 5309 341 5343 375
rect 5381 341 5415 375
rect 5453 341 5487 375
rect 5525 341 5559 375
rect 5597 341 5631 375
rect 5669 341 5703 375
rect 5741 341 5775 375
rect 5813 341 5847 375
rect 5885 341 5919 375
rect 5957 341 5991 375
rect 6029 341 6063 375
rect 6101 341 6135 375
rect 6173 341 6207 375
rect 6245 341 6279 375
rect 6317 341 6351 375
rect 6389 341 6423 375
rect 6461 341 6495 375
rect 6533 341 6567 375
rect 6605 341 6639 375
rect 6677 341 6711 375
rect 6749 341 6783 375
rect 6821 341 6855 375
rect 6893 341 6927 375
rect 6965 341 6999 375
rect 7037 341 7071 375
rect 7109 341 7143 375
rect 7181 341 7215 375
rect 7253 341 7287 375
rect 7325 341 7359 375
rect 7397 341 7431 375
rect 7469 341 7503 375
rect 7541 341 7575 375
rect 7613 341 7647 375
rect 7685 341 7719 375
rect 7757 341 7791 375
rect 7829 341 7863 375
rect 7901 341 7935 375
rect 7973 341 8007 375
rect 8045 341 8079 375
rect 8117 341 8151 375
rect 8189 341 8223 375
rect 8261 341 8295 375
rect 8333 341 8367 375
rect 8405 341 8439 375
rect 8477 341 8511 375
rect 8549 341 8583 375
rect 8621 341 8655 375
rect 8693 341 8727 375
rect 8765 341 8799 375
rect 8837 341 8871 375
rect 8909 341 8943 375
rect 8981 341 9015 375
rect 9053 341 9087 375
rect 9125 341 9159 375
rect 9197 341 9231 375
rect 9269 341 9303 375
rect 9341 341 9375 375
rect 9413 341 9447 375
rect 9485 341 9519 375
rect 9557 341 9591 375
rect 9629 341 9663 375
rect 9701 341 9735 375
rect 9773 341 9807 375
rect 9845 341 9879 375
rect 9917 341 9951 375
rect 9989 341 10023 375
rect 10061 341 10095 375
rect 10133 341 10167 375
rect 10205 341 10239 375
rect 10277 341 10311 375
rect 10349 341 10383 375
rect 10421 341 10455 375
rect 10493 341 10527 375
rect 10565 341 10599 375
rect 10637 341 10671 375
rect 10709 341 10743 375
rect 10781 341 10815 375
rect 10853 341 10887 375
rect 10925 341 10959 375
rect 10997 341 11031 375
rect 11069 341 11103 375
rect 11141 341 11175 375
rect 11213 341 11247 375
rect 11285 341 11319 375
rect 11357 341 11391 375
rect 11429 341 11463 375
rect 11501 341 11535 375
rect 11573 341 11607 375
rect 11645 341 11679 375
rect 11717 341 11751 375
rect 11789 341 11823 375
rect 11861 341 11895 375
rect 11933 341 11967 375
rect 12005 341 12039 375
rect 12077 341 12111 375
rect 12149 341 12183 375
rect 12221 341 12255 375
rect 12293 341 12327 375
rect 12365 341 12399 375
rect 12437 341 12471 375
rect 12509 341 12543 375
rect 12581 341 12615 375
rect 12653 341 12687 375
rect 12725 341 12759 375
rect 12797 341 12831 375
rect 12869 341 12903 375
rect 12941 341 12975 375
rect 13013 341 13047 375
rect 13085 341 13119 375
rect 13157 341 13191 375
rect 13229 341 13263 375
rect 13301 341 13335 375
rect 13373 341 13407 375
rect 13445 341 13479 375
rect 13517 341 13551 375
rect 13589 341 13623 375
rect 13661 341 13695 375
rect 13733 341 13767 375
rect 13805 341 13839 375
rect 13877 341 13911 375
rect 13949 341 13983 375
rect 14021 341 14055 375
rect 14093 341 14127 375
rect 14165 341 14199 375
rect 14237 341 14271 375
rect 14309 341 14343 375
rect 14381 341 14415 375
rect 14453 341 14487 375
rect 14525 341 14559 375
rect 14597 341 14631 375
rect 14669 341 14703 375
rect 14741 341 14775 375
<< metal1 >>
rect 39 5111 15097 5118
rect 39 5077 361 5111
rect 395 5077 434 5111
rect 468 5077 507 5111
rect 541 5077 580 5111
rect 614 5077 653 5111
rect 687 5077 726 5111
rect 760 5077 799 5111
rect 833 5077 872 5111
rect 906 5077 945 5111
rect 979 5077 1018 5111
rect 1052 5077 1091 5111
rect 1125 5077 1164 5111
rect 1198 5077 1237 5111
rect 1271 5077 1310 5111
rect 1344 5077 1383 5111
rect 1417 5077 1456 5111
rect 1490 5077 1529 5111
rect 1563 5077 1602 5111
rect 1636 5077 1675 5111
rect 1709 5077 1748 5111
rect 1782 5077 1821 5111
rect 1855 5077 1894 5111
rect 1928 5077 1967 5111
rect 2001 5077 2040 5111
rect 2074 5077 2113 5111
rect 2147 5077 2186 5111
rect 2220 5077 2259 5111
rect 2293 5077 2332 5111
rect 2366 5077 2405 5111
rect 2439 5077 2478 5111
rect 2512 5077 2551 5111
rect 2585 5077 2624 5111
rect 2658 5077 2697 5111
rect 2731 5077 2770 5111
rect 2804 5077 2843 5111
rect 2877 5077 2916 5111
rect 2950 5077 2989 5111
rect 3023 5077 3062 5111
rect 3096 5077 3135 5111
rect 3169 5077 3208 5111
rect 3242 5077 3281 5111
rect 3315 5077 3354 5111
rect 3388 5077 3427 5111
rect 3461 5077 3500 5111
rect 3534 5077 3573 5111
rect 3607 5077 3646 5111
rect 3680 5077 3719 5111
rect 3753 5077 3792 5111
rect 3826 5077 3865 5111
rect 3899 5077 3938 5111
rect 3972 5077 4011 5111
rect 4045 5077 4084 5111
rect 4118 5077 4157 5111
rect 4191 5077 4229 5111
rect 4263 5077 4301 5111
rect 4335 5077 4373 5111
rect 4407 5077 4445 5111
rect 4479 5077 4517 5111
rect 4551 5077 4589 5111
rect 4623 5077 4661 5111
rect 4695 5077 4733 5111
rect 4767 5077 4805 5111
rect 4839 5077 4877 5111
rect 4911 5077 4949 5111
rect 4983 5077 5021 5111
rect 5055 5077 5093 5111
rect 5127 5077 5165 5111
rect 5199 5077 5237 5111
rect 5271 5077 5309 5111
rect 5343 5077 5381 5111
rect 5415 5077 5453 5111
rect 5487 5077 5525 5111
rect 5559 5077 5597 5111
rect 5631 5077 5669 5111
rect 5703 5077 5741 5111
rect 5775 5077 5813 5111
rect 5847 5077 5885 5111
rect 5919 5077 5957 5111
rect 5991 5077 6029 5111
rect 6063 5077 6101 5111
rect 6135 5077 6173 5111
rect 6207 5077 6245 5111
rect 6279 5077 6317 5111
rect 6351 5077 6389 5111
rect 6423 5077 6461 5111
rect 6495 5077 6533 5111
rect 6567 5077 6605 5111
rect 6639 5077 6677 5111
rect 6711 5077 6749 5111
rect 6783 5077 6821 5111
rect 6855 5077 6893 5111
rect 6927 5077 6965 5111
rect 6999 5077 7037 5111
rect 7071 5077 7109 5111
rect 7143 5077 7181 5111
rect 7215 5077 7253 5111
rect 7287 5077 7325 5111
rect 7359 5077 7397 5111
rect 7431 5077 7469 5111
rect 7503 5077 7541 5111
rect 7575 5077 7613 5111
rect 7647 5077 7685 5111
rect 7719 5077 7757 5111
rect 7791 5077 7829 5111
rect 7863 5077 7901 5111
rect 7935 5077 7973 5111
rect 8007 5077 8045 5111
rect 8079 5077 8117 5111
rect 8151 5077 8189 5111
rect 8223 5077 8261 5111
rect 8295 5077 8333 5111
rect 8367 5077 8405 5111
rect 8439 5077 8477 5111
rect 8511 5077 8549 5111
rect 8583 5077 8621 5111
rect 8655 5077 8693 5111
rect 8727 5077 8765 5111
rect 8799 5077 8837 5111
rect 8871 5077 8909 5111
rect 8943 5077 8981 5111
rect 9015 5077 9053 5111
rect 9087 5077 9125 5111
rect 9159 5077 9197 5111
rect 9231 5077 9269 5111
rect 9303 5077 9341 5111
rect 9375 5077 9413 5111
rect 9447 5077 9485 5111
rect 9519 5077 9557 5111
rect 9591 5077 9629 5111
rect 9663 5077 9701 5111
rect 9735 5077 9773 5111
rect 9807 5077 9845 5111
rect 9879 5077 9917 5111
rect 9951 5077 9989 5111
rect 10023 5077 10061 5111
rect 10095 5077 10133 5111
rect 10167 5077 10205 5111
rect 10239 5077 10277 5111
rect 10311 5077 10349 5111
rect 10383 5077 10421 5111
rect 10455 5077 10493 5111
rect 10527 5077 10565 5111
rect 10599 5077 10637 5111
rect 10671 5077 10709 5111
rect 10743 5077 10781 5111
rect 10815 5077 10853 5111
rect 10887 5077 10925 5111
rect 10959 5077 10997 5111
rect 11031 5077 11069 5111
rect 11103 5077 11141 5111
rect 11175 5077 11213 5111
rect 11247 5077 11285 5111
rect 11319 5077 11357 5111
rect 11391 5077 11429 5111
rect 11463 5077 11501 5111
rect 11535 5077 11573 5111
rect 11607 5077 11645 5111
rect 11679 5077 11717 5111
rect 11751 5077 11789 5111
rect 11823 5077 11861 5111
rect 11895 5077 11933 5111
rect 11967 5077 12005 5111
rect 12039 5077 12077 5111
rect 12111 5077 12149 5111
rect 12183 5077 12221 5111
rect 12255 5077 12293 5111
rect 12327 5077 12365 5111
rect 12399 5077 12437 5111
rect 12471 5077 12509 5111
rect 12543 5077 12581 5111
rect 12615 5077 12653 5111
rect 12687 5077 12725 5111
rect 12759 5077 12797 5111
rect 12831 5077 12869 5111
rect 12903 5077 12941 5111
rect 12975 5077 13013 5111
rect 13047 5077 13085 5111
rect 13119 5077 13157 5111
rect 13191 5077 13229 5111
rect 13263 5077 13301 5111
rect 13335 5077 13373 5111
rect 13407 5077 13445 5111
rect 13479 5077 13517 5111
rect 13551 5077 13589 5111
rect 13623 5077 13661 5111
rect 13695 5077 13733 5111
rect 13767 5077 13805 5111
rect 13839 5077 13877 5111
rect 13911 5077 13949 5111
rect 13983 5077 14021 5111
rect 14055 5077 14093 5111
rect 14127 5077 14165 5111
rect 14199 5077 14237 5111
rect 14271 5077 14309 5111
rect 14343 5077 14381 5111
rect 14415 5077 14453 5111
rect 14487 5077 14525 5111
rect 14559 5077 14597 5111
rect 14631 5077 14669 5111
rect 14703 5077 14741 5111
rect 14775 5077 15097 5111
rect 39 5062 15097 5077
rect 39 5045 14907 5062
rect 39 331 125 5045
rect 231 5035 14907 5045
rect 231 5029 361 5035
rect 231 4995 269 5029
rect 303 5001 361 5029
rect 395 5001 434 5035
rect 468 5001 507 5035
rect 541 5001 580 5035
rect 614 5001 653 5035
rect 687 5001 726 5035
rect 760 5001 799 5035
rect 833 5001 872 5035
rect 906 5001 945 5035
rect 979 5001 1018 5035
rect 1052 5001 1091 5035
rect 1125 5001 1164 5035
rect 1198 5001 1237 5035
rect 1271 5001 1310 5035
rect 1344 5001 1383 5035
rect 1417 5001 1456 5035
rect 1490 5001 1529 5035
rect 1563 5001 1602 5035
rect 1636 5001 1675 5035
rect 1709 5001 1748 5035
rect 1782 5001 1821 5035
rect 1855 5001 1894 5035
rect 1928 5001 1967 5035
rect 2001 5001 2040 5035
rect 2074 5001 2113 5035
rect 2147 5001 2186 5035
rect 2220 5001 2259 5035
rect 2293 5001 2332 5035
rect 2366 5001 2405 5035
rect 2439 5001 2478 5035
rect 2512 5001 2551 5035
rect 2585 5001 2624 5035
rect 2658 5001 2697 5035
rect 2731 5001 2770 5035
rect 2804 5001 2843 5035
rect 2877 5001 2916 5035
rect 2950 5001 2989 5035
rect 3023 5001 3062 5035
rect 3096 5001 3135 5035
rect 3169 5001 3208 5035
rect 3242 5001 3281 5035
rect 3315 5001 3354 5035
rect 3388 5001 3427 5035
rect 3461 5001 3500 5035
rect 3534 5001 3573 5035
rect 3607 5001 3646 5035
rect 3680 5001 3719 5035
rect 3753 5001 3792 5035
rect 3826 5001 3865 5035
rect 3899 5001 3938 5035
rect 3972 5001 4011 5035
rect 4045 5001 4084 5035
rect 4118 5001 4157 5035
rect 4191 5001 4229 5035
rect 4263 5001 4301 5035
rect 4335 5001 4373 5035
rect 4407 5001 4445 5035
rect 4479 5001 4517 5035
rect 4551 5001 4589 5035
rect 4623 5001 4661 5035
rect 4695 5001 4733 5035
rect 4767 5001 4805 5035
rect 4839 5001 4877 5035
rect 4911 5001 4949 5035
rect 4983 5001 5021 5035
rect 5055 5001 5093 5035
rect 5127 5001 5165 5035
rect 5199 5001 5237 5035
rect 5271 5001 5309 5035
rect 5343 5001 5381 5035
rect 5415 5001 5453 5035
rect 5487 5001 5525 5035
rect 5559 5001 5597 5035
rect 5631 5001 5669 5035
rect 5703 5001 5741 5035
rect 5775 5001 5813 5035
rect 5847 5001 5885 5035
rect 5919 5001 5957 5035
rect 5991 5001 6029 5035
rect 6063 5001 6101 5035
rect 6135 5001 6173 5035
rect 6207 5001 6245 5035
rect 6279 5001 6317 5035
rect 6351 5001 6389 5035
rect 6423 5001 6461 5035
rect 6495 5001 6533 5035
rect 6567 5001 6605 5035
rect 6639 5001 6677 5035
rect 6711 5001 6749 5035
rect 6783 5001 6821 5035
rect 6855 5001 6893 5035
rect 6927 5001 6965 5035
rect 6999 5001 7037 5035
rect 7071 5001 7109 5035
rect 7143 5001 7181 5035
rect 7215 5001 7253 5035
rect 7287 5001 7325 5035
rect 7359 5001 7397 5035
rect 7431 5001 7469 5035
rect 7503 5001 7541 5035
rect 7575 5001 7613 5035
rect 7647 5001 7685 5035
rect 7719 5001 7757 5035
rect 7791 5001 7829 5035
rect 7863 5001 7901 5035
rect 7935 5001 7973 5035
rect 8007 5001 8045 5035
rect 8079 5001 8117 5035
rect 8151 5001 8189 5035
rect 8223 5001 8261 5035
rect 8295 5001 8333 5035
rect 8367 5001 8405 5035
rect 8439 5001 8477 5035
rect 8511 5001 8549 5035
rect 8583 5001 8621 5035
rect 8655 5001 8693 5035
rect 8727 5001 8765 5035
rect 8799 5001 8837 5035
rect 8871 5001 8909 5035
rect 8943 5001 8981 5035
rect 9015 5001 9053 5035
rect 9087 5001 9125 5035
rect 9159 5001 9197 5035
rect 9231 5001 9269 5035
rect 9303 5001 9341 5035
rect 9375 5001 9413 5035
rect 9447 5001 9485 5035
rect 9519 5001 9557 5035
rect 9591 5001 9629 5035
rect 9663 5001 9701 5035
rect 9735 5001 9773 5035
rect 9807 5001 9845 5035
rect 9879 5001 9917 5035
rect 9951 5001 9989 5035
rect 10023 5001 10061 5035
rect 10095 5001 10133 5035
rect 10167 5001 10205 5035
rect 10239 5001 10277 5035
rect 10311 5001 10349 5035
rect 10383 5001 10421 5035
rect 10455 5001 10493 5035
rect 10527 5001 10565 5035
rect 10599 5001 10637 5035
rect 10671 5001 10709 5035
rect 10743 5001 10781 5035
rect 10815 5001 10853 5035
rect 10887 5001 10925 5035
rect 10959 5001 10997 5035
rect 11031 5001 11069 5035
rect 11103 5001 11141 5035
rect 11175 5001 11213 5035
rect 11247 5001 11285 5035
rect 11319 5001 11357 5035
rect 11391 5001 11429 5035
rect 11463 5001 11501 5035
rect 11535 5001 11573 5035
rect 11607 5001 11645 5035
rect 11679 5001 11717 5035
rect 11751 5001 11789 5035
rect 11823 5001 11861 5035
rect 11895 5001 11933 5035
rect 11967 5001 12005 5035
rect 12039 5001 12077 5035
rect 12111 5001 12149 5035
rect 12183 5001 12221 5035
rect 12255 5001 12293 5035
rect 12327 5001 12365 5035
rect 12399 5001 12437 5035
rect 12471 5001 12509 5035
rect 12543 5001 12581 5035
rect 12615 5001 12653 5035
rect 12687 5001 12725 5035
rect 12759 5001 12797 5035
rect 12831 5001 12869 5035
rect 12903 5001 12941 5035
rect 12975 5001 13013 5035
rect 13047 5001 13085 5035
rect 13119 5001 13157 5035
rect 13191 5001 13229 5035
rect 13263 5001 13301 5035
rect 13335 5001 13373 5035
rect 13407 5001 13445 5035
rect 13479 5001 13517 5035
rect 13551 5001 13589 5035
rect 13623 5001 13661 5035
rect 13695 5001 13733 5035
rect 13767 5001 13805 5035
rect 13839 5001 13877 5035
rect 13911 5001 13949 5035
rect 13983 5001 14021 5035
rect 14055 5001 14093 5035
rect 14127 5001 14165 5035
rect 14199 5001 14237 5035
rect 14271 5001 14309 5035
rect 14343 5001 14381 5035
rect 14415 5001 14453 5035
rect 14487 5001 14525 5035
rect 14559 5001 14597 5035
rect 14631 5001 14669 5035
rect 14703 5001 14741 5035
rect 14775 5030 14907 5035
rect 14775 5001 14835 5030
rect 303 4995 14835 5001
rect 231 4959 14835 4995
rect 231 4956 361 4959
rect 231 4922 269 4956
rect 303 4925 361 4956
rect 395 4925 434 4959
rect 468 4925 507 4959
rect 541 4925 580 4959
rect 614 4925 653 4959
rect 687 4925 726 4959
rect 760 4925 799 4959
rect 833 4925 872 4959
rect 906 4925 945 4959
rect 979 4925 1018 4959
rect 1052 4925 1091 4959
rect 1125 4925 1164 4959
rect 1198 4925 1237 4959
rect 1271 4925 1310 4959
rect 1344 4925 1383 4959
rect 1417 4925 1456 4959
rect 1490 4925 1529 4959
rect 1563 4925 1602 4959
rect 1636 4925 1675 4959
rect 1709 4925 1748 4959
rect 1782 4925 1821 4959
rect 1855 4925 1894 4959
rect 1928 4925 1967 4959
rect 2001 4925 2040 4959
rect 2074 4925 2113 4959
rect 2147 4925 2186 4959
rect 2220 4925 2259 4959
rect 2293 4925 2332 4959
rect 2366 4925 2405 4959
rect 2439 4925 2478 4959
rect 2512 4925 2551 4959
rect 2585 4925 2624 4959
rect 2658 4925 2697 4959
rect 2731 4925 2770 4959
rect 2804 4925 2843 4959
rect 2877 4925 2916 4959
rect 2950 4925 2989 4959
rect 3023 4925 3062 4959
rect 3096 4925 3135 4959
rect 3169 4925 3208 4959
rect 3242 4925 3281 4959
rect 3315 4925 3354 4959
rect 3388 4925 3427 4959
rect 3461 4925 3500 4959
rect 3534 4925 3573 4959
rect 3607 4925 3646 4959
rect 3680 4925 3719 4959
rect 3753 4925 3792 4959
rect 3826 4925 3865 4959
rect 3899 4925 3938 4959
rect 3972 4925 4011 4959
rect 4045 4925 4084 4959
rect 4118 4925 4157 4959
rect 4191 4925 4229 4959
rect 4263 4925 4301 4959
rect 4335 4925 4373 4959
rect 4407 4925 4445 4959
rect 4479 4925 4517 4959
rect 4551 4925 4589 4959
rect 4623 4925 4661 4959
rect 4695 4925 4733 4959
rect 4767 4925 4805 4959
rect 4839 4925 4877 4959
rect 4911 4925 4949 4959
rect 4983 4925 5021 4959
rect 5055 4925 5093 4959
rect 5127 4925 5165 4959
rect 5199 4925 5237 4959
rect 5271 4925 5309 4959
rect 5343 4925 5381 4959
rect 5415 4925 5453 4959
rect 5487 4925 5525 4959
rect 5559 4925 5597 4959
rect 5631 4925 5669 4959
rect 5703 4925 5741 4959
rect 5775 4925 5813 4959
rect 5847 4925 5885 4959
rect 5919 4925 5957 4959
rect 5991 4925 6029 4959
rect 6063 4925 6101 4959
rect 6135 4925 6173 4959
rect 6207 4925 6245 4959
rect 6279 4925 6317 4959
rect 6351 4925 6389 4959
rect 6423 4925 6461 4959
rect 6495 4925 6533 4959
rect 6567 4925 6605 4959
rect 6639 4925 6677 4959
rect 6711 4925 6749 4959
rect 6783 4925 6821 4959
rect 6855 4925 6893 4959
rect 6927 4925 6965 4959
rect 6999 4925 7037 4959
rect 7071 4925 7109 4959
rect 7143 4925 7181 4959
rect 7215 4925 7253 4959
rect 7287 4925 7325 4959
rect 7359 4925 7397 4959
rect 7431 4925 7469 4959
rect 7503 4925 7541 4959
rect 7575 4925 7613 4959
rect 7647 4925 7685 4959
rect 7719 4925 7757 4959
rect 7791 4925 7829 4959
rect 7863 4925 7901 4959
rect 7935 4925 7973 4959
rect 8007 4925 8045 4959
rect 8079 4925 8117 4959
rect 8151 4925 8189 4959
rect 8223 4925 8261 4959
rect 8295 4925 8333 4959
rect 8367 4925 8405 4959
rect 8439 4925 8477 4959
rect 8511 4925 8549 4959
rect 8583 4925 8621 4959
rect 8655 4925 8693 4959
rect 8727 4925 8765 4959
rect 8799 4925 8837 4959
rect 8871 4925 8909 4959
rect 8943 4925 8981 4959
rect 9015 4925 9053 4959
rect 9087 4925 9125 4959
rect 9159 4925 9197 4959
rect 9231 4925 9269 4959
rect 9303 4925 9341 4959
rect 9375 4925 9413 4959
rect 9447 4925 9485 4959
rect 9519 4925 9557 4959
rect 9591 4925 9629 4959
rect 9663 4925 9701 4959
rect 9735 4925 9773 4959
rect 9807 4925 9845 4959
rect 9879 4925 9917 4959
rect 9951 4925 9989 4959
rect 10023 4925 10061 4959
rect 10095 4925 10133 4959
rect 10167 4925 10205 4959
rect 10239 4925 10277 4959
rect 10311 4925 10349 4959
rect 10383 4925 10421 4959
rect 10455 4925 10493 4959
rect 10527 4925 10565 4959
rect 10599 4925 10637 4959
rect 10671 4925 10709 4959
rect 10743 4925 10781 4959
rect 10815 4925 10853 4959
rect 10887 4925 10925 4959
rect 10959 4925 10997 4959
rect 11031 4925 11069 4959
rect 11103 4925 11141 4959
rect 11175 4925 11213 4959
rect 11247 4925 11285 4959
rect 11319 4925 11357 4959
rect 11391 4925 11429 4959
rect 11463 4925 11501 4959
rect 11535 4925 11573 4959
rect 11607 4925 11645 4959
rect 11679 4925 11717 4959
rect 11751 4925 11789 4959
rect 11823 4925 11861 4959
rect 11895 4925 11933 4959
rect 11967 4925 12005 4959
rect 12039 4925 12077 4959
rect 12111 4925 12149 4959
rect 12183 4925 12221 4959
rect 12255 4925 12293 4959
rect 12327 4925 12365 4959
rect 12399 4925 12437 4959
rect 12471 4925 12509 4959
rect 12543 4925 12581 4959
rect 12615 4925 12653 4959
rect 12687 4925 12725 4959
rect 12759 4925 12797 4959
rect 12831 4925 12869 4959
rect 12903 4925 12941 4959
rect 12975 4925 13013 4959
rect 13047 4925 13085 4959
rect 13119 4925 13157 4959
rect 13191 4925 13229 4959
rect 13263 4925 13301 4959
rect 13335 4925 13373 4959
rect 13407 4925 13445 4959
rect 13479 4925 13517 4959
rect 13551 4925 13589 4959
rect 13623 4925 13661 4959
rect 13695 4925 13733 4959
rect 13767 4925 13805 4959
rect 13839 4925 13877 4959
rect 13911 4925 13949 4959
rect 13983 4925 14021 4959
rect 14055 4925 14093 4959
rect 14127 4925 14165 4959
rect 14199 4925 14237 4959
rect 14271 4925 14309 4959
rect 14343 4925 14381 4959
rect 14415 4925 14453 4959
rect 14487 4925 14525 4959
rect 14559 4925 14597 4959
rect 14631 4925 14669 4959
rect 14703 4925 14741 4959
rect 14775 4925 14835 4959
rect 303 4922 14835 4925
rect 231 4918 14835 4922
rect 231 4883 491 4918
rect 231 4849 269 4883
rect 303 4849 491 4883
rect 231 4810 491 4849
rect 231 4776 269 4810
rect 303 4776 491 4810
rect 231 4737 491 4776
rect 231 4703 269 4737
rect 303 4703 491 4737
rect 231 4664 491 4703
rect 231 4630 269 4664
rect 303 4630 491 4664
rect 231 4618 491 4630
tri 491 4618 791 4918 nw
tri 14335 4618 14635 4918 ne
rect 14635 4618 14835 4918
rect 231 4606 479 4618
tri 479 4606 491 4618 nw
tri 621 4606 633 4618 se
rect 633 4606 14502 4618
rect 231 4591 373 4606
rect 231 4557 269 4591
rect 303 4557 373 4591
rect 231 4518 373 4557
rect 231 4484 269 4518
rect 303 4500 373 4518
tri 373 4500 479 4606 nw
tri 517 4502 621 4606 se
rect 621 4502 709 4606
rect 517 4500 709 4502
rect 14207 4572 14246 4606
rect 14280 4572 14319 4606
rect 14353 4572 14392 4606
rect 14426 4572 14502 4606
rect 14207 4534 14502 4572
rect 14207 4500 14246 4534
rect 14280 4500 14319 4534
rect 14353 4500 14392 4534
rect 14426 4502 14502 4534
tri 14502 4502 14618 4618 sw
rect 14426 4500 14618 4502
rect 303 4484 329 4500
rect 231 4445 329 4484
tri 329 4456 373 4500 nw
rect 517 4488 14618 4500
rect 517 4456 946 4488
tri 946 4456 978 4488 nw
tri 14157 4468 14177 4488 ne
rect 14177 4468 14618 4488
tri 14177 4456 14189 4468 ne
rect 14189 4456 14618 4468
rect 231 4411 269 4445
rect 303 4411 329 4445
rect 231 4372 329 4411
rect 231 4338 269 4372
rect 303 4338 329 4372
rect 231 4299 329 4338
rect 231 4265 269 4299
rect 303 4265 329 4299
rect 231 4226 329 4265
rect 231 4192 269 4226
rect 303 4192 329 4226
rect 231 4153 329 4192
rect 231 4119 269 4153
rect 303 4119 329 4153
rect 231 4080 329 4119
rect 231 4046 269 4080
rect 303 4046 329 4080
rect 231 4007 329 4046
rect 231 3973 269 4007
rect 303 3973 329 4007
rect 231 3934 329 3973
rect 231 3900 269 3934
rect 303 3900 329 3934
rect 231 3861 329 3900
rect 231 3827 269 3861
rect 303 3827 329 3861
rect 231 3788 329 3827
rect 231 3754 269 3788
rect 303 3754 329 3788
rect 231 3715 329 3754
rect 231 3681 269 3715
rect 303 3681 329 3715
rect 231 3642 329 3681
rect 231 3608 269 3642
rect 303 3608 329 3642
rect 231 3569 329 3608
rect 231 3535 269 3569
rect 303 3535 329 3569
rect 231 3496 329 3535
rect 231 3462 269 3496
rect 303 3462 329 3496
rect 231 3423 329 3462
rect 231 3389 269 3423
rect 303 3389 329 3423
rect 231 3350 329 3389
rect 231 3316 269 3350
rect 303 3316 329 3350
rect 231 3277 329 3316
rect 231 3243 269 3277
rect 303 3243 329 3277
rect 231 3204 329 3243
rect 231 3170 269 3204
rect 303 3170 329 3204
rect 231 3131 329 3170
rect 231 3097 269 3131
rect 303 3097 329 3131
rect 231 3058 329 3097
rect 231 3024 269 3058
rect 303 3024 329 3058
rect 231 2985 329 3024
rect 231 2951 269 2985
rect 303 2951 329 2985
rect 231 2912 329 2951
rect 231 2878 269 2912
rect 303 2878 329 2912
rect 231 2839 329 2878
rect 231 2805 269 2839
rect 303 2805 329 2839
rect 231 2766 329 2805
rect 231 2732 269 2766
rect 303 2732 329 2766
rect 231 2693 329 2732
rect 231 2659 269 2693
rect 303 2659 329 2693
rect 231 2620 329 2659
rect 231 2586 269 2620
rect 303 2586 329 2620
rect 231 2547 329 2586
rect 231 2513 269 2547
rect 303 2513 329 2547
rect 231 2474 329 2513
rect 231 2440 269 2474
rect 303 2440 329 2474
rect 231 2401 329 2440
rect 231 2367 269 2401
rect 303 2367 329 2401
rect 231 2328 329 2367
rect 231 2294 269 2328
rect 303 2294 329 2328
rect 231 2255 329 2294
rect 231 2221 269 2255
rect 303 2221 329 2255
rect 231 2182 329 2221
rect 231 2148 269 2182
rect 303 2148 329 2182
rect 231 2109 329 2148
rect 231 2075 269 2109
rect 303 2075 329 2109
rect 231 2036 329 2075
rect 231 2002 269 2036
rect 303 2002 329 2036
rect 231 1963 329 2002
rect 231 1929 269 1963
rect 303 1929 329 1963
rect 231 1890 329 1929
rect 231 1856 269 1890
rect 303 1856 329 1890
rect 231 1817 329 1856
rect 231 1783 269 1817
rect 303 1783 329 1817
rect 231 1744 329 1783
rect 231 1710 269 1744
rect 303 1710 329 1744
rect 231 1671 329 1710
rect 231 1637 269 1671
rect 303 1637 329 1671
rect 231 1598 329 1637
rect 231 1564 269 1598
rect 303 1564 329 1598
rect 231 1525 329 1564
rect 231 1491 269 1525
rect 303 1491 329 1525
rect 231 1452 329 1491
rect 231 1418 269 1452
rect 303 1418 329 1452
rect 231 1379 329 1418
rect 231 1345 269 1379
rect 303 1345 329 1379
rect 231 1306 329 1345
rect 231 1272 269 1306
rect 303 1272 329 1306
rect 231 1233 329 1272
rect 231 1199 269 1233
rect 303 1199 329 1233
rect 231 1159 329 1199
rect 231 1125 269 1159
rect 303 1125 329 1159
rect 231 1085 329 1125
rect 231 1051 269 1085
rect 303 1051 329 1085
rect 231 1011 329 1051
rect 231 977 269 1011
rect 303 977 329 1011
rect 231 937 329 977
rect 231 903 269 937
rect 303 903 329 937
rect 231 863 329 903
rect 517 4404 518 4456
rect 570 4404 590 4456
rect 642 4404 662 4456
rect 714 4445 734 4456
rect 786 4448 938 4456
tri 938 4448 946 4456 nw
tri 14189 4448 14197 4456 ne
rect 14197 4448 14428 4456
rect 786 4432 922 4448
tri 922 4432 938 4448 nw
tri 14197 4444 14201 4448 ne
rect 14201 4444 14428 4448
tri 14201 4432 14213 4444 ne
rect 14213 4432 14428 4444
rect 786 4404 888 4432
rect 517 4392 529 4404
rect 563 4392 601 4404
rect 635 4392 674 4404
rect 517 4390 674 4392
rect 780 4398 888 4404
tri 888 4398 922 4432 nw
tri 14213 4398 14247 4432 ne
rect 14247 4398 14356 4432
rect 14390 4398 14428 4432
rect 14462 4426 14618 4456
tri 14635 4446 14807 4618 ne
rect 780 4390 849 4398
rect 517 4338 518 4390
rect 570 4338 590 4390
rect 642 4338 662 4390
rect 786 4359 849 4390
tri 849 4359 888 4398 nw
tri 14247 4359 14286 4398 ne
rect 14286 4359 14428 4398
rect 786 4338 815 4359
rect 517 4325 529 4338
rect 563 4325 601 4338
rect 635 4325 674 4338
rect 780 4325 815 4338
tri 815 4325 849 4359 nw
tri 14286 4325 14320 4359 ne
rect 14320 4325 14356 4359
rect 14390 4325 14428 4359
rect 517 4273 518 4325
rect 570 4273 590 4325
rect 642 4273 662 4325
tri 786 4296 815 4325 nw
tri 14320 4296 14349 4325 ne
rect 14349 4296 14428 4325
tri 14349 4295 14350 4296 ne
rect 517 4260 529 4273
rect 563 4260 601 4273
rect 635 4260 674 4273
rect 780 4260 786 4273
rect 517 4208 518 4260
rect 570 4208 590 4260
rect 642 4208 662 4260
rect 517 4201 674 4208
rect 517 4195 529 4201
rect 563 4195 601 4201
rect 635 4195 674 4201
rect 780 4195 786 4208
rect 517 4143 518 4195
rect 570 4143 590 4195
rect 642 4143 662 4195
rect 517 4130 674 4143
rect 780 4130 786 4143
rect 14350 4286 14428 4296
rect 14350 4252 14356 4286
rect 14390 4252 14428 4286
rect 14350 4213 14428 4252
rect 14350 4179 14356 4213
rect 14390 4179 14428 4213
rect 14350 4140 14428 4179
rect 517 4078 518 4130
rect 570 4078 590 4130
rect 642 4078 662 4130
rect 517 4065 674 4078
rect 780 4065 786 4078
rect 517 4013 518 4065
rect 570 4013 590 4065
rect 642 4013 662 4065
rect 517 4000 674 4013
rect 780 4000 786 4013
rect 517 3948 518 4000
rect 570 3948 590 4000
rect 642 3948 662 4000
rect 517 3944 529 3948
rect 563 3944 601 3948
rect 635 3944 674 3948
rect 517 3935 674 3944
rect 780 3935 786 3948
rect 517 3883 518 3935
rect 570 3883 590 3935
rect 642 3883 662 3935
rect 517 3870 529 3883
rect 563 3870 601 3883
rect 635 3870 674 3883
rect 780 3870 786 3883
rect 517 3818 518 3870
rect 570 3818 590 3870
rect 642 3818 662 3870
rect 517 3805 674 3818
rect 780 3805 786 3818
rect 517 3753 518 3805
rect 570 3753 590 3805
rect 642 3753 662 3805
rect 517 3740 674 3753
rect 780 3740 786 3753
rect 517 3688 518 3740
rect 570 3688 590 3740
rect 642 3688 662 3740
rect 517 3686 529 3688
rect 563 3686 601 3688
rect 635 3686 674 3688
rect 517 3675 674 3686
rect 780 3675 786 3688
rect 517 3623 518 3675
rect 570 3623 590 3675
rect 642 3623 662 3675
rect 517 3612 529 3623
rect 563 3612 601 3623
rect 635 3612 674 3623
rect 517 3610 674 3612
rect 780 3610 786 3623
rect 517 3558 518 3610
rect 570 3558 590 3610
rect 642 3558 662 3610
rect 517 3545 529 3558
rect 563 3545 601 3558
rect 635 3545 674 3558
rect 780 3545 786 3558
rect 517 3493 518 3545
rect 570 3493 590 3545
rect 642 3493 662 3545
rect 517 3480 529 3493
rect 563 3480 601 3493
rect 635 3480 674 3493
rect 780 3480 786 3493
rect 517 3428 518 3480
rect 570 3428 590 3480
rect 642 3428 662 3480
rect 517 3424 674 3428
rect 517 3415 529 3424
rect 563 3415 601 3424
rect 635 3415 674 3424
rect 780 3415 786 3428
rect 517 3363 518 3415
rect 570 3363 590 3415
rect 642 3363 662 3415
rect 517 3350 674 3363
rect 780 3350 786 3363
rect 517 3298 518 3350
rect 570 3298 590 3350
rect 642 3298 662 3350
rect 517 3285 674 3298
rect 780 3285 786 3298
rect 517 3233 518 3285
rect 570 3233 590 3285
rect 642 3233 662 3285
rect 517 3220 674 3233
rect 780 3220 786 3233
rect 517 3168 518 3220
rect 570 3168 590 3220
rect 642 3168 662 3220
rect 517 3155 674 3168
rect 780 3155 786 3168
rect 517 3103 518 3155
rect 570 3103 590 3155
rect 642 3103 662 3155
rect 517 3094 529 3103
rect 563 3094 601 3103
rect 635 3094 674 3103
rect 517 3090 674 3094
rect 780 3090 786 3103
rect 517 3038 518 3090
rect 570 3038 590 3090
rect 642 3038 662 3090
rect 517 3025 529 3038
rect 563 3025 601 3038
rect 635 3025 674 3038
rect 780 3025 786 3038
rect 517 2973 518 3025
rect 570 2973 590 3025
rect 642 2973 662 3025
rect 517 2960 529 2973
rect 563 2960 601 2973
rect 635 2960 674 2973
rect 780 2960 786 2973
rect 517 2908 518 2960
rect 570 2908 590 2960
rect 642 2908 662 2960
rect 517 2906 674 2908
rect 517 2895 529 2906
rect 563 2895 601 2906
rect 635 2895 674 2906
rect 780 2895 786 2908
rect 517 2843 518 2895
rect 570 2843 590 2895
rect 642 2843 662 2895
rect 517 2832 674 2843
rect 517 2830 529 2832
rect 563 2830 601 2832
rect 635 2830 674 2832
rect 780 2830 786 2843
rect 517 2778 518 2830
rect 570 2778 590 2830
rect 642 2778 662 2830
rect 517 2765 674 2778
rect 780 2765 786 2778
rect 517 2713 518 2765
rect 570 2713 590 2765
rect 642 2713 662 2765
rect 517 2700 674 2713
rect 780 2700 786 2713
rect 517 2648 518 2700
rect 570 2648 590 2700
rect 642 2648 662 2700
rect 517 2635 674 2648
rect 780 2635 786 2648
rect 517 2583 518 2635
rect 570 2583 590 2635
rect 642 2583 662 2635
rect 517 2576 529 2583
rect 563 2576 601 2583
rect 635 2576 674 2583
rect 517 2570 674 2576
rect 780 2570 786 2583
rect 517 2518 518 2570
rect 570 2518 590 2570
rect 642 2518 662 2570
rect 517 2505 529 2518
rect 563 2505 601 2518
rect 635 2505 674 2518
rect 780 2505 786 2518
rect 517 2453 518 2505
rect 570 2453 590 2505
rect 642 2453 662 2505
rect 517 2440 529 2453
rect 563 2440 601 2453
rect 635 2440 674 2453
rect 780 2440 786 2453
rect 517 2388 518 2440
rect 570 2388 590 2440
rect 642 2388 662 2440
rect 517 2375 529 2388
rect 563 2375 601 2388
rect 635 2375 674 2388
rect 780 2375 786 2388
rect 517 2323 518 2375
rect 570 2323 590 2375
rect 642 2323 662 2375
rect 517 2316 674 2323
rect 517 2310 529 2316
rect 563 2310 601 2316
rect 635 2310 674 2316
rect 780 2310 786 2323
rect 517 2258 518 2310
rect 570 2258 590 2310
rect 642 2258 662 2310
rect 517 2245 674 2258
rect 780 2245 786 2258
rect 517 2193 518 2245
rect 570 2193 590 2245
rect 642 2193 662 2245
rect 517 2180 674 2193
rect 780 2180 786 2193
rect 517 2128 518 2180
rect 570 2128 590 2180
rect 642 2128 662 2180
rect 517 2115 674 2128
rect 780 2115 786 2128
rect 517 2063 518 2115
rect 570 2063 590 2115
rect 642 2063 662 2115
rect 517 2050 674 2063
rect 780 2050 786 2063
rect 517 1998 518 2050
rect 570 1998 590 2050
rect 642 1998 662 2050
rect 517 1990 529 1998
rect 563 1990 601 1998
rect 635 1990 674 1998
rect 517 1985 674 1990
rect 780 1985 786 1998
rect 517 1933 518 1985
rect 570 1933 590 1985
rect 642 1933 662 1985
rect 517 1920 529 1933
rect 563 1920 601 1933
rect 635 1920 674 1933
rect 780 1920 786 1933
rect 517 1868 518 1920
rect 570 1868 590 1920
rect 642 1868 662 1920
rect 517 1855 529 1868
rect 563 1855 601 1868
rect 635 1855 674 1868
rect 780 1855 786 1868
rect 517 1803 518 1855
rect 570 1803 590 1855
rect 642 1803 662 1855
rect 517 1790 529 1803
rect 563 1790 601 1803
rect 635 1790 674 1803
rect 780 1790 786 1803
rect 517 1738 518 1790
rect 570 1738 590 1790
rect 642 1738 662 1790
rect 517 1732 674 1738
rect 517 1725 529 1732
rect 563 1725 601 1732
rect 635 1725 674 1732
rect 780 1725 786 1738
rect 517 1673 518 1725
rect 570 1673 590 1725
rect 642 1673 662 1725
rect 517 1660 674 1673
rect 780 1660 786 1673
rect 517 1608 518 1660
rect 570 1608 590 1660
rect 642 1608 662 1660
rect 517 1595 674 1608
rect 780 1595 786 1608
rect 517 1543 518 1595
rect 570 1543 590 1595
rect 642 1543 662 1595
rect 1060 4119 1252 4125
rect 1060 4067 1066 4119
rect 1118 4067 1130 4119
rect 1182 4067 1194 4119
rect 1246 4067 1252 4119
rect 1060 4064 1067 4067
rect 1101 4064 1139 4067
rect 1173 4064 1211 4067
rect 1245 4064 1252 4067
rect 1060 4054 1252 4064
rect 1060 4002 1066 4054
rect 1118 4002 1130 4054
rect 1182 4002 1194 4054
rect 1246 4002 1252 4054
rect 1060 3991 1067 4002
rect 1101 3991 1139 4002
rect 1173 3991 1211 4002
rect 1245 3991 1252 4002
rect 1060 3989 1252 3991
rect 1060 3937 1066 3989
rect 1118 3937 1130 3989
rect 1182 3937 1194 3989
rect 1246 3937 1252 3989
rect 1060 3924 1067 3937
rect 1101 3924 1139 3937
rect 1173 3924 1211 3937
rect 1245 3924 1252 3937
rect 1060 1568 1066 3924
rect 1246 1568 1252 3924
rect 1060 1562 1252 1568
rect 1556 4124 1748 4130
rect 1556 4072 1562 4124
rect 1614 4092 1626 4124
rect 1678 4092 1690 4124
rect 1742 4072 1748 4124
rect 1556 4059 1563 4072
rect 1741 4059 1748 4072
rect 1556 4007 1562 4059
rect 1742 4007 1748 4059
rect 1556 3994 1563 4007
rect 1741 3994 1748 4007
rect 1556 3942 1562 3994
rect 1742 3942 1748 3994
rect 1556 3929 1563 3942
rect 1741 3929 1748 3942
rect 1556 3877 1562 3929
rect 1742 3877 1748 3929
rect 1556 3864 1563 3877
rect 1741 3864 1748 3877
rect 1556 3812 1562 3864
rect 1742 3812 1748 3864
rect 1556 3799 1563 3812
rect 1741 3799 1748 3812
rect 1556 3747 1562 3799
rect 1742 3747 1748 3799
rect 1556 3734 1563 3747
rect 1741 3734 1748 3747
rect 1556 3682 1562 3734
rect 1742 3682 1748 3734
rect 1556 3669 1563 3682
rect 1741 3669 1748 3682
rect 1556 3617 1562 3669
rect 1742 3617 1748 3669
rect 1556 3604 1563 3617
rect 1741 3604 1748 3617
rect 1556 1568 1562 3604
rect 1742 1568 1748 3604
rect 1556 1562 1748 1568
rect 2052 4119 2244 4125
rect 2052 4067 2058 4119
rect 2110 4067 2122 4119
rect 2174 4067 2186 4119
rect 2238 4067 2244 4119
rect 2052 4064 2059 4067
rect 2093 4064 2131 4067
rect 2165 4064 2203 4067
rect 2237 4064 2244 4067
rect 2052 4054 2244 4064
rect 2052 4002 2058 4054
rect 2110 4002 2122 4054
rect 2174 4002 2186 4054
rect 2238 4002 2244 4054
rect 2052 3991 2059 4002
rect 2093 3991 2131 4002
rect 2165 3991 2203 4002
rect 2237 3991 2244 4002
rect 2052 3989 2244 3991
rect 2052 3937 2058 3989
rect 2110 3937 2122 3989
rect 2174 3937 2186 3989
rect 2238 3937 2244 3989
rect 2052 3924 2059 3937
rect 2093 3924 2131 3937
rect 2165 3924 2203 3937
rect 2237 3924 2244 3937
rect 2052 1568 2058 3924
rect 2238 1568 2244 3924
rect 2052 1562 2244 1568
rect 2548 4124 2740 4130
rect 2548 4072 2554 4124
rect 2606 4092 2618 4124
rect 2670 4092 2682 4124
rect 2734 4072 2740 4124
rect 2548 4059 2555 4072
rect 2733 4059 2740 4072
rect 2548 4007 2554 4059
rect 2734 4007 2740 4059
rect 2548 3994 2555 4007
rect 2733 3994 2740 4007
rect 2548 3942 2554 3994
rect 2734 3942 2740 3994
rect 2548 3929 2555 3942
rect 2733 3929 2740 3942
rect 2548 3877 2554 3929
rect 2734 3877 2740 3929
rect 2548 3864 2555 3877
rect 2733 3864 2740 3877
rect 2548 3812 2554 3864
rect 2734 3812 2740 3864
rect 2548 3799 2555 3812
rect 2733 3799 2740 3812
rect 2548 3747 2554 3799
rect 2734 3747 2740 3799
rect 2548 3734 2555 3747
rect 2733 3734 2740 3747
rect 2548 3682 2554 3734
rect 2734 3682 2740 3734
rect 2548 3669 2555 3682
rect 2733 3669 2740 3682
rect 2548 3617 2554 3669
rect 2734 3617 2740 3669
rect 2548 3604 2555 3617
rect 2733 3604 2740 3617
rect 2548 1568 2554 3604
rect 2734 1568 2740 3604
rect 2548 1562 2740 1568
rect 3044 4119 3236 4125
rect 3044 4067 3050 4119
rect 3102 4067 3114 4119
rect 3166 4067 3178 4119
rect 3230 4067 3236 4119
rect 3044 4064 3051 4067
rect 3085 4064 3123 4067
rect 3157 4064 3195 4067
rect 3229 4064 3236 4067
rect 3044 4054 3236 4064
rect 3044 4002 3050 4054
rect 3102 4002 3114 4054
rect 3166 4002 3178 4054
rect 3230 4002 3236 4054
rect 3044 3991 3051 4002
rect 3085 3991 3123 4002
rect 3157 3991 3195 4002
rect 3229 3991 3236 4002
rect 3044 3989 3236 3991
rect 3044 3937 3050 3989
rect 3102 3937 3114 3989
rect 3166 3937 3178 3989
rect 3230 3937 3236 3989
rect 3044 3924 3051 3937
rect 3085 3924 3123 3937
rect 3157 3924 3195 3937
rect 3229 3924 3236 3937
rect 3044 1568 3050 3924
rect 3230 1568 3236 3924
rect 3044 1562 3236 1568
rect 3540 4124 3732 4130
rect 3540 4072 3546 4124
rect 3598 4092 3610 4124
rect 3662 4092 3674 4124
rect 3726 4072 3732 4124
rect 3540 4059 3547 4072
rect 3725 4059 3732 4072
rect 3540 4007 3546 4059
rect 3726 4007 3732 4059
rect 3540 3994 3547 4007
rect 3725 3994 3732 4007
rect 3540 3942 3546 3994
rect 3726 3942 3732 3994
rect 3540 3929 3547 3942
rect 3725 3929 3732 3942
rect 3540 3877 3546 3929
rect 3726 3877 3732 3929
rect 3540 3864 3547 3877
rect 3725 3864 3732 3877
rect 3540 3812 3546 3864
rect 3726 3812 3732 3864
rect 3540 3799 3547 3812
rect 3725 3799 3732 3812
rect 3540 3747 3546 3799
rect 3726 3747 3732 3799
rect 3540 3734 3547 3747
rect 3725 3734 3732 3747
rect 3540 3682 3546 3734
rect 3726 3682 3732 3734
rect 3540 3669 3547 3682
rect 3725 3669 3732 3682
rect 3540 3617 3546 3669
rect 3726 3617 3732 3669
rect 3540 3604 3547 3617
rect 3725 3604 3732 3617
rect 3540 1568 3546 3604
rect 3726 1568 3732 3604
rect 3540 1562 3732 1568
rect 4036 4119 4228 4125
rect 4036 4067 4042 4119
rect 4094 4067 4106 4119
rect 4158 4067 4170 4119
rect 4222 4067 4228 4119
rect 4036 4064 4043 4067
rect 4077 4064 4115 4067
rect 4149 4064 4187 4067
rect 4221 4064 4228 4067
rect 4036 4054 4228 4064
rect 4036 4002 4042 4054
rect 4094 4002 4106 4054
rect 4158 4002 4170 4054
rect 4222 4002 4228 4054
rect 4036 3991 4043 4002
rect 4077 3991 4115 4002
rect 4149 3991 4187 4002
rect 4221 3991 4228 4002
rect 4036 3989 4228 3991
rect 4036 3937 4042 3989
rect 4094 3937 4106 3989
rect 4158 3937 4170 3989
rect 4222 3937 4228 3989
rect 4036 3924 4043 3937
rect 4077 3924 4115 3937
rect 4149 3924 4187 3937
rect 4221 3924 4228 3937
rect 4036 1568 4042 3924
rect 4222 1568 4228 3924
rect 4036 1562 4228 1568
rect 4532 4124 4724 4130
rect 4532 4072 4538 4124
rect 4590 4092 4602 4124
rect 4654 4092 4666 4124
rect 4718 4072 4724 4124
rect 4532 4059 4539 4072
rect 4717 4059 4724 4072
rect 4532 4007 4538 4059
rect 4718 4007 4724 4059
rect 4532 3994 4539 4007
rect 4717 3994 4724 4007
rect 4532 3942 4538 3994
rect 4718 3942 4724 3994
rect 4532 3929 4539 3942
rect 4717 3929 4724 3942
rect 4532 3877 4538 3929
rect 4718 3877 4724 3929
rect 4532 3864 4539 3877
rect 4717 3864 4724 3877
rect 4532 3812 4538 3864
rect 4718 3812 4724 3864
rect 4532 3799 4539 3812
rect 4717 3799 4724 3812
rect 4532 3747 4538 3799
rect 4718 3747 4724 3799
rect 4532 3734 4539 3747
rect 4717 3734 4724 3747
rect 4532 3682 4538 3734
rect 4718 3682 4724 3734
rect 4532 3669 4539 3682
rect 4717 3669 4724 3682
rect 4532 3617 4538 3669
rect 4718 3617 4724 3669
rect 4532 3604 4539 3617
rect 4717 3604 4724 3617
rect 4532 1568 4538 3604
rect 4718 1568 4724 3604
rect 4532 1562 4724 1568
rect 5028 4119 5220 4125
rect 5028 4067 5034 4119
rect 5086 4067 5098 4119
rect 5150 4067 5162 4119
rect 5214 4067 5220 4119
rect 5028 4064 5035 4067
rect 5069 4064 5107 4067
rect 5141 4064 5179 4067
rect 5213 4064 5220 4067
rect 5028 4054 5220 4064
rect 5028 4002 5034 4054
rect 5086 4002 5098 4054
rect 5150 4002 5162 4054
rect 5214 4002 5220 4054
rect 5028 3991 5035 4002
rect 5069 3991 5107 4002
rect 5141 3991 5179 4002
rect 5213 3991 5220 4002
rect 5028 3989 5220 3991
rect 5028 3937 5034 3989
rect 5086 3937 5098 3989
rect 5150 3937 5162 3989
rect 5214 3937 5220 3989
rect 5028 3924 5035 3937
rect 5069 3924 5107 3937
rect 5141 3924 5179 3937
rect 5213 3924 5220 3937
rect 5028 1568 5034 3924
rect 5214 1568 5220 3924
rect 5028 1562 5220 1568
rect 5524 4124 5716 4130
rect 5524 4072 5530 4124
rect 5582 4092 5594 4124
rect 5646 4092 5658 4124
rect 5710 4072 5716 4124
rect 5524 4059 5531 4072
rect 5709 4059 5716 4072
rect 5524 4007 5530 4059
rect 5710 4007 5716 4059
rect 5524 3994 5531 4007
rect 5709 3994 5716 4007
rect 5524 3942 5530 3994
rect 5710 3942 5716 3994
rect 5524 3929 5531 3942
rect 5709 3929 5716 3942
rect 5524 3877 5530 3929
rect 5710 3877 5716 3929
rect 5524 3864 5531 3877
rect 5709 3864 5716 3877
rect 5524 3812 5530 3864
rect 5710 3812 5716 3864
rect 5524 3799 5531 3812
rect 5709 3799 5716 3812
rect 5524 3747 5530 3799
rect 5710 3747 5716 3799
rect 5524 3734 5531 3747
rect 5709 3734 5716 3747
rect 5524 3682 5530 3734
rect 5710 3682 5716 3734
rect 5524 3669 5531 3682
rect 5709 3669 5716 3682
rect 5524 3617 5530 3669
rect 5710 3617 5716 3669
rect 5524 3604 5531 3617
rect 5709 3604 5716 3617
rect 5524 1568 5530 3604
rect 5710 1568 5716 3604
rect 5524 1562 5716 1568
rect 6020 4119 6212 4125
rect 6020 4067 6026 4119
rect 6078 4067 6090 4119
rect 6142 4067 6154 4119
rect 6206 4067 6212 4119
rect 6020 4064 6027 4067
rect 6061 4064 6099 4067
rect 6133 4064 6171 4067
rect 6205 4064 6212 4067
rect 6020 4054 6212 4064
rect 6020 4002 6026 4054
rect 6078 4002 6090 4054
rect 6142 4002 6154 4054
rect 6206 4002 6212 4054
rect 6020 3991 6027 4002
rect 6061 3991 6099 4002
rect 6133 3991 6171 4002
rect 6205 3991 6212 4002
rect 6020 3989 6212 3991
rect 6020 3937 6026 3989
rect 6078 3937 6090 3989
rect 6142 3937 6154 3989
rect 6206 3937 6212 3989
rect 6020 3924 6027 3937
rect 6061 3924 6099 3937
rect 6133 3924 6171 3937
rect 6205 3924 6212 3937
rect 6020 1568 6026 3924
rect 6206 1568 6212 3924
rect 6020 1562 6212 1568
rect 6516 4124 6708 4130
rect 6516 4072 6522 4124
rect 6574 4092 6586 4124
rect 6638 4092 6650 4124
rect 6702 4072 6708 4124
rect 6516 4059 6523 4072
rect 6701 4059 6708 4072
rect 6516 4007 6522 4059
rect 6702 4007 6708 4059
rect 6516 3994 6523 4007
rect 6701 3994 6708 4007
rect 6516 3942 6522 3994
rect 6702 3942 6708 3994
rect 6516 3929 6523 3942
rect 6701 3929 6708 3942
rect 6516 3877 6522 3929
rect 6702 3877 6708 3929
rect 6516 3864 6523 3877
rect 6701 3864 6708 3877
rect 6516 3812 6522 3864
rect 6702 3812 6708 3864
rect 6516 3799 6523 3812
rect 6701 3799 6708 3812
rect 6516 3747 6522 3799
rect 6702 3747 6708 3799
rect 6516 3734 6523 3747
rect 6701 3734 6708 3747
rect 6516 3682 6522 3734
rect 6702 3682 6708 3734
rect 6516 3669 6523 3682
rect 6701 3669 6708 3682
rect 6516 3617 6522 3669
rect 6702 3617 6708 3669
rect 6516 3604 6523 3617
rect 6701 3604 6708 3617
rect 6516 1568 6522 3604
rect 6702 1568 6708 3604
rect 6516 1562 6708 1568
rect 7012 4119 7204 4125
rect 7012 4067 7018 4119
rect 7070 4067 7082 4119
rect 7134 4067 7146 4119
rect 7198 4067 7204 4119
rect 7012 4064 7019 4067
rect 7053 4064 7091 4067
rect 7125 4064 7163 4067
rect 7197 4064 7204 4067
rect 7012 4054 7204 4064
rect 7012 4002 7018 4054
rect 7070 4002 7082 4054
rect 7134 4002 7146 4054
rect 7198 4002 7204 4054
rect 7012 3991 7019 4002
rect 7053 3991 7091 4002
rect 7125 3991 7163 4002
rect 7197 3991 7204 4002
rect 7012 3989 7204 3991
rect 7012 3937 7018 3989
rect 7070 3937 7082 3989
rect 7134 3937 7146 3989
rect 7198 3937 7204 3989
rect 7012 3924 7019 3937
rect 7053 3924 7091 3937
rect 7125 3924 7163 3937
rect 7197 3924 7204 3937
rect 7012 1568 7018 3924
rect 7198 1568 7204 3924
rect 7012 1562 7204 1568
rect 7508 4124 7700 4130
rect 7508 4072 7514 4124
rect 7566 4092 7578 4124
rect 7630 4092 7642 4124
rect 7694 4072 7700 4124
rect 7508 4059 7515 4072
rect 7693 4059 7700 4072
rect 7508 4007 7514 4059
rect 7694 4007 7700 4059
rect 7508 3994 7515 4007
rect 7693 3994 7700 4007
rect 7508 3942 7514 3994
rect 7694 3942 7700 3994
rect 7508 3929 7515 3942
rect 7693 3929 7700 3942
rect 7508 3877 7514 3929
rect 7694 3877 7700 3929
rect 7508 3864 7515 3877
rect 7693 3864 7700 3877
rect 7508 3812 7514 3864
rect 7694 3812 7700 3864
rect 7508 3799 7515 3812
rect 7693 3799 7700 3812
rect 7508 3747 7514 3799
rect 7694 3747 7700 3799
rect 7508 3734 7515 3747
rect 7693 3734 7700 3747
rect 7508 3682 7514 3734
rect 7694 3682 7700 3734
rect 7508 3669 7515 3682
rect 7693 3669 7700 3682
rect 7508 3617 7514 3669
rect 7694 3617 7700 3669
rect 7508 3604 7515 3617
rect 7693 3604 7700 3617
rect 7508 1568 7514 3604
rect 7694 1568 7700 3604
rect 7508 1562 7700 1568
rect 8004 4119 8196 4125
rect 8004 4067 8010 4119
rect 8062 4067 8074 4119
rect 8126 4067 8138 4119
rect 8190 4067 8196 4119
rect 8004 4064 8011 4067
rect 8045 4064 8083 4067
rect 8117 4064 8155 4067
rect 8189 4064 8196 4067
rect 8004 4054 8196 4064
rect 8004 4002 8010 4054
rect 8062 4002 8074 4054
rect 8126 4002 8138 4054
rect 8190 4002 8196 4054
rect 8004 3991 8011 4002
rect 8045 3991 8083 4002
rect 8117 3991 8155 4002
rect 8189 3991 8196 4002
rect 8004 3989 8196 3991
rect 8004 3937 8010 3989
rect 8062 3937 8074 3989
rect 8126 3937 8138 3989
rect 8190 3937 8196 3989
rect 8004 3924 8011 3937
rect 8045 3924 8083 3937
rect 8117 3924 8155 3937
rect 8189 3924 8196 3937
rect 8004 1568 8010 3924
rect 8190 1568 8196 3924
rect 8004 1562 8196 1568
rect 8500 4124 8692 4130
rect 8500 4072 8506 4124
rect 8558 4092 8570 4124
rect 8622 4092 8634 4124
rect 8686 4072 8692 4124
rect 8500 4059 8507 4072
rect 8685 4059 8692 4072
rect 8500 4007 8506 4059
rect 8686 4007 8692 4059
rect 8500 3994 8507 4007
rect 8685 3994 8692 4007
rect 8500 3942 8506 3994
rect 8686 3942 8692 3994
rect 8500 3929 8507 3942
rect 8685 3929 8692 3942
rect 8500 3877 8506 3929
rect 8686 3877 8692 3929
rect 8500 3864 8507 3877
rect 8685 3864 8692 3877
rect 8500 3812 8506 3864
rect 8686 3812 8692 3864
rect 8500 3799 8507 3812
rect 8685 3799 8692 3812
rect 8500 3747 8506 3799
rect 8686 3747 8692 3799
rect 8500 3734 8507 3747
rect 8685 3734 8692 3747
rect 8500 3682 8506 3734
rect 8686 3682 8692 3734
rect 8500 3669 8507 3682
rect 8685 3669 8692 3682
rect 8500 3617 8506 3669
rect 8686 3617 8692 3669
rect 8500 3604 8507 3617
rect 8685 3604 8692 3617
rect 8500 1568 8506 3604
rect 8686 1568 8692 3604
rect 8500 1562 8692 1568
rect 8996 4119 9188 4125
rect 8996 4067 9002 4119
rect 9054 4067 9066 4119
rect 9118 4067 9130 4119
rect 9182 4067 9188 4119
rect 8996 4064 9003 4067
rect 9037 4064 9075 4067
rect 9109 4064 9147 4067
rect 9181 4064 9188 4067
rect 8996 4054 9188 4064
rect 8996 4002 9002 4054
rect 9054 4002 9066 4054
rect 9118 4002 9130 4054
rect 9182 4002 9188 4054
rect 8996 3991 9003 4002
rect 9037 3991 9075 4002
rect 9109 3991 9147 4002
rect 9181 3991 9188 4002
rect 8996 3989 9188 3991
rect 8996 3937 9002 3989
rect 9054 3937 9066 3989
rect 9118 3937 9130 3989
rect 9182 3937 9188 3989
rect 8996 3924 9003 3937
rect 9037 3924 9075 3937
rect 9109 3924 9147 3937
rect 9181 3924 9188 3937
rect 8996 1568 9002 3924
rect 9182 1568 9188 3924
rect 8996 1562 9188 1568
rect 9492 4124 9684 4130
rect 9492 4072 9498 4124
rect 9550 4092 9562 4124
rect 9614 4092 9626 4124
rect 9678 4072 9684 4124
rect 9492 4059 9499 4072
rect 9677 4059 9684 4072
rect 9492 4007 9498 4059
rect 9678 4007 9684 4059
rect 9492 3994 9499 4007
rect 9677 3994 9684 4007
rect 9492 3942 9498 3994
rect 9678 3942 9684 3994
rect 9492 3929 9499 3942
rect 9677 3929 9684 3942
rect 9492 3877 9498 3929
rect 9678 3877 9684 3929
rect 9492 3864 9499 3877
rect 9677 3864 9684 3877
rect 9492 3812 9498 3864
rect 9678 3812 9684 3864
rect 9492 3799 9499 3812
rect 9677 3799 9684 3812
rect 9492 3747 9498 3799
rect 9678 3747 9684 3799
rect 9492 3734 9499 3747
rect 9677 3734 9684 3747
rect 9492 3682 9498 3734
rect 9678 3682 9684 3734
rect 9492 3669 9499 3682
rect 9677 3669 9684 3682
rect 9492 3617 9498 3669
rect 9678 3617 9684 3669
rect 9492 3604 9499 3617
rect 9677 3604 9684 3617
rect 9492 1568 9498 3604
rect 9678 1568 9684 3604
rect 9492 1562 9684 1568
rect 9988 4119 10180 4125
rect 9988 4067 9994 4119
rect 10046 4067 10058 4119
rect 10110 4067 10122 4119
rect 10174 4067 10180 4119
rect 9988 4064 9995 4067
rect 10029 4064 10067 4067
rect 10101 4064 10139 4067
rect 10173 4064 10180 4067
rect 9988 4054 10180 4064
rect 9988 4002 9994 4054
rect 10046 4002 10058 4054
rect 10110 4002 10122 4054
rect 10174 4002 10180 4054
rect 9988 3991 9995 4002
rect 10029 3991 10067 4002
rect 10101 3991 10139 4002
rect 10173 3991 10180 4002
rect 9988 3989 10180 3991
rect 9988 3937 9994 3989
rect 10046 3937 10058 3989
rect 10110 3937 10122 3989
rect 10174 3937 10180 3989
rect 9988 3924 9995 3937
rect 10029 3924 10067 3937
rect 10101 3924 10139 3937
rect 10173 3924 10180 3937
rect 9988 1568 9994 3924
rect 10174 1568 10180 3924
rect 9988 1562 10180 1568
rect 10484 4124 10676 4130
rect 10484 4072 10490 4124
rect 10542 4092 10554 4124
rect 10606 4092 10618 4124
rect 10670 4072 10676 4124
rect 10484 4059 10491 4072
rect 10669 4059 10676 4072
rect 10484 4007 10490 4059
rect 10670 4007 10676 4059
rect 10484 3994 10491 4007
rect 10669 3994 10676 4007
rect 10484 3942 10490 3994
rect 10670 3942 10676 3994
rect 10484 3929 10491 3942
rect 10669 3929 10676 3942
rect 10484 3877 10490 3929
rect 10670 3877 10676 3929
rect 10484 3864 10491 3877
rect 10669 3864 10676 3877
rect 10484 3812 10490 3864
rect 10670 3812 10676 3864
rect 10484 3799 10491 3812
rect 10669 3799 10676 3812
rect 10484 3747 10490 3799
rect 10670 3747 10676 3799
rect 10484 3734 10491 3747
rect 10669 3734 10676 3747
rect 10484 3682 10490 3734
rect 10670 3682 10676 3734
rect 10484 3669 10491 3682
rect 10669 3669 10676 3682
rect 10484 3617 10490 3669
rect 10670 3617 10676 3669
rect 10484 3604 10491 3617
rect 10669 3604 10676 3617
rect 10484 1568 10490 3604
rect 10670 1568 10676 3604
rect 10484 1562 10676 1568
rect 10980 4119 11172 4125
rect 10980 4067 10986 4119
rect 11038 4067 11050 4119
rect 11102 4067 11114 4119
rect 11166 4067 11172 4119
rect 10980 4064 10987 4067
rect 11021 4064 11059 4067
rect 11093 4064 11131 4067
rect 11165 4064 11172 4067
rect 10980 4054 11172 4064
rect 10980 4002 10986 4054
rect 11038 4002 11050 4054
rect 11102 4002 11114 4054
rect 11166 4002 11172 4054
rect 10980 3991 10987 4002
rect 11021 3991 11059 4002
rect 11093 3991 11131 4002
rect 11165 3991 11172 4002
rect 10980 3989 11172 3991
rect 10980 3937 10986 3989
rect 11038 3937 11050 3989
rect 11102 3937 11114 3989
rect 11166 3937 11172 3989
rect 10980 3924 10987 3937
rect 11021 3924 11059 3937
rect 11093 3924 11131 3937
rect 11165 3924 11172 3937
rect 10980 1568 10986 3924
rect 11166 1568 11172 3924
rect 10980 1562 11172 1568
rect 11476 4124 11668 4130
rect 11476 4072 11482 4124
rect 11534 4092 11546 4124
rect 11598 4092 11610 4124
rect 11662 4072 11668 4124
rect 11476 4059 11483 4072
rect 11661 4059 11668 4072
rect 11476 4007 11482 4059
rect 11662 4007 11668 4059
rect 11476 3994 11483 4007
rect 11661 3994 11668 4007
rect 11476 3942 11482 3994
rect 11662 3942 11668 3994
rect 11476 3929 11483 3942
rect 11661 3929 11668 3942
rect 11476 3877 11482 3929
rect 11662 3877 11668 3929
rect 11476 3864 11483 3877
rect 11661 3864 11668 3877
rect 11476 3812 11482 3864
rect 11662 3812 11668 3864
rect 11476 3799 11483 3812
rect 11661 3799 11668 3812
rect 11476 3747 11482 3799
rect 11662 3747 11668 3799
rect 11476 3734 11483 3747
rect 11661 3734 11668 3747
rect 11476 3682 11482 3734
rect 11662 3682 11668 3734
rect 11476 3669 11483 3682
rect 11661 3669 11668 3682
rect 11476 3617 11482 3669
rect 11662 3617 11668 3669
rect 11476 3604 11483 3617
rect 11661 3604 11668 3617
rect 11476 1568 11482 3604
rect 11662 1568 11668 3604
rect 11476 1562 11668 1568
rect 11972 4119 12164 4125
rect 11972 4067 11978 4119
rect 12030 4067 12042 4119
rect 12094 4067 12106 4119
rect 12158 4067 12164 4119
rect 11972 4064 11979 4067
rect 12013 4064 12051 4067
rect 12085 4064 12123 4067
rect 12157 4064 12164 4067
rect 11972 4054 12164 4064
rect 11972 4002 11978 4054
rect 12030 4002 12042 4054
rect 12094 4002 12106 4054
rect 12158 4002 12164 4054
rect 11972 3991 11979 4002
rect 12013 3991 12051 4002
rect 12085 3991 12123 4002
rect 12157 3991 12164 4002
rect 11972 3989 12164 3991
rect 11972 3937 11978 3989
rect 12030 3937 12042 3989
rect 12094 3937 12106 3989
rect 12158 3937 12164 3989
rect 11972 3924 11979 3937
rect 12013 3924 12051 3937
rect 12085 3924 12123 3937
rect 12157 3924 12164 3937
rect 11972 1568 11978 3924
rect 12158 1568 12164 3924
rect 11972 1562 12164 1568
rect 12468 4124 12660 4130
rect 12468 4072 12474 4124
rect 12526 4092 12538 4124
rect 12590 4092 12602 4124
rect 12654 4072 12660 4124
rect 12468 4059 12475 4072
rect 12653 4059 12660 4072
rect 12468 4007 12474 4059
rect 12654 4007 12660 4059
rect 12468 3994 12475 4007
rect 12653 3994 12660 4007
rect 12468 3942 12474 3994
rect 12654 3942 12660 3994
rect 12468 3929 12475 3942
rect 12653 3929 12660 3942
rect 12468 3877 12474 3929
rect 12654 3877 12660 3929
rect 12468 3864 12475 3877
rect 12653 3864 12660 3877
rect 12468 3812 12474 3864
rect 12654 3812 12660 3864
rect 12468 3799 12475 3812
rect 12653 3799 12660 3812
rect 12468 3747 12474 3799
rect 12654 3747 12660 3799
rect 12468 3734 12475 3747
rect 12653 3734 12660 3747
rect 12468 3682 12474 3734
rect 12654 3682 12660 3734
rect 12468 3669 12475 3682
rect 12653 3669 12660 3682
rect 12468 3617 12474 3669
rect 12654 3617 12660 3669
rect 12468 3604 12475 3617
rect 12653 3604 12660 3617
rect 12468 1568 12474 3604
rect 12654 1568 12660 3604
rect 12468 1562 12660 1568
rect 12964 4119 13156 4125
rect 12964 4067 12970 4119
rect 13022 4067 13034 4119
rect 13086 4067 13098 4119
rect 13150 4067 13156 4119
rect 12964 4064 12971 4067
rect 13005 4064 13043 4067
rect 13077 4064 13115 4067
rect 13149 4064 13156 4067
rect 12964 4054 13156 4064
rect 12964 4002 12970 4054
rect 13022 4002 13034 4054
rect 13086 4002 13098 4054
rect 13150 4002 13156 4054
rect 12964 3991 12971 4002
rect 13005 3991 13043 4002
rect 13077 3991 13115 4002
rect 13149 3991 13156 4002
rect 12964 3989 13156 3991
rect 12964 3937 12970 3989
rect 13022 3937 13034 3989
rect 13086 3937 13098 3989
rect 13150 3937 13156 3989
rect 12964 3924 12971 3937
rect 13005 3924 13043 3937
rect 13077 3924 13115 3937
rect 13149 3924 13156 3937
rect 12964 1568 12970 3924
rect 13150 1568 13156 3924
rect 12964 1562 13156 1568
rect 13460 4124 13652 4130
rect 13460 4072 13466 4124
rect 13518 4092 13530 4124
rect 13582 4092 13594 4124
rect 13646 4072 13652 4124
rect 13460 4059 13467 4072
rect 13645 4059 13652 4072
rect 13460 4007 13466 4059
rect 13646 4007 13652 4059
rect 13460 3994 13467 4007
rect 13645 3994 13652 4007
rect 13460 3942 13466 3994
rect 13646 3942 13652 3994
rect 13460 3929 13467 3942
rect 13645 3929 13652 3942
rect 13460 3877 13466 3929
rect 13646 3877 13652 3929
rect 13460 3864 13467 3877
rect 13645 3864 13652 3877
rect 13460 3812 13466 3864
rect 13646 3812 13652 3864
rect 13460 3799 13467 3812
rect 13645 3799 13652 3812
rect 13460 3747 13466 3799
rect 13646 3747 13652 3799
rect 13460 3734 13467 3747
rect 13645 3734 13652 3747
rect 13460 3682 13466 3734
rect 13646 3682 13652 3734
rect 13460 3669 13467 3682
rect 13645 3669 13652 3682
rect 13460 3617 13466 3669
rect 13646 3617 13652 3669
rect 13460 3604 13467 3617
rect 13645 3604 13652 3617
rect 13460 1568 13466 3604
rect 13646 1568 13652 3604
rect 13460 1562 13652 1568
rect 13957 4124 14135 4130
rect 13957 4098 13991 4124
rect 14043 4098 14083 4124
rect 13957 4064 13963 4098
rect 14069 4072 14083 4098
rect 13997 4064 14035 4072
rect 14069 4064 14135 4072
rect 13957 4060 14135 4064
rect 13957 4024 13991 4060
rect 14043 4024 14083 4060
rect 13957 3990 13963 4024
rect 14069 4008 14083 4024
rect 13997 3996 14035 4008
rect 14069 3996 14135 4008
rect 14069 3990 14083 3996
rect 13957 3950 13991 3990
rect 14043 3950 14083 3990
rect 13957 3916 13963 3950
rect 14069 3944 14083 3950
rect 13997 3932 14035 3944
rect 14069 3932 14135 3944
rect 14069 3916 14083 3932
rect 13957 3880 13991 3916
rect 14043 3880 14083 3916
rect 13957 3876 14135 3880
rect 13957 3842 13963 3876
rect 13997 3868 14035 3876
rect 14069 3868 14135 3876
rect 14069 3842 14083 3868
rect 13957 3816 13991 3842
rect 14043 3816 14083 3842
rect 13957 3804 14135 3816
rect 13957 3802 13991 3804
rect 14043 3802 14083 3804
rect 13957 3768 13963 3802
rect 14069 3768 14083 3802
rect 13957 3752 13991 3768
rect 14043 3752 14083 3768
rect 13957 3740 14135 3752
rect 13957 3728 13991 3740
rect 14043 3728 14083 3740
rect 13957 3694 13963 3728
rect 14069 3694 14083 3728
rect 13957 3688 13991 3694
rect 14043 3688 14083 3694
rect 13957 3676 14135 3688
rect 13957 3654 13991 3676
rect 14043 3654 14083 3676
rect 13957 3620 13963 3654
rect 14069 3624 14083 3654
rect 13997 3620 14035 3624
rect 14069 3620 14135 3624
rect 13957 3612 14135 3620
rect 13957 3580 13991 3612
rect 14043 3580 14083 3612
rect 13957 3546 13963 3580
rect 14069 3560 14083 3580
rect 13997 3548 14035 3560
rect 14069 3548 14135 3560
rect 14069 3546 14083 3548
rect 13957 3506 13991 3546
rect 14043 3506 14083 3546
rect 13957 3472 13963 3506
rect 14069 3496 14083 3506
rect 13997 3484 14035 3496
rect 14069 3484 14135 3496
rect 14069 3472 14083 3484
rect 13957 3432 13991 3472
rect 14043 3432 14083 3472
rect 13957 3398 13963 3432
rect 13997 3420 14035 3432
rect 14069 3420 14135 3432
rect 14069 3398 14083 3420
rect 13957 3368 13991 3398
rect 14043 3368 14083 3398
rect 13957 3358 14135 3368
rect 13957 3324 13963 3358
rect 13997 3356 14035 3358
rect 14069 3356 14135 3358
rect 14069 3324 14083 3356
rect 13957 3304 13991 3324
rect 14043 3304 14083 3324
rect 13957 3292 14135 3304
rect 13957 3284 13991 3292
rect 14043 3284 14083 3292
rect 13957 3250 13963 3284
rect 14069 3250 14083 3284
rect 13957 3240 13991 3250
rect 14043 3240 14083 3250
rect 13957 3228 14135 3240
rect 13957 3210 13991 3228
rect 14043 3210 14083 3228
rect 13957 3176 13963 3210
rect 14069 3176 14083 3210
rect 13957 3164 14135 3176
rect 13957 3136 13991 3164
rect 14043 3136 14083 3164
rect 13957 3102 13963 3136
rect 14069 3112 14083 3136
rect 13997 3102 14035 3112
rect 14069 3102 14135 3112
rect 13957 3100 14135 3102
rect 13957 3062 13991 3100
rect 14043 3062 14083 3100
rect 13957 3028 13963 3062
rect 14069 3048 14083 3062
rect 13997 3036 14035 3048
rect 14069 3036 14135 3048
rect 14069 3028 14083 3036
rect 13957 2988 13991 3028
rect 14043 2988 14083 3028
rect 13957 2954 13963 2988
rect 14069 2984 14083 2988
rect 13997 2972 14035 2984
rect 14069 2972 14135 2984
rect 14069 2954 14083 2972
rect 13957 2920 13991 2954
rect 14043 2920 14083 2954
rect 13957 2914 14135 2920
rect 13957 2880 13963 2914
rect 13997 2908 14035 2914
rect 14069 2908 14135 2914
rect 14069 2880 14083 2908
rect 13957 2856 13991 2880
rect 14043 2856 14083 2880
rect 13957 2844 14135 2856
rect 13957 2840 13991 2844
rect 14043 2840 14083 2844
rect 13957 2806 13963 2840
rect 14069 2806 14083 2840
rect 13957 2792 13991 2806
rect 14043 2792 14083 2806
rect 13957 2780 14135 2792
rect 13957 2766 13991 2780
rect 14043 2766 14083 2780
rect 13957 2732 13963 2766
rect 14069 2732 14083 2766
rect 13957 2728 13991 2732
rect 14043 2728 14083 2732
rect 13957 2716 14135 2728
rect 13957 2692 13991 2716
rect 14043 2692 14083 2716
rect 13957 2658 13963 2692
rect 14069 2664 14083 2692
rect 13997 2658 14035 2664
rect 14069 2658 14135 2664
rect 13957 2652 14135 2658
rect 13957 2618 13991 2652
rect 14043 2618 14083 2652
rect 13957 2584 13963 2618
rect 14069 2600 14083 2618
rect 13997 2588 14035 2600
rect 14069 2588 14135 2600
rect 14069 2584 14083 2588
rect 13957 2544 13991 2584
rect 14043 2544 14083 2584
rect 13957 2510 13963 2544
rect 14069 2536 14083 2544
rect 13997 2524 14035 2536
rect 14069 2524 14135 2536
rect 14069 2510 14083 2524
rect 13957 2472 13991 2510
rect 14043 2472 14083 2510
rect 13957 2470 14135 2472
rect 13957 2436 13963 2470
rect 13997 2460 14035 2470
rect 14069 2460 14135 2470
rect 14069 2436 14083 2460
rect 13957 2408 13991 2436
rect 14043 2408 14083 2436
rect 13957 2396 14135 2408
rect 13957 2362 13963 2396
rect 14069 2362 14083 2396
rect 13957 2344 13991 2362
rect 14043 2344 14083 2362
rect 13957 2332 14135 2344
rect 13957 2322 13991 2332
rect 14043 2322 14083 2332
rect 13957 2288 13963 2322
rect 14069 2288 14083 2322
rect 13957 2280 13991 2288
rect 14043 2280 14083 2288
rect 13957 2268 14135 2280
rect 13957 2248 13991 2268
rect 14043 2248 14083 2268
rect 13957 2214 13963 2248
rect 14069 2216 14083 2248
rect 13997 2214 14035 2216
rect 14069 2214 14135 2216
rect 13957 2204 14135 2214
rect 13957 2174 13991 2204
rect 14043 2174 14083 2204
rect 13957 2140 13963 2174
rect 14069 2152 14083 2174
rect 13997 2140 14035 2152
rect 14069 2140 14135 2152
rect 13957 2100 13991 2140
rect 14043 2100 14083 2140
rect 13957 2066 13963 2100
rect 14069 2088 14083 2100
rect 13997 2075 14035 2088
rect 14069 2075 14135 2088
rect 14069 2066 14083 2075
rect 13957 2026 13991 2066
rect 14043 2026 14083 2066
rect 13957 1992 13963 2026
rect 14069 2023 14083 2026
rect 13997 2010 14035 2023
rect 14069 2010 14135 2023
rect 14069 1992 14083 2010
rect 13957 1958 13991 1992
rect 14043 1958 14083 1992
rect 13957 1952 14135 1958
rect 13957 1918 13963 1952
rect 13997 1945 14035 1952
rect 14069 1945 14135 1952
rect 14069 1918 14083 1945
rect 13957 1893 13991 1918
rect 14043 1893 14083 1918
rect 13957 1880 14135 1893
rect 13957 1878 13991 1880
rect 14043 1878 14083 1880
rect 13957 1844 13963 1878
rect 14069 1844 14083 1878
rect 13957 1828 13991 1844
rect 14043 1828 14083 1844
rect 13957 1815 14135 1828
rect 13957 1804 13991 1815
rect 14043 1804 14083 1815
rect 13957 1770 13963 1804
rect 14069 1770 14083 1804
rect 13957 1763 13991 1770
rect 14043 1763 14083 1770
rect 13957 1750 14135 1763
rect 13957 1730 13991 1750
rect 14043 1730 14083 1750
rect 13957 1696 13963 1730
rect 14069 1698 14083 1730
rect 13997 1696 14035 1698
rect 14069 1696 14135 1698
rect 13957 1685 14135 1696
rect 13957 1656 13991 1685
rect 14043 1656 14083 1685
rect 13957 1622 13963 1656
rect 14069 1633 14083 1656
rect 13997 1622 14035 1633
rect 14069 1622 14135 1633
rect 13957 1620 14135 1622
rect 13957 1582 13991 1620
rect 14043 1582 14083 1620
rect 517 1530 674 1543
rect 780 1530 786 1543
rect 13957 1548 13963 1582
rect 14069 1568 14083 1582
rect 13997 1548 14035 1568
rect 14069 1548 14135 1568
rect 13957 1536 14135 1548
rect 14350 4124 14356 4140
rect 14390 4124 14428 4140
rect 14606 4124 14618 4426
rect 14402 4072 14422 4124
rect 14350 4067 14428 4072
rect 14350 4059 14356 4067
rect 14390 4059 14428 4067
rect 14606 4059 14618 4072
rect 14402 4007 14422 4059
rect 14350 3994 14428 4007
rect 14606 3994 14618 4007
rect 14402 3942 14422 3994
rect 14474 3942 14494 3960
rect 14546 3942 14566 3960
rect 14350 3929 14428 3942
rect 14462 3929 14618 3942
rect 14402 3877 14422 3929
rect 14474 3877 14494 3929
rect 14546 3877 14566 3929
rect 14350 3864 14428 3877
rect 14462 3864 14618 3877
rect 14402 3812 14422 3864
rect 14474 3812 14494 3864
rect 14546 3812 14566 3864
rect 14350 3808 14618 3812
rect 14350 3799 14428 3808
rect 14462 3799 14618 3808
rect 14402 3747 14422 3799
rect 14474 3747 14494 3799
rect 14546 3747 14566 3799
rect 14350 3741 14356 3747
rect 14390 3741 14500 3747
rect 14534 3741 14572 3747
rect 14606 3741 14618 3747
rect 14350 3736 14618 3741
rect 14350 3734 14428 3736
rect 14462 3734 14618 3736
rect 14402 3682 14422 3734
rect 14474 3682 14494 3734
rect 14546 3682 14566 3734
rect 14350 3669 14356 3682
rect 14390 3669 14500 3682
rect 14534 3669 14572 3682
rect 14606 3669 14618 3682
rect 14402 3617 14422 3669
rect 14474 3617 14494 3669
rect 14546 3617 14566 3669
rect 14350 3604 14356 3617
rect 14390 3604 14500 3617
rect 14534 3604 14572 3617
rect 14606 3604 14618 3617
rect 14402 3552 14422 3604
rect 14474 3552 14494 3604
rect 14546 3552 14566 3604
rect 14350 3540 14356 3552
rect 14390 3540 14500 3552
rect 14534 3540 14572 3552
rect 14606 3540 14618 3552
rect 14402 3488 14422 3540
rect 14474 3488 14494 3540
rect 14546 3488 14566 3540
rect 14350 3486 14428 3488
rect 14462 3486 14618 3488
rect 14350 3483 14618 3486
rect 14350 3476 14356 3483
rect 14390 3476 14500 3483
rect 14534 3476 14572 3483
rect 14606 3476 14618 3483
rect 14402 3424 14422 3476
rect 14474 3424 14494 3476
rect 14546 3424 14566 3476
rect 14350 3414 14428 3424
rect 14462 3414 14618 3424
rect 14350 3412 14618 3414
rect 14402 3360 14422 3412
rect 14474 3360 14494 3412
rect 14546 3360 14566 3412
rect 14350 3348 14428 3360
rect 14462 3348 14618 3360
rect 14402 3296 14422 3348
rect 14474 3296 14494 3348
rect 14546 3296 14566 3348
rect 14350 3284 14428 3296
rect 14462 3284 14618 3296
rect 14402 3232 14422 3284
rect 14474 3232 14494 3284
rect 14546 3232 14566 3284
rect 14350 3230 14356 3232
rect 14390 3230 14428 3232
rect 14350 3220 14428 3230
rect 14462 3230 14500 3232
rect 14534 3230 14572 3232
rect 14606 3230 14618 3232
rect 14462 3220 14618 3230
rect 14402 3168 14422 3220
rect 14474 3168 14494 3220
rect 14546 3168 14566 3220
rect 14350 3157 14356 3168
rect 14390 3160 14500 3168
rect 14390 3157 14428 3160
rect 14350 3156 14428 3157
rect 14462 3157 14500 3160
rect 14534 3157 14572 3168
rect 14606 3157 14618 3168
rect 14462 3156 14618 3157
rect 14402 3104 14422 3156
rect 14474 3104 14494 3156
rect 14546 3104 14566 3156
rect 14350 3092 14356 3104
rect 14390 3092 14500 3104
rect 14534 3092 14572 3104
rect 14606 3092 14618 3104
rect 14402 3040 14422 3092
rect 14474 3040 14494 3092
rect 14546 3040 14566 3092
rect 14350 3028 14356 3040
rect 14390 3028 14500 3040
rect 14534 3028 14572 3040
rect 14606 3028 14618 3040
rect 14402 2976 14422 3028
rect 14474 2976 14494 3028
rect 14546 2976 14566 3028
rect 14350 2972 14618 2976
rect 14350 2964 14356 2972
rect 14390 2964 14500 2972
rect 14534 2964 14572 2972
rect 14606 2964 14618 2972
rect 14402 2912 14422 2964
rect 14474 2912 14494 2964
rect 14546 2912 14566 2964
rect 14350 2910 14428 2912
rect 14462 2910 14618 2912
rect 14350 2900 14618 2910
rect 14402 2848 14422 2900
rect 14474 2848 14494 2900
rect 14546 2848 14566 2900
rect 14350 2838 14428 2848
rect 14462 2838 14618 2848
rect 14350 2836 14618 2838
rect 14402 2784 14422 2836
rect 14474 2784 14494 2836
rect 14546 2784 14566 2836
rect 14350 2772 14428 2784
rect 14462 2772 14618 2784
rect 14402 2720 14422 2772
rect 14474 2720 14494 2772
rect 14546 2720 14566 2772
rect 14350 2719 14356 2720
rect 14390 2719 14428 2720
rect 14350 2708 14428 2719
rect 14462 2719 14500 2720
rect 14534 2719 14572 2720
rect 14606 2719 14618 2720
rect 14462 2708 14618 2719
rect 14402 2656 14422 2708
rect 14474 2656 14494 2708
rect 14546 2656 14566 2708
rect 14350 2646 14356 2656
rect 14390 2646 14428 2656
rect 14350 2644 14428 2646
rect 14462 2646 14500 2656
rect 14534 2646 14572 2656
rect 14606 2646 14618 2656
rect 14462 2644 14618 2646
rect 14402 2592 14422 2644
rect 14474 2592 14494 2644
rect 14546 2592 14566 2644
rect 14350 2580 14356 2592
rect 14390 2584 14500 2592
rect 14390 2580 14428 2584
rect 14462 2580 14500 2584
rect 14534 2580 14572 2592
rect 14606 2580 14618 2592
rect 14402 2528 14422 2580
rect 14474 2528 14494 2580
rect 14546 2528 14566 2580
rect 14350 2516 14356 2528
rect 14390 2516 14500 2528
rect 14534 2516 14572 2528
rect 14606 2516 14618 2528
rect 14402 2464 14422 2516
rect 14474 2464 14494 2516
rect 14546 2464 14566 2516
rect 14350 2461 14618 2464
rect 14350 2452 14356 2461
rect 14390 2452 14500 2461
rect 14534 2452 14572 2461
rect 14606 2452 14618 2461
rect 14402 2400 14422 2452
rect 14474 2400 14494 2452
rect 14546 2400 14566 2452
rect 14350 2388 14618 2400
rect 14402 2336 14422 2388
rect 14474 2336 14494 2388
rect 14546 2336 14566 2388
rect 14350 2334 14428 2336
rect 14462 2334 14618 2336
rect 14350 2324 14618 2334
rect 14402 2272 14422 2324
rect 14474 2272 14494 2324
rect 14546 2272 14566 2324
rect 14350 2262 14428 2272
rect 14462 2262 14618 2272
rect 14350 2260 14618 2262
rect 14402 2208 14422 2260
rect 14474 2208 14494 2260
rect 14546 2208 14566 2260
rect 14350 2196 14428 2208
rect 14462 2196 14618 2208
rect 14402 2144 14422 2196
rect 14474 2144 14494 2196
rect 14546 2144 14566 2196
rect 14350 2135 14356 2144
rect 14390 2135 14428 2144
rect 14350 2132 14428 2135
rect 14462 2135 14500 2144
rect 14534 2135 14572 2144
rect 14606 2135 14618 2144
rect 14462 2132 14618 2135
rect 14402 2080 14422 2132
rect 14474 2080 14494 2132
rect 14546 2080 14566 2132
rect 14350 2068 14356 2080
rect 14390 2068 14428 2080
rect 14462 2068 14500 2080
rect 14534 2068 14572 2080
rect 14606 2068 14618 2080
rect 14402 2016 14422 2068
rect 14474 2016 14494 2068
rect 14546 2016 14566 2068
rect 14350 2004 14356 2016
rect 14390 2008 14500 2016
rect 14390 2004 14428 2008
rect 14462 2004 14500 2008
rect 14534 2004 14572 2016
rect 14606 2004 14618 2016
rect 14402 1952 14422 2004
rect 14474 1952 14494 2004
rect 14546 1952 14566 2004
rect 14350 1950 14618 1952
rect 14350 1940 14356 1950
rect 14390 1940 14500 1950
rect 14534 1940 14572 1950
rect 14606 1940 14618 1950
rect 14402 1888 14422 1940
rect 14474 1888 14494 1940
rect 14546 1888 14566 1940
rect 14350 1877 14618 1888
rect 14350 1876 14356 1877
rect 14390 1876 14500 1877
rect 14534 1876 14572 1877
rect 14606 1876 14618 1877
rect 14402 1824 14422 1876
rect 14474 1824 14494 1876
rect 14546 1824 14566 1876
rect 14350 1812 14618 1824
rect 14402 1760 14422 1812
rect 14474 1760 14494 1812
rect 14546 1760 14566 1812
rect 14350 1758 14428 1760
rect 14462 1758 14618 1760
rect 14350 1748 14618 1758
rect 14402 1696 14422 1748
rect 14474 1696 14494 1748
rect 14546 1696 14566 1748
rect 14350 1686 14428 1696
rect 14462 1686 14618 1696
rect 14350 1684 14618 1686
rect 14402 1632 14422 1684
rect 14474 1632 14494 1684
rect 14546 1632 14566 1684
rect 14350 1623 14356 1632
rect 14390 1623 14428 1632
rect 14350 1620 14428 1623
rect 14462 1624 14500 1632
rect 14534 1624 14572 1632
rect 14606 1624 14618 1632
rect 14462 1620 14618 1624
rect 14402 1568 14422 1620
rect 14474 1568 14494 1620
rect 14546 1568 14566 1620
rect 14350 1549 14356 1568
rect 14390 1549 14428 1568
rect 14350 1542 14428 1549
rect 14462 1551 14500 1568
rect 14534 1551 14572 1568
rect 14606 1551 14618 1568
rect 14462 1542 14618 1551
rect 517 1478 518 1530
rect 570 1478 590 1530
rect 642 1478 662 1530
rect 517 1465 674 1478
rect 780 1465 786 1478
rect 517 1413 518 1465
rect 570 1413 590 1465
rect 642 1413 662 1465
rect 517 1406 529 1413
rect 563 1406 601 1413
rect 635 1406 674 1413
rect 517 1400 674 1406
rect 780 1400 786 1413
rect 517 1348 518 1400
rect 570 1348 590 1400
rect 642 1348 662 1400
rect 517 1335 529 1348
rect 563 1335 601 1348
rect 635 1335 674 1348
rect 780 1335 786 1348
rect 517 1283 518 1335
rect 570 1283 590 1335
rect 642 1283 662 1335
rect 517 1270 529 1283
rect 563 1270 601 1283
rect 635 1270 674 1283
rect 780 1270 786 1283
rect 517 1218 518 1270
rect 570 1218 590 1270
rect 642 1218 662 1270
rect 14350 1512 14618 1542
rect 14350 1509 14500 1512
rect 14350 1475 14356 1509
rect 14390 1504 14500 1509
rect 14390 1475 14428 1504
rect 14350 1470 14428 1475
rect 14462 1478 14500 1504
rect 14534 1478 14572 1512
rect 14606 1478 14618 1512
rect 14462 1470 14618 1478
rect 14350 1439 14618 1470
rect 14350 1435 14500 1439
rect 14350 1401 14356 1435
rect 14390 1432 14500 1435
rect 14390 1401 14428 1432
rect 14350 1398 14428 1401
rect 14462 1405 14500 1432
rect 14534 1405 14572 1439
rect 14606 1405 14618 1439
rect 14462 1398 14618 1405
rect 14350 1366 14618 1398
rect 14350 1361 14500 1366
rect 14350 1327 14356 1361
rect 14390 1360 14500 1361
rect 14390 1327 14428 1360
rect 14350 1326 14428 1327
rect 14462 1332 14500 1360
rect 14534 1332 14572 1366
rect 14606 1332 14618 1366
rect 14462 1326 14618 1332
rect 14350 1293 14618 1326
rect 14350 1288 14500 1293
rect 14350 1287 14428 1288
rect 517 1205 529 1218
rect 563 1205 601 1218
rect 635 1205 674 1218
rect 780 1205 786 1218
rect 517 1153 518 1205
rect 570 1153 590 1205
rect 642 1153 662 1205
rect 517 1148 674 1153
rect 517 1140 529 1148
rect 563 1140 601 1148
rect 635 1140 674 1148
rect 780 1140 786 1153
rect 517 1088 518 1140
rect 570 1088 590 1140
rect 642 1088 662 1140
rect 912 1250 970 1262
rect 912 1216 924 1250
rect 958 1216 970 1250
rect 912 1178 970 1216
rect 912 1144 924 1178
rect 958 1144 970 1178
rect 912 1132 970 1144
rect 1306 1250 1436 1262
rect 1306 1144 1318 1250
rect 1424 1144 1436 1250
rect 1306 1132 1436 1144
rect 1868 1250 1998 1262
rect 1868 1144 1880 1250
rect 1986 1144 1998 1250
rect 1868 1132 1998 1144
rect 2298 1250 2428 1262
rect 2298 1144 2310 1250
rect 2416 1144 2428 1250
rect 2298 1132 2428 1144
rect 2860 1250 2990 1262
rect 2860 1144 2872 1250
rect 2978 1144 2990 1250
rect 2860 1132 2990 1144
rect 3290 1250 3420 1262
rect 3290 1144 3302 1250
rect 3408 1144 3420 1250
rect 3290 1132 3420 1144
rect 3852 1250 3982 1262
rect 3852 1144 3864 1250
rect 3970 1144 3982 1250
rect 3852 1132 3982 1144
rect 4282 1250 4412 1262
rect 4282 1144 4294 1250
rect 4400 1144 4412 1250
rect 4282 1132 4412 1144
rect 4844 1250 4974 1262
rect 4844 1144 4856 1250
rect 4962 1144 4974 1250
rect 4844 1132 4974 1144
rect 5274 1250 5404 1262
rect 5274 1144 5286 1250
rect 5392 1144 5404 1250
rect 5274 1132 5404 1144
rect 5836 1250 5966 1262
rect 5836 1144 5848 1250
rect 5954 1144 5966 1250
rect 5836 1132 5966 1144
rect 6266 1250 6396 1262
rect 6266 1144 6278 1250
rect 6384 1144 6396 1250
rect 6266 1132 6396 1144
rect 6828 1250 6958 1262
rect 6828 1144 6840 1250
rect 6946 1144 6958 1250
rect 6828 1132 6958 1144
rect 7258 1250 7388 1262
rect 7258 1144 7270 1250
rect 7376 1144 7388 1250
rect 7258 1132 7388 1144
rect 7820 1250 7950 1262
rect 7820 1144 7832 1250
rect 7938 1144 7950 1250
rect 7820 1132 7950 1144
rect 8250 1250 8380 1262
rect 8250 1144 8262 1250
rect 8368 1144 8380 1250
rect 8250 1132 8380 1144
rect 8812 1250 8942 1262
rect 8812 1144 8824 1250
rect 8930 1144 8942 1250
rect 8812 1132 8942 1144
rect 9242 1250 9372 1262
rect 9242 1144 9254 1250
rect 9360 1144 9372 1250
rect 9242 1132 9372 1144
rect 9804 1250 9934 1262
rect 9804 1144 9816 1250
rect 9922 1144 9934 1250
rect 9804 1132 9934 1144
rect 10234 1250 10364 1262
rect 10234 1144 10246 1250
rect 10352 1144 10364 1250
rect 10234 1132 10364 1144
rect 10796 1250 10926 1262
rect 10796 1144 10808 1250
rect 10914 1144 10926 1250
rect 10796 1132 10926 1144
rect 11226 1250 11356 1262
rect 11226 1144 11238 1250
rect 11344 1144 11356 1250
rect 11226 1132 11356 1144
rect 11788 1250 11918 1262
rect 11788 1144 11800 1250
rect 11906 1144 11918 1250
rect 11788 1132 11918 1144
rect 12218 1250 12348 1262
rect 12218 1144 12230 1250
rect 12336 1144 12348 1250
rect 12218 1132 12348 1144
rect 12780 1250 12910 1262
rect 12780 1144 12792 1250
rect 12898 1144 12910 1250
rect 12780 1132 12910 1144
rect 13210 1250 13340 1262
rect 13210 1144 13222 1250
rect 13328 1144 13340 1250
rect 13210 1132 13340 1144
rect 13772 1250 13902 1262
rect 13772 1144 13784 1250
rect 13890 1144 13902 1250
rect 13772 1132 13902 1144
rect 14130 1250 14260 1262
rect 14130 1144 14142 1250
rect 14248 1144 14260 1250
rect 14130 1132 14260 1144
rect 14350 1253 14356 1287
rect 14390 1254 14428 1287
rect 14462 1259 14500 1288
rect 14534 1259 14572 1293
rect 14606 1259 14618 1293
rect 14462 1254 14618 1259
rect 14390 1253 14618 1254
rect 14350 1220 14618 1253
rect 14350 1216 14500 1220
rect 14350 1213 14428 1216
rect 14350 1179 14356 1213
rect 14390 1182 14428 1213
rect 14462 1186 14500 1216
rect 14534 1186 14572 1220
rect 14606 1186 14618 1220
rect 14462 1182 14618 1186
rect 14390 1179 14618 1182
rect 14350 1147 14618 1179
rect 14350 1144 14500 1147
rect 14350 1139 14428 1144
rect 517 1075 674 1088
rect 780 1075 786 1088
rect 517 1023 518 1075
rect 570 1023 590 1075
rect 642 1023 662 1075
rect 14350 1105 14356 1139
rect 14390 1110 14428 1139
rect 14462 1113 14500 1144
rect 14534 1113 14572 1147
rect 14606 1113 14618 1147
rect 14462 1110 14618 1113
rect 14390 1105 14618 1110
rect 14350 1074 14618 1105
rect 14350 1072 14500 1074
rect 14350 1065 14428 1072
rect 14350 1031 14356 1065
rect 14390 1038 14428 1065
rect 14462 1040 14500 1072
rect 14534 1040 14572 1074
rect 14606 1040 14618 1074
rect 14462 1038 14618 1040
rect 14390 1031 14618 1038
tri 14349 1024 14350 1025 se
rect 14350 1024 14618 1031
rect 517 1010 674 1023
rect 780 1010 786 1023
rect 517 958 518 1010
rect 570 958 590 1010
rect 642 958 662 1010
tri 786 1001 809 1024 sw
tri 14326 1001 14349 1024 se
rect 14349 1001 14618 1024
rect 786 1000 809 1001
tri 809 1000 810 1001 sw
tri 14325 1000 14326 1001 se
rect 14326 1000 14500 1001
rect 786 991 810 1000
tri 810 991 819 1000 sw
tri 14316 991 14325 1000 se
rect 14325 991 14428 1000
rect 786 958 819 991
rect 517 945 674 958
rect 780 957 819 958
tri 819 957 853 991 sw
tri 14282 957 14316 991 se
rect 14316 957 14356 991
rect 14390 966 14428 991
rect 14462 967 14500 1000
rect 14534 967 14572 1001
rect 14606 967 14618 1001
rect 14462 966 14618 967
rect 14390 957 14618 966
rect 780 945 853 957
rect 517 893 518 945
rect 570 893 590 945
rect 642 893 662 945
rect 714 893 734 894
rect 786 928 853 945
tri 853 928 882 957 sw
tri 14253 928 14282 957 se
rect 14282 928 14618 957
rect 786 917 882 928
tri 882 917 893 928 sw
tri 14242 917 14253 928 se
rect 14253 917 14428 928
rect 786 893 893 917
rect 517 883 746 893
rect 780 883 893 893
tri 893 883 927 917 sw
tri 14208 883 14242 917 se
rect 14242 883 14356 917
rect 14390 894 14428 917
rect 14462 894 14500 928
rect 14534 894 14572 928
rect 14606 894 14618 928
rect 14390 883 14618 894
rect 231 829 269 863
rect 303 845 329 863
tri 329 845 366 882 sw
rect 517 880 927 883
rect 303 829 366 845
rect 231 820 366 829
tri 366 820 391 845 sw
rect 517 828 518 880
rect 570 828 590 880
rect 642 828 662 880
rect 714 828 734 880
rect 786 872 927 880
tri 927 872 938 883 sw
tri 14197 872 14208 883 se
rect 14208 872 14618 883
rect 786 845 938 872
tri 938 845 965 872 sw
tri 14196 871 14197 872 se
rect 14197 871 14618 872
tri 14184 859 14196 871 se
rect 14196 859 14618 871
rect 14807 1468 14835 4618
rect 14807 1429 14907 1468
rect 14807 1395 14835 1429
rect 14869 1395 14907 1429
rect 14807 1356 14907 1395
rect 14807 1322 14835 1356
rect 14869 1322 14907 1356
rect 14807 1283 14907 1322
rect 14807 1249 14835 1283
rect 14869 1249 14907 1283
rect 14807 1210 14907 1249
rect 14807 1176 14835 1210
rect 14869 1176 14907 1210
rect 14807 1137 14907 1176
rect 14807 1103 14835 1137
rect 14869 1103 14907 1137
rect 14807 1064 14907 1103
rect 14807 1030 14835 1064
rect 14869 1030 14907 1064
rect 14807 991 14907 1030
rect 14807 957 14835 991
rect 14869 957 14907 991
rect 14807 918 14907 957
rect 14807 884 14835 918
rect 14869 884 14907 918
tri 14170 845 14184 859 se
rect 14184 845 14618 859
tri 14793 845 14807 859 se
rect 14807 845 14907 884
rect 786 832 965 845
tri 965 832 978 845 sw
tri 14157 832 14170 845 se
rect 14170 832 14618 845
rect 786 828 14618 832
rect 517 820 14618 828
rect 231 818 391 820
tri 391 818 393 820 sw
rect 517 818 709 820
rect 231 789 393 818
rect 231 755 269 789
rect 303 786 393 789
tri 393 786 425 818 sw
tri 517 786 549 818 ne
rect 549 786 709 818
rect 743 786 782 820
rect 816 786 855 820
rect 889 786 928 820
rect 303 755 425 786
rect 231 748 425 755
tri 425 748 463 786 sw
tri 549 748 587 786 ne
rect 587 748 928 786
rect 231 715 463 748
rect 231 681 269 715
rect 303 714 463 715
tri 463 714 497 748 sw
tri 587 714 621 748 ne
rect 621 714 709 748
rect 743 714 782 748
rect 816 714 855 748
rect 889 714 928 748
rect 14426 818 14618 820
rect 14426 811 14611 818
tri 14611 811 14618 818 nw
tri 14759 811 14793 845 se
rect 14793 811 14835 845
rect 14869 811 14907 845
rect 14426 772 14572 811
tri 14572 772 14611 811 nw
tri 14720 772 14759 811 se
rect 14759 772 14907 811
rect 14426 738 14538 772
tri 14538 738 14572 772 nw
tri 14686 738 14720 772 se
rect 14720 738 14835 772
rect 14869 738 14907 772
rect 14426 714 14502 738
rect 303 702 497 714
tri 497 702 509 714 sw
tri 621 702 633 714 ne
rect 633 702 14502 714
tri 14502 702 14538 738 nw
tri 14650 702 14686 738 se
rect 14686 702 14907 738
rect 303 699 509 702
tri 509 699 512 702 sw
tri 14647 699 14650 702 se
rect 14650 699 14907 702
rect 303 681 512 699
rect 231 665 512 681
tri 512 665 546 699 sw
tri 14613 665 14647 699 se
rect 14647 665 14835 699
rect 14869 665 14907 699
rect 231 641 546 665
rect 231 607 269 641
rect 303 626 546 641
tri 546 626 585 665 sw
tri 14574 626 14613 665 se
rect 14613 626 14907 665
rect 303 607 585 626
rect 231 592 585 607
tri 585 592 619 626 sw
tri 14540 592 14574 626 se
rect 14574 592 14835 626
rect 14869 592 14907 626
rect 231 567 619 592
rect 231 533 269 567
rect 303 553 619 567
tri 619 553 658 592 sw
tri 14501 553 14540 592 se
rect 14540 553 14907 592
rect 303 533 658 553
rect 231 519 658 533
tri 658 519 692 553 sw
tri 14467 519 14501 553 se
rect 14501 519 14835 553
rect 14869 519 14907 553
rect 231 505 692 519
tri 692 505 706 519 sw
tri 14453 505 14467 519 se
rect 14467 505 14907 519
rect 231 497 706 505
rect 231 463 343 497
rect 377 463 419 497
rect 453 463 495 497
rect 529 463 571 497
rect 605 463 648 497
rect 682 481 706 497
tri 706 481 730 505 sw
tri 14435 487 14453 505 se
rect 14453 487 14907 505
tri 14429 481 14435 487 se
rect 14435 481 14907 487
rect 682 463 730 481
rect 231 447 730 463
tri 730 447 764 481 sw
tri 14395 447 14429 481 se
rect 14429 447 14468 481
rect 14502 447 14542 481
rect 14576 447 14616 481
rect 14650 447 14689 481
rect 14723 447 14762 481
rect 14796 447 14907 481
rect 231 420 764 447
tri 764 420 791 447 sw
tri 14389 441 14395 447 se
rect 14395 441 14907 447
tri 14368 420 14389 441 se
rect 14389 420 14907 441
rect 15013 420 15097 5062
rect 231 402 791 420
tri 791 402 809 420 sw
tri 14350 402 14368 420 se
rect 14368 402 15097 420
rect 231 375 15097 402
rect 231 341 361 375
rect 395 341 434 375
rect 468 341 507 375
rect 541 341 580 375
rect 614 341 653 375
rect 687 341 726 375
rect 760 341 799 375
rect 833 341 872 375
rect 906 341 945 375
rect 979 341 1018 375
rect 1052 341 1091 375
rect 1125 341 1164 375
rect 1198 341 1237 375
rect 1271 341 1310 375
rect 1344 341 1383 375
rect 1417 341 1456 375
rect 1490 341 1529 375
rect 1563 341 1602 375
rect 1636 341 1675 375
rect 1709 341 1748 375
rect 1782 341 1821 375
rect 1855 341 1894 375
rect 1928 341 1967 375
rect 2001 341 2040 375
rect 2074 341 2113 375
rect 2147 341 2186 375
rect 2220 341 2259 375
rect 2293 341 2332 375
rect 2366 341 2405 375
rect 2439 341 2478 375
rect 2512 341 2551 375
rect 2585 341 2624 375
rect 2658 341 2697 375
rect 2731 341 2770 375
rect 2804 341 2843 375
rect 2877 341 2916 375
rect 2950 341 2989 375
rect 3023 341 3062 375
rect 3096 341 3135 375
rect 3169 341 3208 375
rect 3242 341 3281 375
rect 3315 341 3354 375
rect 3388 341 3427 375
rect 3461 341 3500 375
rect 3534 341 3573 375
rect 3607 341 3646 375
rect 3680 341 3719 375
rect 3753 341 3792 375
rect 3826 341 3865 375
rect 3899 341 3938 375
rect 3972 341 4011 375
rect 4045 341 4084 375
rect 4118 341 4157 375
rect 4191 341 4229 375
rect 4263 341 4301 375
rect 4335 341 4373 375
rect 4407 341 4445 375
rect 4479 341 4517 375
rect 4551 341 4589 375
rect 4623 341 4661 375
rect 4695 341 4733 375
rect 4767 341 4805 375
rect 4839 341 4877 375
rect 4911 341 4949 375
rect 4983 341 5021 375
rect 5055 341 5093 375
rect 5127 341 5165 375
rect 5199 341 5237 375
rect 5271 341 5309 375
rect 5343 341 5381 375
rect 5415 341 5453 375
rect 5487 341 5525 375
rect 5559 341 5597 375
rect 5631 341 5669 375
rect 5703 341 5741 375
rect 5775 341 5813 375
rect 5847 341 5885 375
rect 5919 341 5957 375
rect 5991 341 6029 375
rect 6063 341 6101 375
rect 6135 341 6173 375
rect 6207 341 6245 375
rect 6279 341 6317 375
rect 6351 341 6389 375
rect 6423 341 6461 375
rect 6495 341 6533 375
rect 6567 341 6605 375
rect 6639 341 6677 375
rect 6711 341 6749 375
rect 6783 341 6821 375
rect 6855 341 6893 375
rect 6927 341 6965 375
rect 6999 341 7037 375
rect 7071 341 7109 375
rect 7143 341 7181 375
rect 7215 341 7253 375
rect 7287 341 7325 375
rect 7359 341 7397 375
rect 7431 341 7469 375
rect 7503 341 7541 375
rect 7575 341 7613 375
rect 7647 341 7685 375
rect 7719 341 7757 375
rect 7791 341 7829 375
rect 7863 341 7901 375
rect 7935 341 7973 375
rect 8007 341 8045 375
rect 8079 341 8117 375
rect 8151 341 8189 375
rect 8223 341 8261 375
rect 8295 341 8333 375
rect 8367 341 8405 375
rect 8439 341 8477 375
rect 8511 341 8549 375
rect 8583 341 8621 375
rect 8655 341 8693 375
rect 8727 341 8765 375
rect 8799 341 8837 375
rect 8871 341 8909 375
rect 8943 341 8981 375
rect 9015 341 9053 375
rect 9087 341 9125 375
rect 9159 341 9197 375
rect 9231 341 9269 375
rect 9303 341 9341 375
rect 9375 341 9413 375
rect 9447 341 9485 375
rect 9519 341 9557 375
rect 9591 341 9629 375
rect 9663 341 9701 375
rect 9735 341 9773 375
rect 9807 341 9845 375
rect 9879 341 9917 375
rect 9951 341 9989 375
rect 10023 341 10061 375
rect 10095 341 10133 375
rect 10167 341 10205 375
rect 10239 341 10277 375
rect 10311 341 10349 375
rect 10383 341 10421 375
rect 10455 341 10493 375
rect 10527 341 10565 375
rect 10599 341 10637 375
rect 10671 341 10709 375
rect 10743 341 10781 375
rect 10815 341 10853 375
rect 10887 341 10925 375
rect 10959 341 10997 375
rect 11031 341 11069 375
rect 11103 341 11141 375
rect 11175 341 11213 375
rect 11247 341 11285 375
rect 11319 341 11357 375
rect 11391 341 11429 375
rect 11463 341 11501 375
rect 11535 341 11573 375
rect 11607 341 11645 375
rect 11679 341 11717 375
rect 11751 341 11789 375
rect 11823 341 11861 375
rect 11895 341 11933 375
rect 11967 341 12005 375
rect 12039 341 12077 375
rect 12111 341 12149 375
rect 12183 341 12221 375
rect 12255 341 12293 375
rect 12327 341 12365 375
rect 12399 341 12437 375
rect 12471 341 12509 375
rect 12543 341 12581 375
rect 12615 341 12653 375
rect 12687 341 12725 375
rect 12759 341 12797 375
rect 12831 341 12869 375
rect 12903 341 12941 375
rect 12975 341 13013 375
rect 13047 341 13085 375
rect 13119 341 13157 375
rect 13191 341 13229 375
rect 13263 341 13301 375
rect 13335 341 13373 375
rect 13407 341 13445 375
rect 13479 341 13517 375
rect 13551 341 13589 375
rect 13623 341 13661 375
rect 13695 341 13733 375
rect 13767 341 13805 375
rect 13839 341 13877 375
rect 13911 341 13949 375
rect 13983 341 14021 375
rect 14055 341 14093 375
rect 14127 341 14165 375
rect 14199 341 14237 375
rect 14271 341 14309 375
rect 14343 341 14381 375
rect 14415 341 14453 375
rect 14487 341 14525 375
rect 14559 341 14597 375
rect 14631 341 14669 375
rect 14703 341 14741 375
rect 14775 341 15097 375
rect 231 331 15097 341
rect 39 314 15097 331
<< via1 >>
rect 518 4426 570 4456
rect 518 4404 529 4426
rect 529 4404 563 4426
rect 563 4404 570 4426
rect 590 4426 642 4456
rect 590 4404 601 4426
rect 601 4404 635 4426
rect 635 4404 642 4426
rect 662 4404 674 4456
rect 674 4445 708 4456
rect 708 4445 714 4456
rect 734 4445 786 4456
rect 674 4404 714 4445
rect 734 4404 780 4445
rect 780 4404 786 4445
rect 518 4351 570 4390
rect 518 4338 529 4351
rect 529 4338 563 4351
rect 563 4338 570 4351
rect 590 4351 642 4390
rect 590 4338 601 4351
rect 601 4338 635 4351
rect 635 4338 642 4351
rect 662 4338 674 4390
rect 674 4338 714 4390
rect 734 4338 780 4390
rect 780 4338 786 4390
rect 518 4317 529 4325
rect 529 4317 563 4325
rect 563 4317 570 4325
rect 518 4276 570 4317
rect 518 4273 529 4276
rect 529 4273 563 4276
rect 563 4273 570 4276
rect 590 4317 601 4325
rect 601 4317 635 4325
rect 635 4317 642 4325
rect 590 4276 642 4317
rect 590 4273 601 4276
rect 601 4273 635 4276
rect 635 4273 642 4276
rect 662 4273 674 4325
rect 674 4273 714 4325
rect 734 4273 780 4325
rect 780 4273 786 4325
rect 518 4242 529 4260
rect 529 4242 563 4260
rect 563 4242 570 4260
rect 518 4208 570 4242
rect 590 4242 601 4260
rect 601 4242 635 4260
rect 635 4242 642 4260
rect 590 4208 642 4242
rect 662 4208 674 4260
rect 674 4208 714 4260
rect 734 4208 780 4260
rect 780 4208 786 4260
rect 518 4167 529 4195
rect 529 4167 563 4195
rect 563 4167 570 4195
rect 518 4143 570 4167
rect 590 4167 601 4195
rect 601 4167 635 4195
rect 635 4167 642 4195
rect 590 4143 642 4167
rect 662 4143 674 4195
rect 674 4143 714 4195
rect 734 4143 780 4195
rect 780 4143 786 4195
rect 518 4126 570 4130
rect 518 4092 529 4126
rect 529 4092 563 4126
rect 563 4092 570 4126
rect 518 4078 570 4092
rect 590 4126 642 4130
rect 590 4092 601 4126
rect 601 4092 635 4126
rect 635 4092 642 4126
rect 590 4078 642 4092
rect 662 4078 674 4130
rect 674 4078 714 4130
rect 734 4078 780 4130
rect 780 4078 786 4130
rect 518 4052 570 4065
rect 518 4018 529 4052
rect 529 4018 563 4052
rect 563 4018 570 4052
rect 518 4013 570 4018
rect 590 4052 642 4065
rect 590 4018 601 4052
rect 601 4018 635 4052
rect 635 4018 642 4052
rect 590 4013 642 4018
rect 662 4013 674 4065
rect 674 4013 714 4065
rect 734 4013 780 4065
rect 780 4013 786 4065
rect 518 3978 570 4000
rect 518 3948 529 3978
rect 529 3948 563 3978
rect 563 3948 570 3978
rect 590 3978 642 4000
rect 590 3948 601 3978
rect 601 3948 635 3978
rect 635 3948 642 3978
rect 662 3948 674 4000
rect 674 3948 714 4000
rect 734 3948 780 4000
rect 780 3948 786 4000
rect 518 3904 570 3935
rect 518 3883 529 3904
rect 529 3883 563 3904
rect 563 3883 570 3904
rect 590 3904 642 3935
rect 590 3883 601 3904
rect 601 3883 635 3904
rect 635 3883 642 3904
rect 662 3883 674 3935
rect 674 3883 714 3935
rect 734 3883 780 3935
rect 780 3883 786 3935
rect 518 3818 570 3870
rect 590 3818 642 3870
rect 662 3818 674 3870
rect 674 3818 714 3870
rect 734 3818 780 3870
rect 780 3818 786 3870
rect 518 3794 570 3805
rect 518 3760 529 3794
rect 529 3760 563 3794
rect 563 3760 570 3794
rect 518 3753 570 3760
rect 590 3794 642 3805
rect 590 3760 601 3794
rect 601 3760 635 3794
rect 635 3760 642 3794
rect 590 3753 642 3760
rect 662 3753 674 3805
rect 674 3753 714 3805
rect 734 3753 780 3805
rect 780 3753 786 3805
rect 518 3720 570 3740
rect 518 3688 529 3720
rect 529 3688 563 3720
rect 563 3688 570 3720
rect 590 3720 642 3740
rect 590 3688 601 3720
rect 601 3688 635 3720
rect 635 3688 642 3720
rect 662 3688 674 3740
rect 674 3688 714 3740
rect 734 3688 780 3740
rect 780 3688 786 3740
rect 518 3646 570 3675
rect 518 3623 529 3646
rect 529 3623 563 3646
rect 563 3623 570 3646
rect 590 3646 642 3675
rect 590 3623 601 3646
rect 601 3623 635 3646
rect 635 3623 642 3646
rect 662 3623 674 3675
rect 674 3623 714 3675
rect 734 3623 780 3675
rect 780 3623 786 3675
rect 518 3572 570 3610
rect 518 3558 529 3572
rect 529 3558 563 3572
rect 563 3558 570 3572
rect 590 3572 642 3610
rect 590 3558 601 3572
rect 601 3558 635 3572
rect 635 3558 642 3572
rect 662 3558 674 3610
rect 674 3558 714 3610
rect 734 3558 780 3610
rect 780 3558 786 3610
rect 518 3538 529 3545
rect 529 3538 563 3545
rect 563 3538 570 3545
rect 518 3498 570 3538
rect 518 3493 529 3498
rect 529 3493 563 3498
rect 563 3493 570 3498
rect 590 3538 601 3545
rect 601 3538 635 3545
rect 635 3538 642 3545
rect 590 3498 642 3538
rect 590 3493 601 3498
rect 601 3493 635 3498
rect 635 3493 642 3498
rect 662 3493 674 3545
rect 674 3493 714 3545
rect 734 3493 780 3545
rect 780 3493 786 3545
rect 518 3464 529 3480
rect 529 3464 563 3480
rect 563 3464 570 3480
rect 518 3428 570 3464
rect 590 3464 601 3480
rect 601 3464 635 3480
rect 635 3464 642 3480
rect 590 3428 642 3464
rect 662 3428 674 3480
rect 674 3428 714 3480
rect 734 3428 780 3480
rect 780 3428 786 3480
rect 518 3390 529 3415
rect 529 3390 563 3415
rect 563 3390 570 3415
rect 518 3363 570 3390
rect 590 3390 601 3415
rect 601 3390 635 3415
rect 635 3390 642 3415
rect 590 3363 642 3390
rect 662 3363 674 3415
rect 674 3363 714 3415
rect 734 3363 780 3415
rect 780 3363 786 3415
rect 518 3316 529 3350
rect 529 3316 563 3350
rect 563 3316 570 3350
rect 518 3298 570 3316
rect 590 3316 601 3350
rect 601 3316 635 3350
rect 635 3316 642 3350
rect 590 3298 642 3316
rect 662 3298 674 3350
rect 674 3298 714 3350
rect 734 3298 780 3350
rect 780 3298 786 3350
rect 518 3276 570 3285
rect 518 3242 529 3276
rect 529 3242 563 3276
rect 563 3242 570 3276
rect 518 3233 570 3242
rect 590 3276 642 3285
rect 590 3242 601 3276
rect 601 3242 635 3276
rect 635 3242 642 3276
rect 590 3233 642 3242
rect 662 3233 674 3285
rect 674 3233 714 3285
rect 734 3233 780 3285
rect 780 3233 786 3285
rect 518 3202 570 3220
rect 518 3168 529 3202
rect 529 3168 563 3202
rect 563 3168 570 3202
rect 590 3202 642 3220
rect 590 3168 601 3202
rect 601 3168 635 3202
rect 635 3168 642 3202
rect 662 3168 674 3220
rect 674 3168 714 3220
rect 734 3168 780 3220
rect 780 3168 786 3220
rect 518 3128 570 3155
rect 518 3103 529 3128
rect 529 3103 563 3128
rect 563 3103 570 3128
rect 590 3128 642 3155
rect 590 3103 601 3128
rect 601 3103 635 3128
rect 635 3103 642 3128
rect 662 3103 674 3155
rect 674 3103 714 3155
rect 734 3103 780 3155
rect 780 3103 786 3155
rect 518 3054 570 3090
rect 518 3038 529 3054
rect 529 3038 563 3054
rect 563 3038 570 3054
rect 590 3054 642 3090
rect 590 3038 601 3054
rect 601 3038 635 3054
rect 635 3038 642 3054
rect 662 3038 674 3090
rect 674 3038 714 3090
rect 734 3038 780 3090
rect 780 3038 786 3090
rect 518 3020 529 3025
rect 529 3020 563 3025
rect 563 3020 570 3025
rect 518 2980 570 3020
rect 518 2973 529 2980
rect 529 2973 563 2980
rect 563 2973 570 2980
rect 590 3020 601 3025
rect 601 3020 635 3025
rect 635 3020 642 3025
rect 590 2980 642 3020
rect 590 2973 601 2980
rect 601 2973 635 2980
rect 635 2973 642 2980
rect 662 2973 674 3025
rect 674 2973 714 3025
rect 734 2973 780 3025
rect 780 2973 786 3025
rect 518 2946 529 2960
rect 529 2946 563 2960
rect 563 2946 570 2960
rect 518 2908 570 2946
rect 590 2946 601 2960
rect 601 2946 635 2960
rect 635 2946 642 2960
rect 590 2908 642 2946
rect 662 2908 674 2960
rect 674 2908 714 2960
rect 734 2908 780 2960
rect 780 2908 786 2960
rect 518 2872 529 2895
rect 529 2872 563 2895
rect 563 2872 570 2895
rect 518 2843 570 2872
rect 590 2872 601 2895
rect 601 2872 635 2895
rect 635 2872 642 2895
rect 590 2843 642 2872
rect 662 2843 674 2895
rect 674 2843 714 2895
rect 734 2843 780 2895
rect 780 2843 786 2895
rect 518 2798 529 2830
rect 529 2798 563 2830
rect 563 2798 570 2830
rect 518 2778 570 2798
rect 590 2798 601 2830
rect 601 2798 635 2830
rect 635 2798 642 2830
rect 590 2778 642 2798
rect 662 2778 674 2830
rect 674 2778 714 2830
rect 734 2778 780 2830
rect 780 2778 786 2830
rect 518 2758 570 2765
rect 518 2724 529 2758
rect 529 2724 563 2758
rect 563 2724 570 2758
rect 518 2713 570 2724
rect 590 2758 642 2765
rect 590 2724 601 2758
rect 601 2724 635 2758
rect 635 2724 642 2758
rect 590 2713 642 2724
rect 662 2713 674 2765
rect 674 2713 714 2765
rect 734 2713 780 2765
rect 780 2713 786 2765
rect 518 2684 570 2700
rect 518 2650 529 2684
rect 529 2650 563 2684
rect 563 2650 570 2684
rect 518 2648 570 2650
rect 590 2684 642 2700
rect 590 2650 601 2684
rect 601 2650 635 2684
rect 635 2650 642 2684
rect 590 2648 642 2650
rect 662 2648 674 2700
rect 674 2648 714 2700
rect 734 2648 780 2700
rect 780 2648 786 2700
rect 518 2610 570 2635
rect 518 2583 529 2610
rect 529 2583 563 2610
rect 563 2583 570 2610
rect 590 2610 642 2635
rect 590 2583 601 2610
rect 601 2583 635 2610
rect 635 2583 642 2610
rect 662 2583 674 2635
rect 674 2583 714 2635
rect 734 2583 780 2635
rect 780 2583 786 2635
rect 518 2536 570 2570
rect 518 2518 529 2536
rect 529 2518 563 2536
rect 563 2518 570 2536
rect 590 2536 642 2570
rect 590 2518 601 2536
rect 601 2518 635 2536
rect 635 2518 642 2536
rect 662 2518 674 2570
rect 674 2518 714 2570
rect 734 2518 780 2570
rect 780 2518 786 2570
rect 518 2502 529 2505
rect 529 2502 563 2505
rect 563 2502 570 2505
rect 518 2462 570 2502
rect 518 2453 529 2462
rect 529 2453 563 2462
rect 563 2453 570 2462
rect 590 2502 601 2505
rect 601 2502 635 2505
rect 635 2502 642 2505
rect 590 2462 642 2502
rect 590 2453 601 2462
rect 601 2453 635 2462
rect 635 2453 642 2462
rect 662 2453 674 2505
rect 674 2453 714 2505
rect 734 2453 780 2505
rect 780 2453 786 2505
rect 518 2428 529 2440
rect 529 2428 563 2440
rect 563 2428 570 2440
rect 518 2389 570 2428
rect 518 2388 529 2389
rect 529 2388 563 2389
rect 563 2388 570 2389
rect 590 2428 601 2440
rect 601 2428 635 2440
rect 635 2428 642 2440
rect 590 2389 642 2428
rect 590 2388 601 2389
rect 601 2388 635 2389
rect 635 2388 642 2389
rect 662 2388 674 2440
rect 674 2388 714 2440
rect 734 2388 780 2440
rect 780 2388 786 2440
rect 518 2355 529 2375
rect 529 2355 563 2375
rect 563 2355 570 2375
rect 518 2323 570 2355
rect 590 2355 601 2375
rect 601 2355 635 2375
rect 635 2355 642 2375
rect 590 2323 642 2355
rect 662 2323 674 2375
rect 674 2323 714 2375
rect 734 2323 780 2375
rect 780 2323 786 2375
rect 518 2282 529 2310
rect 529 2282 563 2310
rect 563 2282 570 2310
rect 518 2258 570 2282
rect 590 2282 601 2310
rect 601 2282 635 2310
rect 635 2282 642 2310
rect 590 2258 642 2282
rect 662 2258 674 2310
rect 674 2258 714 2310
rect 734 2258 780 2310
rect 780 2258 786 2310
rect 518 2243 570 2245
rect 518 2209 529 2243
rect 529 2209 563 2243
rect 563 2209 570 2243
rect 518 2193 570 2209
rect 590 2243 642 2245
rect 590 2209 601 2243
rect 601 2209 635 2243
rect 635 2209 642 2243
rect 590 2193 642 2209
rect 662 2193 674 2245
rect 674 2193 714 2245
rect 734 2193 780 2245
rect 780 2193 786 2245
rect 518 2170 570 2180
rect 518 2136 529 2170
rect 529 2136 563 2170
rect 563 2136 570 2170
rect 518 2128 570 2136
rect 590 2170 642 2180
rect 590 2136 601 2170
rect 601 2136 635 2170
rect 635 2136 642 2170
rect 590 2128 642 2136
rect 662 2128 674 2180
rect 674 2128 714 2180
rect 734 2128 780 2180
rect 780 2128 786 2180
rect 518 2097 570 2115
rect 518 2063 529 2097
rect 529 2063 563 2097
rect 563 2063 570 2097
rect 590 2097 642 2115
rect 590 2063 601 2097
rect 601 2063 635 2097
rect 635 2063 642 2097
rect 662 2063 674 2115
rect 674 2063 714 2115
rect 734 2063 780 2115
rect 780 2063 786 2115
rect 518 2024 570 2050
rect 518 1998 529 2024
rect 529 1998 563 2024
rect 563 1998 570 2024
rect 590 2024 642 2050
rect 590 1998 601 2024
rect 601 1998 635 2024
rect 635 1998 642 2024
rect 662 1998 674 2050
rect 674 1998 714 2050
rect 734 1998 780 2050
rect 780 1998 786 2050
rect 518 1951 570 1985
rect 518 1933 529 1951
rect 529 1933 563 1951
rect 563 1933 570 1951
rect 590 1951 642 1985
rect 590 1933 601 1951
rect 601 1933 635 1951
rect 635 1933 642 1951
rect 662 1933 674 1985
rect 674 1933 714 1985
rect 734 1933 780 1985
rect 780 1933 786 1985
rect 518 1917 529 1920
rect 529 1917 563 1920
rect 563 1917 570 1920
rect 518 1878 570 1917
rect 518 1868 529 1878
rect 529 1868 563 1878
rect 563 1868 570 1878
rect 590 1917 601 1920
rect 601 1917 635 1920
rect 635 1917 642 1920
rect 590 1878 642 1917
rect 590 1868 601 1878
rect 601 1868 635 1878
rect 635 1868 642 1878
rect 662 1868 674 1920
rect 674 1868 714 1920
rect 734 1868 780 1920
rect 780 1868 786 1920
rect 518 1844 529 1855
rect 529 1844 563 1855
rect 563 1844 570 1855
rect 518 1805 570 1844
rect 518 1803 529 1805
rect 529 1803 563 1805
rect 563 1803 570 1805
rect 590 1844 601 1855
rect 601 1844 635 1855
rect 635 1844 642 1855
rect 590 1805 642 1844
rect 590 1803 601 1805
rect 601 1803 635 1805
rect 635 1803 642 1805
rect 662 1803 674 1855
rect 674 1803 714 1855
rect 734 1803 780 1855
rect 780 1803 786 1855
rect 518 1771 529 1790
rect 529 1771 563 1790
rect 563 1771 570 1790
rect 518 1738 570 1771
rect 590 1771 601 1790
rect 601 1771 635 1790
rect 635 1771 642 1790
rect 590 1738 642 1771
rect 662 1738 674 1790
rect 674 1738 714 1790
rect 734 1738 780 1790
rect 780 1738 786 1790
rect 518 1698 529 1725
rect 529 1698 563 1725
rect 563 1698 570 1725
rect 518 1673 570 1698
rect 590 1698 601 1725
rect 601 1698 635 1725
rect 635 1698 642 1725
rect 590 1673 642 1698
rect 662 1673 674 1725
rect 674 1673 714 1725
rect 734 1673 780 1725
rect 780 1673 786 1725
rect 518 1659 570 1660
rect 518 1625 529 1659
rect 529 1625 563 1659
rect 563 1625 570 1659
rect 518 1608 570 1625
rect 590 1659 642 1660
rect 590 1625 601 1659
rect 601 1625 635 1659
rect 635 1625 642 1659
rect 590 1608 642 1625
rect 662 1608 674 1660
rect 674 1608 714 1660
rect 734 1608 780 1660
rect 780 1608 786 1660
rect 518 1586 570 1595
rect 518 1552 529 1586
rect 529 1552 563 1586
rect 563 1552 570 1586
rect 518 1543 570 1552
rect 590 1586 642 1595
rect 590 1552 601 1586
rect 601 1552 635 1586
rect 635 1552 642 1586
rect 590 1543 642 1552
rect 662 1543 674 1595
rect 674 1543 714 1595
rect 734 1543 780 1595
rect 780 1543 786 1595
rect 1066 4098 1118 4119
rect 1066 4067 1067 4098
rect 1067 4067 1101 4098
rect 1101 4067 1118 4098
rect 1130 4098 1182 4119
rect 1130 4067 1139 4098
rect 1139 4067 1173 4098
rect 1173 4067 1182 4098
rect 1194 4098 1246 4119
rect 1194 4067 1211 4098
rect 1211 4067 1245 4098
rect 1245 4067 1246 4098
rect 1066 4025 1118 4054
rect 1066 4002 1067 4025
rect 1067 4002 1101 4025
rect 1101 4002 1118 4025
rect 1130 4025 1182 4054
rect 1130 4002 1139 4025
rect 1139 4002 1173 4025
rect 1173 4002 1182 4025
rect 1194 4025 1246 4054
rect 1194 4002 1211 4025
rect 1211 4002 1245 4025
rect 1245 4002 1246 4025
rect 1066 3952 1118 3989
rect 1066 3937 1067 3952
rect 1067 3937 1101 3952
rect 1101 3937 1118 3952
rect 1130 3952 1182 3989
rect 1130 3937 1139 3952
rect 1139 3937 1173 3952
rect 1173 3937 1182 3952
rect 1194 3952 1246 3989
rect 1194 3937 1211 3952
rect 1211 3937 1245 3952
rect 1245 3937 1246 3952
rect 1066 3918 1067 3924
rect 1067 3918 1101 3924
rect 1101 3918 1139 3924
rect 1139 3918 1173 3924
rect 1173 3918 1211 3924
rect 1211 3918 1245 3924
rect 1245 3918 1246 3924
rect 1066 3879 1246 3918
rect 1066 3845 1067 3879
rect 1067 3845 1101 3879
rect 1101 3845 1139 3879
rect 1139 3845 1173 3879
rect 1173 3845 1211 3879
rect 1211 3845 1245 3879
rect 1245 3845 1246 3879
rect 1066 3806 1246 3845
rect 1066 3772 1067 3806
rect 1067 3772 1101 3806
rect 1101 3772 1139 3806
rect 1139 3772 1173 3806
rect 1173 3772 1211 3806
rect 1211 3772 1245 3806
rect 1245 3772 1246 3806
rect 1066 3733 1246 3772
rect 1066 3699 1067 3733
rect 1067 3699 1101 3733
rect 1101 3699 1139 3733
rect 1139 3699 1173 3733
rect 1173 3699 1211 3733
rect 1211 3699 1245 3733
rect 1245 3699 1246 3733
rect 1066 3660 1246 3699
rect 1066 3626 1067 3660
rect 1067 3626 1101 3660
rect 1101 3626 1139 3660
rect 1139 3626 1173 3660
rect 1173 3626 1211 3660
rect 1211 3626 1245 3660
rect 1245 3626 1246 3660
rect 1066 3587 1246 3626
rect 1066 3553 1067 3587
rect 1067 3553 1101 3587
rect 1101 3553 1139 3587
rect 1139 3553 1173 3587
rect 1173 3553 1211 3587
rect 1211 3553 1245 3587
rect 1245 3553 1246 3587
rect 1066 3514 1246 3553
rect 1066 3480 1067 3514
rect 1067 3480 1101 3514
rect 1101 3480 1139 3514
rect 1139 3480 1173 3514
rect 1173 3480 1211 3514
rect 1211 3480 1245 3514
rect 1245 3480 1246 3514
rect 1066 3441 1246 3480
rect 1066 3407 1067 3441
rect 1067 3407 1101 3441
rect 1101 3407 1139 3441
rect 1139 3407 1173 3441
rect 1173 3407 1211 3441
rect 1211 3407 1245 3441
rect 1245 3407 1246 3441
rect 1066 3368 1246 3407
rect 1066 3334 1067 3368
rect 1067 3334 1101 3368
rect 1101 3334 1139 3368
rect 1139 3334 1173 3368
rect 1173 3334 1211 3368
rect 1211 3334 1245 3368
rect 1245 3334 1246 3368
rect 1066 3295 1246 3334
rect 1066 3261 1067 3295
rect 1067 3261 1101 3295
rect 1101 3261 1139 3295
rect 1139 3261 1173 3295
rect 1173 3261 1211 3295
rect 1211 3261 1245 3295
rect 1245 3261 1246 3295
rect 1066 3222 1246 3261
rect 1066 3188 1067 3222
rect 1067 3188 1101 3222
rect 1101 3188 1139 3222
rect 1139 3188 1173 3222
rect 1173 3188 1211 3222
rect 1211 3188 1245 3222
rect 1245 3188 1246 3222
rect 1066 3149 1246 3188
rect 1066 3115 1067 3149
rect 1067 3115 1101 3149
rect 1101 3115 1139 3149
rect 1139 3115 1173 3149
rect 1173 3115 1211 3149
rect 1211 3115 1245 3149
rect 1245 3115 1246 3149
rect 1066 3076 1246 3115
rect 1066 3042 1067 3076
rect 1067 3042 1101 3076
rect 1101 3042 1139 3076
rect 1139 3042 1173 3076
rect 1173 3042 1211 3076
rect 1211 3042 1245 3076
rect 1245 3042 1246 3076
rect 1066 3003 1246 3042
rect 1066 2969 1067 3003
rect 1067 2969 1101 3003
rect 1101 2969 1139 3003
rect 1139 2969 1173 3003
rect 1173 2969 1211 3003
rect 1211 2969 1245 3003
rect 1245 2969 1246 3003
rect 1066 2930 1246 2969
rect 1066 2896 1067 2930
rect 1067 2896 1101 2930
rect 1101 2896 1139 2930
rect 1139 2896 1173 2930
rect 1173 2896 1211 2930
rect 1211 2896 1245 2930
rect 1245 2896 1246 2930
rect 1066 2857 1246 2896
rect 1066 2823 1067 2857
rect 1067 2823 1101 2857
rect 1101 2823 1139 2857
rect 1139 2823 1173 2857
rect 1173 2823 1211 2857
rect 1211 2823 1245 2857
rect 1245 2823 1246 2857
rect 1066 2784 1246 2823
rect 1066 2750 1067 2784
rect 1067 2750 1101 2784
rect 1101 2750 1139 2784
rect 1139 2750 1173 2784
rect 1173 2750 1211 2784
rect 1211 2750 1245 2784
rect 1245 2750 1246 2784
rect 1066 2711 1246 2750
rect 1066 2677 1067 2711
rect 1067 2677 1101 2711
rect 1101 2677 1139 2711
rect 1139 2677 1173 2711
rect 1173 2677 1211 2711
rect 1211 2677 1245 2711
rect 1245 2677 1246 2711
rect 1066 2638 1246 2677
rect 1066 2604 1067 2638
rect 1067 2604 1101 2638
rect 1101 2604 1139 2638
rect 1139 2604 1173 2638
rect 1173 2604 1211 2638
rect 1211 2604 1245 2638
rect 1245 2604 1246 2638
rect 1066 2565 1246 2604
rect 1066 2531 1067 2565
rect 1067 2531 1101 2565
rect 1101 2531 1139 2565
rect 1139 2531 1173 2565
rect 1173 2531 1211 2565
rect 1211 2531 1245 2565
rect 1245 2531 1246 2565
rect 1066 2492 1246 2531
rect 1066 2458 1067 2492
rect 1067 2458 1101 2492
rect 1101 2458 1139 2492
rect 1139 2458 1173 2492
rect 1173 2458 1211 2492
rect 1211 2458 1245 2492
rect 1245 2458 1246 2492
rect 1066 2419 1246 2458
rect 1066 2385 1067 2419
rect 1067 2385 1101 2419
rect 1101 2385 1139 2419
rect 1139 2385 1173 2419
rect 1173 2385 1211 2419
rect 1211 2385 1245 2419
rect 1245 2385 1246 2419
rect 1066 2346 1246 2385
rect 1066 2312 1067 2346
rect 1067 2312 1101 2346
rect 1101 2312 1139 2346
rect 1139 2312 1173 2346
rect 1173 2312 1211 2346
rect 1211 2312 1245 2346
rect 1245 2312 1246 2346
rect 1066 2273 1246 2312
rect 1066 2239 1067 2273
rect 1067 2239 1101 2273
rect 1101 2239 1139 2273
rect 1139 2239 1173 2273
rect 1173 2239 1211 2273
rect 1211 2239 1245 2273
rect 1245 2239 1246 2273
rect 1066 2200 1246 2239
rect 1066 2166 1067 2200
rect 1067 2166 1101 2200
rect 1101 2166 1139 2200
rect 1139 2166 1173 2200
rect 1173 2166 1211 2200
rect 1211 2166 1245 2200
rect 1245 2166 1246 2200
rect 1066 2126 1246 2166
rect 1066 2092 1067 2126
rect 1067 2092 1101 2126
rect 1101 2092 1139 2126
rect 1139 2092 1173 2126
rect 1173 2092 1211 2126
rect 1211 2092 1245 2126
rect 1245 2092 1246 2126
rect 1066 2052 1246 2092
rect 1066 2018 1067 2052
rect 1067 2018 1101 2052
rect 1101 2018 1139 2052
rect 1139 2018 1173 2052
rect 1173 2018 1211 2052
rect 1211 2018 1245 2052
rect 1245 2018 1246 2052
rect 1066 1978 1246 2018
rect 1066 1944 1067 1978
rect 1067 1944 1101 1978
rect 1101 1944 1139 1978
rect 1139 1944 1173 1978
rect 1173 1944 1211 1978
rect 1211 1944 1245 1978
rect 1245 1944 1246 1978
rect 1066 1904 1246 1944
rect 1066 1870 1067 1904
rect 1067 1870 1101 1904
rect 1101 1870 1139 1904
rect 1139 1870 1173 1904
rect 1173 1870 1211 1904
rect 1211 1870 1245 1904
rect 1245 1870 1246 1904
rect 1066 1830 1246 1870
rect 1066 1796 1067 1830
rect 1067 1796 1101 1830
rect 1101 1796 1139 1830
rect 1139 1796 1173 1830
rect 1173 1796 1211 1830
rect 1211 1796 1245 1830
rect 1245 1796 1246 1830
rect 1066 1756 1246 1796
rect 1066 1722 1067 1756
rect 1067 1722 1101 1756
rect 1101 1722 1139 1756
rect 1139 1722 1173 1756
rect 1173 1722 1211 1756
rect 1211 1722 1245 1756
rect 1245 1722 1246 1756
rect 1066 1682 1246 1722
rect 1066 1648 1067 1682
rect 1067 1648 1101 1682
rect 1101 1648 1139 1682
rect 1139 1648 1173 1682
rect 1173 1648 1211 1682
rect 1211 1648 1245 1682
rect 1245 1648 1246 1682
rect 1066 1608 1246 1648
rect 1066 1574 1067 1608
rect 1067 1574 1101 1608
rect 1101 1574 1139 1608
rect 1139 1574 1173 1608
rect 1173 1574 1211 1608
rect 1211 1574 1245 1608
rect 1245 1574 1246 1608
rect 1066 1568 1246 1574
rect 1562 4092 1614 4124
rect 1626 4118 1678 4124
rect 1626 4092 1635 4118
rect 1635 4092 1669 4118
rect 1669 4092 1678 4118
rect 1690 4092 1742 4124
rect 1562 4072 1563 4092
rect 1563 4072 1614 4092
rect 1626 4072 1678 4092
rect 1690 4072 1741 4092
rect 1741 4072 1742 4092
rect 1562 4007 1563 4059
rect 1563 4007 1614 4059
rect 1626 4007 1678 4059
rect 1690 4007 1741 4059
rect 1741 4007 1742 4059
rect 1562 3942 1563 3994
rect 1563 3942 1614 3994
rect 1626 3942 1678 3994
rect 1690 3942 1741 3994
rect 1741 3942 1742 3994
rect 1562 3877 1563 3929
rect 1563 3877 1614 3929
rect 1626 3877 1678 3929
rect 1690 3877 1741 3929
rect 1741 3877 1742 3929
rect 1562 3812 1563 3864
rect 1563 3812 1614 3864
rect 1626 3812 1678 3864
rect 1690 3812 1741 3864
rect 1741 3812 1742 3864
rect 1562 3747 1563 3799
rect 1563 3747 1614 3799
rect 1626 3747 1678 3799
rect 1690 3747 1741 3799
rect 1741 3747 1742 3799
rect 1562 3682 1563 3734
rect 1563 3682 1614 3734
rect 1626 3682 1678 3734
rect 1690 3682 1741 3734
rect 1741 3682 1742 3734
rect 1562 3617 1563 3669
rect 1563 3617 1614 3669
rect 1626 3617 1678 3669
rect 1690 3617 1741 3669
rect 1741 3617 1742 3669
rect 1562 3194 1563 3604
rect 1563 3194 1741 3604
rect 1741 3194 1742 3604
rect 1562 3182 1742 3194
rect 1562 3148 1635 3182
rect 1635 3148 1669 3182
rect 1669 3148 1742 3182
rect 1562 3108 1742 3148
rect 1562 3074 1563 3108
rect 1563 3074 1597 3108
rect 1597 3074 1635 3108
rect 1635 3074 1669 3108
rect 1669 3074 1707 3108
rect 1707 3074 1741 3108
rect 1741 3074 1742 3108
rect 1562 3028 1742 3074
rect 1562 2994 1563 3028
rect 1563 2994 1597 3028
rect 1597 2994 1635 3028
rect 1635 2994 1669 3028
rect 1669 2994 1707 3028
rect 1707 2994 1741 3028
rect 1741 2994 1742 3028
rect 1562 2948 1742 2994
rect 1562 2914 1563 2948
rect 1563 2914 1597 2948
rect 1597 2914 1635 2948
rect 1635 2914 1669 2948
rect 1669 2914 1707 2948
rect 1707 2914 1741 2948
rect 1741 2914 1742 2948
rect 1562 2868 1742 2914
rect 1562 2834 1563 2868
rect 1563 2834 1597 2868
rect 1597 2834 1635 2868
rect 1635 2834 1669 2868
rect 1669 2834 1707 2868
rect 1707 2834 1741 2868
rect 1741 2834 1742 2868
rect 1562 2788 1742 2834
rect 1562 2754 1563 2788
rect 1563 2754 1597 2788
rect 1597 2754 1635 2788
rect 1635 2754 1669 2788
rect 1669 2754 1707 2788
rect 1707 2754 1741 2788
rect 1741 2754 1742 2788
rect 1562 2708 1742 2754
rect 1562 2674 1563 2708
rect 1563 2674 1597 2708
rect 1597 2674 1635 2708
rect 1635 2674 1669 2708
rect 1669 2674 1707 2708
rect 1707 2674 1741 2708
rect 1741 2674 1742 2708
rect 1562 2628 1742 2674
rect 1562 2594 1563 2628
rect 1563 2594 1597 2628
rect 1597 2594 1635 2628
rect 1635 2594 1669 2628
rect 1669 2594 1707 2628
rect 1707 2594 1741 2628
rect 1741 2594 1742 2628
rect 1562 2556 1742 2594
rect 1562 2522 1635 2556
rect 1635 2522 1669 2556
rect 1669 2522 1742 2556
rect 1562 2518 1742 2522
rect 1562 1620 1563 2518
rect 1563 1620 1741 2518
rect 1741 1620 1742 2518
rect 1562 1586 1635 1620
rect 1635 1586 1669 1620
rect 1669 1586 1742 1620
rect 1562 1568 1742 1586
rect 2058 4098 2110 4119
rect 2058 4067 2059 4098
rect 2059 4067 2093 4098
rect 2093 4067 2110 4098
rect 2122 4098 2174 4119
rect 2122 4067 2131 4098
rect 2131 4067 2165 4098
rect 2165 4067 2174 4098
rect 2186 4098 2238 4119
rect 2186 4067 2203 4098
rect 2203 4067 2237 4098
rect 2237 4067 2238 4098
rect 2058 4025 2110 4054
rect 2058 4002 2059 4025
rect 2059 4002 2093 4025
rect 2093 4002 2110 4025
rect 2122 4025 2174 4054
rect 2122 4002 2131 4025
rect 2131 4002 2165 4025
rect 2165 4002 2174 4025
rect 2186 4025 2238 4054
rect 2186 4002 2203 4025
rect 2203 4002 2237 4025
rect 2237 4002 2238 4025
rect 2058 3952 2110 3989
rect 2058 3937 2059 3952
rect 2059 3937 2093 3952
rect 2093 3937 2110 3952
rect 2122 3952 2174 3989
rect 2122 3937 2131 3952
rect 2131 3937 2165 3952
rect 2165 3937 2174 3952
rect 2186 3952 2238 3989
rect 2186 3937 2203 3952
rect 2203 3937 2237 3952
rect 2237 3937 2238 3952
rect 2058 3918 2059 3924
rect 2059 3918 2093 3924
rect 2093 3918 2131 3924
rect 2131 3918 2165 3924
rect 2165 3918 2203 3924
rect 2203 3918 2237 3924
rect 2237 3918 2238 3924
rect 2058 3879 2238 3918
rect 2058 3845 2059 3879
rect 2059 3845 2093 3879
rect 2093 3845 2131 3879
rect 2131 3845 2165 3879
rect 2165 3845 2203 3879
rect 2203 3845 2237 3879
rect 2237 3845 2238 3879
rect 2058 3806 2238 3845
rect 2058 3772 2059 3806
rect 2059 3772 2093 3806
rect 2093 3772 2131 3806
rect 2131 3772 2165 3806
rect 2165 3772 2203 3806
rect 2203 3772 2237 3806
rect 2237 3772 2238 3806
rect 2058 3733 2238 3772
rect 2058 3699 2059 3733
rect 2059 3699 2093 3733
rect 2093 3699 2131 3733
rect 2131 3699 2165 3733
rect 2165 3699 2203 3733
rect 2203 3699 2237 3733
rect 2237 3699 2238 3733
rect 2058 3660 2238 3699
rect 2058 3626 2059 3660
rect 2059 3626 2093 3660
rect 2093 3626 2131 3660
rect 2131 3626 2165 3660
rect 2165 3626 2203 3660
rect 2203 3626 2237 3660
rect 2237 3626 2238 3660
rect 2058 3587 2238 3626
rect 2058 3553 2059 3587
rect 2059 3553 2093 3587
rect 2093 3553 2131 3587
rect 2131 3553 2165 3587
rect 2165 3553 2203 3587
rect 2203 3553 2237 3587
rect 2237 3553 2238 3587
rect 2058 3514 2238 3553
rect 2058 3480 2059 3514
rect 2059 3480 2093 3514
rect 2093 3480 2131 3514
rect 2131 3480 2165 3514
rect 2165 3480 2203 3514
rect 2203 3480 2237 3514
rect 2237 3480 2238 3514
rect 2058 3441 2238 3480
rect 2058 3407 2059 3441
rect 2059 3407 2093 3441
rect 2093 3407 2131 3441
rect 2131 3407 2165 3441
rect 2165 3407 2203 3441
rect 2203 3407 2237 3441
rect 2237 3407 2238 3441
rect 2058 3368 2238 3407
rect 2058 3334 2059 3368
rect 2059 3334 2093 3368
rect 2093 3334 2131 3368
rect 2131 3334 2165 3368
rect 2165 3334 2203 3368
rect 2203 3334 2237 3368
rect 2237 3334 2238 3368
rect 2058 3295 2238 3334
rect 2058 3261 2059 3295
rect 2059 3261 2093 3295
rect 2093 3261 2131 3295
rect 2131 3261 2165 3295
rect 2165 3261 2203 3295
rect 2203 3261 2237 3295
rect 2237 3261 2238 3295
rect 2058 3222 2238 3261
rect 2058 3188 2059 3222
rect 2059 3188 2093 3222
rect 2093 3188 2131 3222
rect 2131 3188 2165 3222
rect 2165 3188 2203 3222
rect 2203 3188 2237 3222
rect 2237 3188 2238 3222
rect 2058 3149 2238 3188
rect 2058 3115 2059 3149
rect 2059 3115 2093 3149
rect 2093 3115 2131 3149
rect 2131 3115 2165 3149
rect 2165 3115 2203 3149
rect 2203 3115 2237 3149
rect 2237 3115 2238 3149
rect 2058 3076 2238 3115
rect 2058 3042 2059 3076
rect 2059 3042 2093 3076
rect 2093 3042 2131 3076
rect 2131 3042 2165 3076
rect 2165 3042 2203 3076
rect 2203 3042 2237 3076
rect 2237 3042 2238 3076
rect 2058 3003 2238 3042
rect 2058 2969 2059 3003
rect 2059 2969 2093 3003
rect 2093 2969 2131 3003
rect 2131 2969 2165 3003
rect 2165 2969 2203 3003
rect 2203 2969 2237 3003
rect 2237 2969 2238 3003
rect 2058 2930 2238 2969
rect 2058 2896 2059 2930
rect 2059 2896 2093 2930
rect 2093 2896 2131 2930
rect 2131 2896 2165 2930
rect 2165 2896 2203 2930
rect 2203 2896 2237 2930
rect 2237 2896 2238 2930
rect 2058 2857 2238 2896
rect 2058 2823 2059 2857
rect 2059 2823 2093 2857
rect 2093 2823 2131 2857
rect 2131 2823 2165 2857
rect 2165 2823 2203 2857
rect 2203 2823 2237 2857
rect 2237 2823 2238 2857
rect 2058 2784 2238 2823
rect 2058 2750 2059 2784
rect 2059 2750 2093 2784
rect 2093 2750 2131 2784
rect 2131 2750 2165 2784
rect 2165 2750 2203 2784
rect 2203 2750 2237 2784
rect 2237 2750 2238 2784
rect 2058 2711 2238 2750
rect 2058 2677 2059 2711
rect 2059 2677 2093 2711
rect 2093 2677 2131 2711
rect 2131 2677 2165 2711
rect 2165 2677 2203 2711
rect 2203 2677 2237 2711
rect 2237 2677 2238 2711
rect 2058 2638 2238 2677
rect 2058 2604 2059 2638
rect 2059 2604 2093 2638
rect 2093 2604 2131 2638
rect 2131 2604 2165 2638
rect 2165 2604 2203 2638
rect 2203 2604 2237 2638
rect 2237 2604 2238 2638
rect 2058 2565 2238 2604
rect 2058 2531 2059 2565
rect 2059 2531 2093 2565
rect 2093 2531 2131 2565
rect 2131 2531 2165 2565
rect 2165 2531 2203 2565
rect 2203 2531 2237 2565
rect 2237 2531 2238 2565
rect 2058 2492 2238 2531
rect 2058 2458 2059 2492
rect 2059 2458 2093 2492
rect 2093 2458 2131 2492
rect 2131 2458 2165 2492
rect 2165 2458 2203 2492
rect 2203 2458 2237 2492
rect 2237 2458 2238 2492
rect 2058 2419 2238 2458
rect 2058 2385 2059 2419
rect 2059 2385 2093 2419
rect 2093 2385 2131 2419
rect 2131 2385 2165 2419
rect 2165 2385 2203 2419
rect 2203 2385 2237 2419
rect 2237 2385 2238 2419
rect 2058 2346 2238 2385
rect 2058 2312 2059 2346
rect 2059 2312 2093 2346
rect 2093 2312 2131 2346
rect 2131 2312 2165 2346
rect 2165 2312 2203 2346
rect 2203 2312 2237 2346
rect 2237 2312 2238 2346
rect 2058 2273 2238 2312
rect 2058 2239 2059 2273
rect 2059 2239 2093 2273
rect 2093 2239 2131 2273
rect 2131 2239 2165 2273
rect 2165 2239 2203 2273
rect 2203 2239 2237 2273
rect 2237 2239 2238 2273
rect 2058 2200 2238 2239
rect 2058 2166 2059 2200
rect 2059 2166 2093 2200
rect 2093 2166 2131 2200
rect 2131 2166 2165 2200
rect 2165 2166 2203 2200
rect 2203 2166 2237 2200
rect 2237 2166 2238 2200
rect 2058 2126 2238 2166
rect 2058 2092 2059 2126
rect 2059 2092 2093 2126
rect 2093 2092 2131 2126
rect 2131 2092 2165 2126
rect 2165 2092 2203 2126
rect 2203 2092 2237 2126
rect 2237 2092 2238 2126
rect 2058 2052 2238 2092
rect 2058 2018 2059 2052
rect 2059 2018 2093 2052
rect 2093 2018 2131 2052
rect 2131 2018 2165 2052
rect 2165 2018 2203 2052
rect 2203 2018 2237 2052
rect 2237 2018 2238 2052
rect 2058 1978 2238 2018
rect 2058 1944 2059 1978
rect 2059 1944 2093 1978
rect 2093 1944 2131 1978
rect 2131 1944 2165 1978
rect 2165 1944 2203 1978
rect 2203 1944 2237 1978
rect 2237 1944 2238 1978
rect 2058 1904 2238 1944
rect 2058 1870 2059 1904
rect 2059 1870 2093 1904
rect 2093 1870 2131 1904
rect 2131 1870 2165 1904
rect 2165 1870 2203 1904
rect 2203 1870 2237 1904
rect 2237 1870 2238 1904
rect 2058 1830 2238 1870
rect 2058 1796 2059 1830
rect 2059 1796 2093 1830
rect 2093 1796 2131 1830
rect 2131 1796 2165 1830
rect 2165 1796 2203 1830
rect 2203 1796 2237 1830
rect 2237 1796 2238 1830
rect 2058 1756 2238 1796
rect 2058 1722 2059 1756
rect 2059 1722 2093 1756
rect 2093 1722 2131 1756
rect 2131 1722 2165 1756
rect 2165 1722 2203 1756
rect 2203 1722 2237 1756
rect 2237 1722 2238 1756
rect 2058 1682 2238 1722
rect 2058 1648 2059 1682
rect 2059 1648 2093 1682
rect 2093 1648 2131 1682
rect 2131 1648 2165 1682
rect 2165 1648 2203 1682
rect 2203 1648 2237 1682
rect 2237 1648 2238 1682
rect 2058 1608 2238 1648
rect 2058 1574 2059 1608
rect 2059 1574 2093 1608
rect 2093 1574 2131 1608
rect 2131 1574 2165 1608
rect 2165 1574 2203 1608
rect 2203 1574 2237 1608
rect 2237 1574 2238 1608
rect 2058 1568 2238 1574
rect 2554 4092 2606 4124
rect 2618 4118 2670 4124
rect 2618 4092 2627 4118
rect 2627 4092 2661 4118
rect 2661 4092 2670 4118
rect 2682 4092 2734 4124
rect 2554 4072 2555 4092
rect 2555 4072 2606 4092
rect 2618 4072 2670 4092
rect 2682 4072 2733 4092
rect 2733 4072 2734 4092
rect 2554 4007 2555 4059
rect 2555 4007 2606 4059
rect 2618 4007 2670 4059
rect 2682 4007 2733 4059
rect 2733 4007 2734 4059
rect 2554 3942 2555 3994
rect 2555 3942 2606 3994
rect 2618 3942 2670 3994
rect 2682 3942 2733 3994
rect 2733 3942 2734 3994
rect 2554 3877 2555 3929
rect 2555 3877 2606 3929
rect 2618 3877 2670 3929
rect 2682 3877 2733 3929
rect 2733 3877 2734 3929
rect 2554 3812 2555 3864
rect 2555 3812 2606 3864
rect 2618 3812 2670 3864
rect 2682 3812 2733 3864
rect 2733 3812 2734 3864
rect 2554 3747 2555 3799
rect 2555 3747 2606 3799
rect 2618 3747 2670 3799
rect 2682 3747 2733 3799
rect 2733 3747 2734 3799
rect 2554 3682 2555 3734
rect 2555 3682 2606 3734
rect 2618 3682 2670 3734
rect 2682 3682 2733 3734
rect 2733 3682 2734 3734
rect 2554 3617 2555 3669
rect 2555 3617 2606 3669
rect 2618 3617 2670 3669
rect 2682 3617 2733 3669
rect 2733 3617 2734 3669
rect 2554 3194 2555 3604
rect 2555 3194 2733 3604
rect 2733 3194 2734 3604
rect 2554 3182 2734 3194
rect 2554 3148 2627 3182
rect 2627 3148 2661 3182
rect 2661 3148 2734 3182
rect 2554 3108 2734 3148
rect 2554 3074 2555 3108
rect 2555 3074 2589 3108
rect 2589 3074 2627 3108
rect 2627 3074 2661 3108
rect 2661 3074 2699 3108
rect 2699 3074 2733 3108
rect 2733 3074 2734 3108
rect 2554 3028 2734 3074
rect 2554 2994 2555 3028
rect 2555 2994 2589 3028
rect 2589 2994 2627 3028
rect 2627 2994 2661 3028
rect 2661 2994 2699 3028
rect 2699 2994 2733 3028
rect 2733 2994 2734 3028
rect 2554 2948 2734 2994
rect 2554 2914 2555 2948
rect 2555 2914 2589 2948
rect 2589 2914 2627 2948
rect 2627 2914 2661 2948
rect 2661 2914 2699 2948
rect 2699 2914 2733 2948
rect 2733 2914 2734 2948
rect 2554 2868 2734 2914
rect 2554 2834 2555 2868
rect 2555 2834 2589 2868
rect 2589 2834 2627 2868
rect 2627 2834 2661 2868
rect 2661 2834 2699 2868
rect 2699 2834 2733 2868
rect 2733 2834 2734 2868
rect 2554 2788 2734 2834
rect 2554 2754 2555 2788
rect 2555 2754 2589 2788
rect 2589 2754 2627 2788
rect 2627 2754 2661 2788
rect 2661 2754 2699 2788
rect 2699 2754 2733 2788
rect 2733 2754 2734 2788
rect 2554 2708 2734 2754
rect 2554 2674 2555 2708
rect 2555 2674 2589 2708
rect 2589 2674 2627 2708
rect 2627 2674 2661 2708
rect 2661 2674 2699 2708
rect 2699 2674 2733 2708
rect 2733 2674 2734 2708
rect 2554 2628 2734 2674
rect 2554 2594 2555 2628
rect 2555 2594 2589 2628
rect 2589 2594 2627 2628
rect 2627 2594 2661 2628
rect 2661 2594 2699 2628
rect 2699 2594 2733 2628
rect 2733 2594 2734 2628
rect 2554 2556 2734 2594
rect 2554 2522 2627 2556
rect 2627 2522 2661 2556
rect 2661 2522 2734 2556
rect 2554 2518 2734 2522
rect 2554 1620 2555 2518
rect 2555 1620 2733 2518
rect 2733 1620 2734 2518
rect 2554 1586 2627 1620
rect 2627 1586 2661 1620
rect 2661 1586 2734 1620
rect 2554 1568 2734 1586
rect 3050 4098 3102 4119
rect 3050 4067 3051 4098
rect 3051 4067 3085 4098
rect 3085 4067 3102 4098
rect 3114 4098 3166 4119
rect 3114 4067 3123 4098
rect 3123 4067 3157 4098
rect 3157 4067 3166 4098
rect 3178 4098 3230 4119
rect 3178 4067 3195 4098
rect 3195 4067 3229 4098
rect 3229 4067 3230 4098
rect 3050 4025 3102 4054
rect 3050 4002 3051 4025
rect 3051 4002 3085 4025
rect 3085 4002 3102 4025
rect 3114 4025 3166 4054
rect 3114 4002 3123 4025
rect 3123 4002 3157 4025
rect 3157 4002 3166 4025
rect 3178 4025 3230 4054
rect 3178 4002 3195 4025
rect 3195 4002 3229 4025
rect 3229 4002 3230 4025
rect 3050 3952 3102 3989
rect 3050 3937 3051 3952
rect 3051 3937 3085 3952
rect 3085 3937 3102 3952
rect 3114 3952 3166 3989
rect 3114 3937 3123 3952
rect 3123 3937 3157 3952
rect 3157 3937 3166 3952
rect 3178 3952 3230 3989
rect 3178 3937 3195 3952
rect 3195 3937 3229 3952
rect 3229 3937 3230 3952
rect 3050 3918 3051 3924
rect 3051 3918 3085 3924
rect 3085 3918 3123 3924
rect 3123 3918 3157 3924
rect 3157 3918 3195 3924
rect 3195 3918 3229 3924
rect 3229 3918 3230 3924
rect 3050 3879 3230 3918
rect 3050 3845 3051 3879
rect 3051 3845 3085 3879
rect 3085 3845 3123 3879
rect 3123 3845 3157 3879
rect 3157 3845 3195 3879
rect 3195 3845 3229 3879
rect 3229 3845 3230 3879
rect 3050 3806 3230 3845
rect 3050 3772 3051 3806
rect 3051 3772 3085 3806
rect 3085 3772 3123 3806
rect 3123 3772 3157 3806
rect 3157 3772 3195 3806
rect 3195 3772 3229 3806
rect 3229 3772 3230 3806
rect 3050 3733 3230 3772
rect 3050 3699 3051 3733
rect 3051 3699 3085 3733
rect 3085 3699 3123 3733
rect 3123 3699 3157 3733
rect 3157 3699 3195 3733
rect 3195 3699 3229 3733
rect 3229 3699 3230 3733
rect 3050 3660 3230 3699
rect 3050 3626 3051 3660
rect 3051 3626 3085 3660
rect 3085 3626 3123 3660
rect 3123 3626 3157 3660
rect 3157 3626 3195 3660
rect 3195 3626 3229 3660
rect 3229 3626 3230 3660
rect 3050 3587 3230 3626
rect 3050 3553 3051 3587
rect 3051 3553 3085 3587
rect 3085 3553 3123 3587
rect 3123 3553 3157 3587
rect 3157 3553 3195 3587
rect 3195 3553 3229 3587
rect 3229 3553 3230 3587
rect 3050 3514 3230 3553
rect 3050 3480 3051 3514
rect 3051 3480 3085 3514
rect 3085 3480 3123 3514
rect 3123 3480 3157 3514
rect 3157 3480 3195 3514
rect 3195 3480 3229 3514
rect 3229 3480 3230 3514
rect 3050 3441 3230 3480
rect 3050 3407 3051 3441
rect 3051 3407 3085 3441
rect 3085 3407 3123 3441
rect 3123 3407 3157 3441
rect 3157 3407 3195 3441
rect 3195 3407 3229 3441
rect 3229 3407 3230 3441
rect 3050 3368 3230 3407
rect 3050 3334 3051 3368
rect 3051 3334 3085 3368
rect 3085 3334 3123 3368
rect 3123 3334 3157 3368
rect 3157 3334 3195 3368
rect 3195 3334 3229 3368
rect 3229 3334 3230 3368
rect 3050 3295 3230 3334
rect 3050 3261 3051 3295
rect 3051 3261 3085 3295
rect 3085 3261 3123 3295
rect 3123 3261 3157 3295
rect 3157 3261 3195 3295
rect 3195 3261 3229 3295
rect 3229 3261 3230 3295
rect 3050 3222 3230 3261
rect 3050 3188 3051 3222
rect 3051 3188 3085 3222
rect 3085 3188 3123 3222
rect 3123 3188 3157 3222
rect 3157 3188 3195 3222
rect 3195 3188 3229 3222
rect 3229 3188 3230 3222
rect 3050 3149 3230 3188
rect 3050 3115 3051 3149
rect 3051 3115 3085 3149
rect 3085 3115 3123 3149
rect 3123 3115 3157 3149
rect 3157 3115 3195 3149
rect 3195 3115 3229 3149
rect 3229 3115 3230 3149
rect 3050 3076 3230 3115
rect 3050 3042 3051 3076
rect 3051 3042 3085 3076
rect 3085 3042 3123 3076
rect 3123 3042 3157 3076
rect 3157 3042 3195 3076
rect 3195 3042 3229 3076
rect 3229 3042 3230 3076
rect 3050 3003 3230 3042
rect 3050 2969 3051 3003
rect 3051 2969 3085 3003
rect 3085 2969 3123 3003
rect 3123 2969 3157 3003
rect 3157 2969 3195 3003
rect 3195 2969 3229 3003
rect 3229 2969 3230 3003
rect 3050 2930 3230 2969
rect 3050 2896 3051 2930
rect 3051 2896 3085 2930
rect 3085 2896 3123 2930
rect 3123 2896 3157 2930
rect 3157 2896 3195 2930
rect 3195 2896 3229 2930
rect 3229 2896 3230 2930
rect 3050 2857 3230 2896
rect 3050 2823 3051 2857
rect 3051 2823 3085 2857
rect 3085 2823 3123 2857
rect 3123 2823 3157 2857
rect 3157 2823 3195 2857
rect 3195 2823 3229 2857
rect 3229 2823 3230 2857
rect 3050 2784 3230 2823
rect 3050 2750 3051 2784
rect 3051 2750 3085 2784
rect 3085 2750 3123 2784
rect 3123 2750 3157 2784
rect 3157 2750 3195 2784
rect 3195 2750 3229 2784
rect 3229 2750 3230 2784
rect 3050 2711 3230 2750
rect 3050 2677 3051 2711
rect 3051 2677 3085 2711
rect 3085 2677 3123 2711
rect 3123 2677 3157 2711
rect 3157 2677 3195 2711
rect 3195 2677 3229 2711
rect 3229 2677 3230 2711
rect 3050 2638 3230 2677
rect 3050 2604 3051 2638
rect 3051 2604 3085 2638
rect 3085 2604 3123 2638
rect 3123 2604 3157 2638
rect 3157 2604 3195 2638
rect 3195 2604 3229 2638
rect 3229 2604 3230 2638
rect 3050 2565 3230 2604
rect 3050 2531 3051 2565
rect 3051 2531 3085 2565
rect 3085 2531 3123 2565
rect 3123 2531 3157 2565
rect 3157 2531 3195 2565
rect 3195 2531 3229 2565
rect 3229 2531 3230 2565
rect 3050 2492 3230 2531
rect 3050 2458 3051 2492
rect 3051 2458 3085 2492
rect 3085 2458 3123 2492
rect 3123 2458 3157 2492
rect 3157 2458 3195 2492
rect 3195 2458 3229 2492
rect 3229 2458 3230 2492
rect 3050 2419 3230 2458
rect 3050 2385 3051 2419
rect 3051 2385 3085 2419
rect 3085 2385 3123 2419
rect 3123 2385 3157 2419
rect 3157 2385 3195 2419
rect 3195 2385 3229 2419
rect 3229 2385 3230 2419
rect 3050 2346 3230 2385
rect 3050 2312 3051 2346
rect 3051 2312 3085 2346
rect 3085 2312 3123 2346
rect 3123 2312 3157 2346
rect 3157 2312 3195 2346
rect 3195 2312 3229 2346
rect 3229 2312 3230 2346
rect 3050 2273 3230 2312
rect 3050 2239 3051 2273
rect 3051 2239 3085 2273
rect 3085 2239 3123 2273
rect 3123 2239 3157 2273
rect 3157 2239 3195 2273
rect 3195 2239 3229 2273
rect 3229 2239 3230 2273
rect 3050 2200 3230 2239
rect 3050 2166 3051 2200
rect 3051 2166 3085 2200
rect 3085 2166 3123 2200
rect 3123 2166 3157 2200
rect 3157 2166 3195 2200
rect 3195 2166 3229 2200
rect 3229 2166 3230 2200
rect 3050 2126 3230 2166
rect 3050 2092 3051 2126
rect 3051 2092 3085 2126
rect 3085 2092 3123 2126
rect 3123 2092 3157 2126
rect 3157 2092 3195 2126
rect 3195 2092 3229 2126
rect 3229 2092 3230 2126
rect 3050 2052 3230 2092
rect 3050 2018 3051 2052
rect 3051 2018 3085 2052
rect 3085 2018 3123 2052
rect 3123 2018 3157 2052
rect 3157 2018 3195 2052
rect 3195 2018 3229 2052
rect 3229 2018 3230 2052
rect 3050 1978 3230 2018
rect 3050 1944 3051 1978
rect 3051 1944 3085 1978
rect 3085 1944 3123 1978
rect 3123 1944 3157 1978
rect 3157 1944 3195 1978
rect 3195 1944 3229 1978
rect 3229 1944 3230 1978
rect 3050 1904 3230 1944
rect 3050 1870 3051 1904
rect 3051 1870 3085 1904
rect 3085 1870 3123 1904
rect 3123 1870 3157 1904
rect 3157 1870 3195 1904
rect 3195 1870 3229 1904
rect 3229 1870 3230 1904
rect 3050 1830 3230 1870
rect 3050 1796 3051 1830
rect 3051 1796 3085 1830
rect 3085 1796 3123 1830
rect 3123 1796 3157 1830
rect 3157 1796 3195 1830
rect 3195 1796 3229 1830
rect 3229 1796 3230 1830
rect 3050 1756 3230 1796
rect 3050 1722 3051 1756
rect 3051 1722 3085 1756
rect 3085 1722 3123 1756
rect 3123 1722 3157 1756
rect 3157 1722 3195 1756
rect 3195 1722 3229 1756
rect 3229 1722 3230 1756
rect 3050 1682 3230 1722
rect 3050 1648 3051 1682
rect 3051 1648 3085 1682
rect 3085 1648 3123 1682
rect 3123 1648 3157 1682
rect 3157 1648 3195 1682
rect 3195 1648 3229 1682
rect 3229 1648 3230 1682
rect 3050 1608 3230 1648
rect 3050 1574 3051 1608
rect 3051 1574 3085 1608
rect 3085 1574 3123 1608
rect 3123 1574 3157 1608
rect 3157 1574 3195 1608
rect 3195 1574 3229 1608
rect 3229 1574 3230 1608
rect 3050 1568 3230 1574
rect 3546 4092 3598 4124
rect 3610 4118 3662 4124
rect 3610 4092 3619 4118
rect 3619 4092 3653 4118
rect 3653 4092 3662 4118
rect 3674 4092 3726 4124
rect 3546 4072 3547 4092
rect 3547 4072 3598 4092
rect 3610 4072 3662 4092
rect 3674 4072 3725 4092
rect 3725 4072 3726 4092
rect 3546 4007 3547 4059
rect 3547 4007 3598 4059
rect 3610 4007 3662 4059
rect 3674 4007 3725 4059
rect 3725 4007 3726 4059
rect 3546 3942 3547 3994
rect 3547 3942 3598 3994
rect 3610 3942 3662 3994
rect 3674 3942 3725 3994
rect 3725 3942 3726 3994
rect 3546 3877 3547 3929
rect 3547 3877 3598 3929
rect 3610 3877 3662 3929
rect 3674 3877 3725 3929
rect 3725 3877 3726 3929
rect 3546 3812 3547 3864
rect 3547 3812 3598 3864
rect 3610 3812 3662 3864
rect 3674 3812 3725 3864
rect 3725 3812 3726 3864
rect 3546 3747 3547 3799
rect 3547 3747 3598 3799
rect 3610 3747 3662 3799
rect 3674 3747 3725 3799
rect 3725 3747 3726 3799
rect 3546 3682 3547 3734
rect 3547 3682 3598 3734
rect 3610 3682 3662 3734
rect 3674 3682 3725 3734
rect 3725 3682 3726 3734
rect 3546 3617 3547 3669
rect 3547 3617 3598 3669
rect 3610 3617 3662 3669
rect 3674 3617 3725 3669
rect 3725 3617 3726 3669
rect 3546 3194 3547 3604
rect 3547 3194 3725 3604
rect 3725 3194 3726 3604
rect 3546 3182 3726 3194
rect 3546 3148 3619 3182
rect 3619 3148 3653 3182
rect 3653 3148 3726 3182
rect 3546 3108 3726 3148
rect 3546 3074 3547 3108
rect 3547 3074 3581 3108
rect 3581 3074 3619 3108
rect 3619 3074 3653 3108
rect 3653 3074 3691 3108
rect 3691 3074 3725 3108
rect 3725 3074 3726 3108
rect 3546 3028 3726 3074
rect 3546 2994 3547 3028
rect 3547 2994 3581 3028
rect 3581 2994 3619 3028
rect 3619 2994 3653 3028
rect 3653 2994 3691 3028
rect 3691 2994 3725 3028
rect 3725 2994 3726 3028
rect 3546 2948 3726 2994
rect 3546 2914 3547 2948
rect 3547 2914 3581 2948
rect 3581 2914 3619 2948
rect 3619 2914 3653 2948
rect 3653 2914 3691 2948
rect 3691 2914 3725 2948
rect 3725 2914 3726 2948
rect 3546 2868 3726 2914
rect 3546 2834 3547 2868
rect 3547 2834 3581 2868
rect 3581 2834 3619 2868
rect 3619 2834 3653 2868
rect 3653 2834 3691 2868
rect 3691 2834 3725 2868
rect 3725 2834 3726 2868
rect 3546 2788 3726 2834
rect 3546 2754 3547 2788
rect 3547 2754 3581 2788
rect 3581 2754 3619 2788
rect 3619 2754 3653 2788
rect 3653 2754 3691 2788
rect 3691 2754 3725 2788
rect 3725 2754 3726 2788
rect 3546 2708 3726 2754
rect 3546 2674 3547 2708
rect 3547 2674 3581 2708
rect 3581 2674 3619 2708
rect 3619 2674 3653 2708
rect 3653 2674 3691 2708
rect 3691 2674 3725 2708
rect 3725 2674 3726 2708
rect 3546 2628 3726 2674
rect 3546 2594 3547 2628
rect 3547 2594 3581 2628
rect 3581 2594 3619 2628
rect 3619 2594 3653 2628
rect 3653 2594 3691 2628
rect 3691 2594 3725 2628
rect 3725 2594 3726 2628
rect 3546 2556 3726 2594
rect 3546 2522 3619 2556
rect 3619 2522 3653 2556
rect 3653 2522 3726 2556
rect 3546 2518 3726 2522
rect 3546 1620 3547 2518
rect 3547 1620 3725 2518
rect 3725 1620 3726 2518
rect 3546 1586 3619 1620
rect 3619 1586 3653 1620
rect 3653 1586 3726 1620
rect 3546 1568 3726 1586
rect 4042 4098 4094 4119
rect 4042 4067 4043 4098
rect 4043 4067 4077 4098
rect 4077 4067 4094 4098
rect 4106 4098 4158 4119
rect 4106 4067 4115 4098
rect 4115 4067 4149 4098
rect 4149 4067 4158 4098
rect 4170 4098 4222 4119
rect 4170 4067 4187 4098
rect 4187 4067 4221 4098
rect 4221 4067 4222 4098
rect 4042 4025 4094 4054
rect 4042 4002 4043 4025
rect 4043 4002 4077 4025
rect 4077 4002 4094 4025
rect 4106 4025 4158 4054
rect 4106 4002 4115 4025
rect 4115 4002 4149 4025
rect 4149 4002 4158 4025
rect 4170 4025 4222 4054
rect 4170 4002 4187 4025
rect 4187 4002 4221 4025
rect 4221 4002 4222 4025
rect 4042 3952 4094 3989
rect 4042 3937 4043 3952
rect 4043 3937 4077 3952
rect 4077 3937 4094 3952
rect 4106 3952 4158 3989
rect 4106 3937 4115 3952
rect 4115 3937 4149 3952
rect 4149 3937 4158 3952
rect 4170 3952 4222 3989
rect 4170 3937 4187 3952
rect 4187 3937 4221 3952
rect 4221 3937 4222 3952
rect 4042 3918 4043 3924
rect 4043 3918 4077 3924
rect 4077 3918 4115 3924
rect 4115 3918 4149 3924
rect 4149 3918 4187 3924
rect 4187 3918 4221 3924
rect 4221 3918 4222 3924
rect 4042 3879 4222 3918
rect 4042 3845 4043 3879
rect 4043 3845 4077 3879
rect 4077 3845 4115 3879
rect 4115 3845 4149 3879
rect 4149 3845 4187 3879
rect 4187 3845 4221 3879
rect 4221 3845 4222 3879
rect 4042 3806 4222 3845
rect 4042 3772 4043 3806
rect 4043 3772 4077 3806
rect 4077 3772 4115 3806
rect 4115 3772 4149 3806
rect 4149 3772 4187 3806
rect 4187 3772 4221 3806
rect 4221 3772 4222 3806
rect 4042 3733 4222 3772
rect 4042 3699 4043 3733
rect 4043 3699 4077 3733
rect 4077 3699 4115 3733
rect 4115 3699 4149 3733
rect 4149 3699 4187 3733
rect 4187 3699 4221 3733
rect 4221 3699 4222 3733
rect 4042 3660 4222 3699
rect 4042 3626 4043 3660
rect 4043 3626 4077 3660
rect 4077 3626 4115 3660
rect 4115 3626 4149 3660
rect 4149 3626 4187 3660
rect 4187 3626 4221 3660
rect 4221 3626 4222 3660
rect 4042 3587 4222 3626
rect 4042 3553 4043 3587
rect 4043 3553 4077 3587
rect 4077 3553 4115 3587
rect 4115 3553 4149 3587
rect 4149 3553 4187 3587
rect 4187 3553 4221 3587
rect 4221 3553 4222 3587
rect 4042 3514 4222 3553
rect 4042 3480 4043 3514
rect 4043 3480 4077 3514
rect 4077 3480 4115 3514
rect 4115 3480 4149 3514
rect 4149 3480 4187 3514
rect 4187 3480 4221 3514
rect 4221 3480 4222 3514
rect 4042 3441 4222 3480
rect 4042 3407 4043 3441
rect 4043 3407 4077 3441
rect 4077 3407 4115 3441
rect 4115 3407 4149 3441
rect 4149 3407 4187 3441
rect 4187 3407 4221 3441
rect 4221 3407 4222 3441
rect 4042 3368 4222 3407
rect 4042 3334 4043 3368
rect 4043 3334 4077 3368
rect 4077 3334 4115 3368
rect 4115 3334 4149 3368
rect 4149 3334 4187 3368
rect 4187 3334 4221 3368
rect 4221 3334 4222 3368
rect 4042 3295 4222 3334
rect 4042 3261 4043 3295
rect 4043 3261 4077 3295
rect 4077 3261 4115 3295
rect 4115 3261 4149 3295
rect 4149 3261 4187 3295
rect 4187 3261 4221 3295
rect 4221 3261 4222 3295
rect 4042 3222 4222 3261
rect 4042 3188 4043 3222
rect 4043 3188 4077 3222
rect 4077 3188 4115 3222
rect 4115 3188 4149 3222
rect 4149 3188 4187 3222
rect 4187 3188 4221 3222
rect 4221 3188 4222 3222
rect 4042 3149 4222 3188
rect 4042 3115 4043 3149
rect 4043 3115 4077 3149
rect 4077 3115 4115 3149
rect 4115 3115 4149 3149
rect 4149 3115 4187 3149
rect 4187 3115 4221 3149
rect 4221 3115 4222 3149
rect 4042 3076 4222 3115
rect 4042 3042 4043 3076
rect 4043 3042 4077 3076
rect 4077 3042 4115 3076
rect 4115 3042 4149 3076
rect 4149 3042 4187 3076
rect 4187 3042 4221 3076
rect 4221 3042 4222 3076
rect 4042 3003 4222 3042
rect 4042 2969 4043 3003
rect 4043 2969 4077 3003
rect 4077 2969 4115 3003
rect 4115 2969 4149 3003
rect 4149 2969 4187 3003
rect 4187 2969 4221 3003
rect 4221 2969 4222 3003
rect 4042 2930 4222 2969
rect 4042 2896 4043 2930
rect 4043 2896 4077 2930
rect 4077 2896 4115 2930
rect 4115 2896 4149 2930
rect 4149 2896 4187 2930
rect 4187 2896 4221 2930
rect 4221 2896 4222 2930
rect 4042 2857 4222 2896
rect 4042 2823 4043 2857
rect 4043 2823 4077 2857
rect 4077 2823 4115 2857
rect 4115 2823 4149 2857
rect 4149 2823 4187 2857
rect 4187 2823 4221 2857
rect 4221 2823 4222 2857
rect 4042 2784 4222 2823
rect 4042 2750 4043 2784
rect 4043 2750 4077 2784
rect 4077 2750 4115 2784
rect 4115 2750 4149 2784
rect 4149 2750 4187 2784
rect 4187 2750 4221 2784
rect 4221 2750 4222 2784
rect 4042 2711 4222 2750
rect 4042 2677 4043 2711
rect 4043 2677 4077 2711
rect 4077 2677 4115 2711
rect 4115 2677 4149 2711
rect 4149 2677 4187 2711
rect 4187 2677 4221 2711
rect 4221 2677 4222 2711
rect 4042 2638 4222 2677
rect 4042 2604 4043 2638
rect 4043 2604 4077 2638
rect 4077 2604 4115 2638
rect 4115 2604 4149 2638
rect 4149 2604 4187 2638
rect 4187 2604 4221 2638
rect 4221 2604 4222 2638
rect 4042 2565 4222 2604
rect 4042 2531 4043 2565
rect 4043 2531 4077 2565
rect 4077 2531 4115 2565
rect 4115 2531 4149 2565
rect 4149 2531 4187 2565
rect 4187 2531 4221 2565
rect 4221 2531 4222 2565
rect 4042 2492 4222 2531
rect 4042 2458 4043 2492
rect 4043 2458 4077 2492
rect 4077 2458 4115 2492
rect 4115 2458 4149 2492
rect 4149 2458 4187 2492
rect 4187 2458 4221 2492
rect 4221 2458 4222 2492
rect 4042 2419 4222 2458
rect 4042 2385 4043 2419
rect 4043 2385 4077 2419
rect 4077 2385 4115 2419
rect 4115 2385 4149 2419
rect 4149 2385 4187 2419
rect 4187 2385 4221 2419
rect 4221 2385 4222 2419
rect 4042 2346 4222 2385
rect 4042 2312 4043 2346
rect 4043 2312 4077 2346
rect 4077 2312 4115 2346
rect 4115 2312 4149 2346
rect 4149 2312 4187 2346
rect 4187 2312 4221 2346
rect 4221 2312 4222 2346
rect 4042 2273 4222 2312
rect 4042 2239 4043 2273
rect 4043 2239 4077 2273
rect 4077 2239 4115 2273
rect 4115 2239 4149 2273
rect 4149 2239 4187 2273
rect 4187 2239 4221 2273
rect 4221 2239 4222 2273
rect 4042 2200 4222 2239
rect 4042 2166 4043 2200
rect 4043 2166 4077 2200
rect 4077 2166 4115 2200
rect 4115 2166 4149 2200
rect 4149 2166 4187 2200
rect 4187 2166 4221 2200
rect 4221 2166 4222 2200
rect 4042 2126 4222 2166
rect 4042 2092 4043 2126
rect 4043 2092 4077 2126
rect 4077 2092 4115 2126
rect 4115 2092 4149 2126
rect 4149 2092 4187 2126
rect 4187 2092 4221 2126
rect 4221 2092 4222 2126
rect 4042 2052 4222 2092
rect 4042 2018 4043 2052
rect 4043 2018 4077 2052
rect 4077 2018 4115 2052
rect 4115 2018 4149 2052
rect 4149 2018 4187 2052
rect 4187 2018 4221 2052
rect 4221 2018 4222 2052
rect 4042 1978 4222 2018
rect 4042 1944 4043 1978
rect 4043 1944 4077 1978
rect 4077 1944 4115 1978
rect 4115 1944 4149 1978
rect 4149 1944 4187 1978
rect 4187 1944 4221 1978
rect 4221 1944 4222 1978
rect 4042 1904 4222 1944
rect 4042 1870 4043 1904
rect 4043 1870 4077 1904
rect 4077 1870 4115 1904
rect 4115 1870 4149 1904
rect 4149 1870 4187 1904
rect 4187 1870 4221 1904
rect 4221 1870 4222 1904
rect 4042 1830 4222 1870
rect 4042 1796 4043 1830
rect 4043 1796 4077 1830
rect 4077 1796 4115 1830
rect 4115 1796 4149 1830
rect 4149 1796 4187 1830
rect 4187 1796 4221 1830
rect 4221 1796 4222 1830
rect 4042 1756 4222 1796
rect 4042 1722 4043 1756
rect 4043 1722 4077 1756
rect 4077 1722 4115 1756
rect 4115 1722 4149 1756
rect 4149 1722 4187 1756
rect 4187 1722 4221 1756
rect 4221 1722 4222 1756
rect 4042 1682 4222 1722
rect 4042 1648 4043 1682
rect 4043 1648 4077 1682
rect 4077 1648 4115 1682
rect 4115 1648 4149 1682
rect 4149 1648 4187 1682
rect 4187 1648 4221 1682
rect 4221 1648 4222 1682
rect 4042 1608 4222 1648
rect 4042 1574 4043 1608
rect 4043 1574 4077 1608
rect 4077 1574 4115 1608
rect 4115 1574 4149 1608
rect 4149 1574 4187 1608
rect 4187 1574 4221 1608
rect 4221 1574 4222 1608
rect 4042 1568 4222 1574
rect 4538 4092 4590 4124
rect 4602 4118 4654 4124
rect 4602 4092 4611 4118
rect 4611 4092 4645 4118
rect 4645 4092 4654 4118
rect 4666 4092 4718 4124
rect 4538 4072 4539 4092
rect 4539 4072 4590 4092
rect 4602 4072 4654 4092
rect 4666 4072 4717 4092
rect 4717 4072 4718 4092
rect 4538 4007 4539 4059
rect 4539 4007 4590 4059
rect 4602 4007 4654 4059
rect 4666 4007 4717 4059
rect 4717 4007 4718 4059
rect 4538 3942 4539 3994
rect 4539 3942 4590 3994
rect 4602 3942 4654 3994
rect 4666 3942 4717 3994
rect 4717 3942 4718 3994
rect 4538 3877 4539 3929
rect 4539 3877 4590 3929
rect 4602 3877 4654 3929
rect 4666 3877 4717 3929
rect 4717 3877 4718 3929
rect 4538 3812 4539 3864
rect 4539 3812 4590 3864
rect 4602 3812 4654 3864
rect 4666 3812 4717 3864
rect 4717 3812 4718 3864
rect 4538 3747 4539 3799
rect 4539 3747 4590 3799
rect 4602 3747 4654 3799
rect 4666 3747 4717 3799
rect 4717 3747 4718 3799
rect 4538 3682 4539 3734
rect 4539 3682 4590 3734
rect 4602 3682 4654 3734
rect 4666 3682 4717 3734
rect 4717 3682 4718 3734
rect 4538 3617 4539 3669
rect 4539 3617 4590 3669
rect 4602 3617 4654 3669
rect 4666 3617 4717 3669
rect 4717 3617 4718 3669
rect 4538 3194 4539 3604
rect 4539 3194 4717 3604
rect 4717 3194 4718 3604
rect 4538 3182 4718 3194
rect 4538 3148 4611 3182
rect 4611 3148 4645 3182
rect 4645 3148 4718 3182
rect 4538 3108 4718 3148
rect 4538 3074 4539 3108
rect 4539 3074 4573 3108
rect 4573 3074 4611 3108
rect 4611 3074 4645 3108
rect 4645 3074 4683 3108
rect 4683 3074 4717 3108
rect 4717 3074 4718 3108
rect 4538 3028 4718 3074
rect 4538 2994 4539 3028
rect 4539 2994 4573 3028
rect 4573 2994 4611 3028
rect 4611 2994 4645 3028
rect 4645 2994 4683 3028
rect 4683 2994 4717 3028
rect 4717 2994 4718 3028
rect 4538 2948 4718 2994
rect 4538 2914 4539 2948
rect 4539 2914 4573 2948
rect 4573 2914 4611 2948
rect 4611 2914 4645 2948
rect 4645 2914 4683 2948
rect 4683 2914 4717 2948
rect 4717 2914 4718 2948
rect 4538 2868 4718 2914
rect 4538 2834 4539 2868
rect 4539 2834 4573 2868
rect 4573 2834 4611 2868
rect 4611 2834 4645 2868
rect 4645 2834 4683 2868
rect 4683 2834 4717 2868
rect 4717 2834 4718 2868
rect 4538 2788 4718 2834
rect 4538 2754 4539 2788
rect 4539 2754 4573 2788
rect 4573 2754 4611 2788
rect 4611 2754 4645 2788
rect 4645 2754 4683 2788
rect 4683 2754 4717 2788
rect 4717 2754 4718 2788
rect 4538 2708 4718 2754
rect 4538 2674 4539 2708
rect 4539 2674 4573 2708
rect 4573 2674 4611 2708
rect 4611 2674 4645 2708
rect 4645 2674 4683 2708
rect 4683 2674 4717 2708
rect 4717 2674 4718 2708
rect 4538 2628 4718 2674
rect 4538 2594 4539 2628
rect 4539 2594 4573 2628
rect 4573 2594 4611 2628
rect 4611 2594 4645 2628
rect 4645 2594 4683 2628
rect 4683 2594 4717 2628
rect 4717 2594 4718 2628
rect 4538 2556 4718 2594
rect 4538 2522 4611 2556
rect 4611 2522 4645 2556
rect 4645 2522 4718 2556
rect 4538 2518 4718 2522
rect 4538 1620 4539 2518
rect 4539 1620 4717 2518
rect 4717 1620 4718 2518
rect 4538 1586 4611 1620
rect 4611 1586 4645 1620
rect 4645 1586 4718 1620
rect 4538 1568 4718 1586
rect 5034 4098 5086 4119
rect 5034 4067 5035 4098
rect 5035 4067 5069 4098
rect 5069 4067 5086 4098
rect 5098 4098 5150 4119
rect 5098 4067 5107 4098
rect 5107 4067 5141 4098
rect 5141 4067 5150 4098
rect 5162 4098 5214 4119
rect 5162 4067 5179 4098
rect 5179 4067 5213 4098
rect 5213 4067 5214 4098
rect 5034 4025 5086 4054
rect 5034 4002 5035 4025
rect 5035 4002 5069 4025
rect 5069 4002 5086 4025
rect 5098 4025 5150 4054
rect 5098 4002 5107 4025
rect 5107 4002 5141 4025
rect 5141 4002 5150 4025
rect 5162 4025 5214 4054
rect 5162 4002 5179 4025
rect 5179 4002 5213 4025
rect 5213 4002 5214 4025
rect 5034 3952 5086 3989
rect 5034 3937 5035 3952
rect 5035 3937 5069 3952
rect 5069 3937 5086 3952
rect 5098 3952 5150 3989
rect 5098 3937 5107 3952
rect 5107 3937 5141 3952
rect 5141 3937 5150 3952
rect 5162 3952 5214 3989
rect 5162 3937 5179 3952
rect 5179 3937 5213 3952
rect 5213 3937 5214 3952
rect 5034 3918 5035 3924
rect 5035 3918 5069 3924
rect 5069 3918 5107 3924
rect 5107 3918 5141 3924
rect 5141 3918 5179 3924
rect 5179 3918 5213 3924
rect 5213 3918 5214 3924
rect 5034 3879 5214 3918
rect 5034 3845 5035 3879
rect 5035 3845 5069 3879
rect 5069 3845 5107 3879
rect 5107 3845 5141 3879
rect 5141 3845 5179 3879
rect 5179 3845 5213 3879
rect 5213 3845 5214 3879
rect 5034 3806 5214 3845
rect 5034 3772 5035 3806
rect 5035 3772 5069 3806
rect 5069 3772 5107 3806
rect 5107 3772 5141 3806
rect 5141 3772 5179 3806
rect 5179 3772 5213 3806
rect 5213 3772 5214 3806
rect 5034 3733 5214 3772
rect 5034 3699 5035 3733
rect 5035 3699 5069 3733
rect 5069 3699 5107 3733
rect 5107 3699 5141 3733
rect 5141 3699 5179 3733
rect 5179 3699 5213 3733
rect 5213 3699 5214 3733
rect 5034 3660 5214 3699
rect 5034 3626 5035 3660
rect 5035 3626 5069 3660
rect 5069 3626 5107 3660
rect 5107 3626 5141 3660
rect 5141 3626 5179 3660
rect 5179 3626 5213 3660
rect 5213 3626 5214 3660
rect 5034 3587 5214 3626
rect 5034 3553 5035 3587
rect 5035 3553 5069 3587
rect 5069 3553 5107 3587
rect 5107 3553 5141 3587
rect 5141 3553 5179 3587
rect 5179 3553 5213 3587
rect 5213 3553 5214 3587
rect 5034 3514 5214 3553
rect 5034 3480 5035 3514
rect 5035 3480 5069 3514
rect 5069 3480 5107 3514
rect 5107 3480 5141 3514
rect 5141 3480 5179 3514
rect 5179 3480 5213 3514
rect 5213 3480 5214 3514
rect 5034 3441 5214 3480
rect 5034 3407 5035 3441
rect 5035 3407 5069 3441
rect 5069 3407 5107 3441
rect 5107 3407 5141 3441
rect 5141 3407 5179 3441
rect 5179 3407 5213 3441
rect 5213 3407 5214 3441
rect 5034 3368 5214 3407
rect 5034 3334 5035 3368
rect 5035 3334 5069 3368
rect 5069 3334 5107 3368
rect 5107 3334 5141 3368
rect 5141 3334 5179 3368
rect 5179 3334 5213 3368
rect 5213 3334 5214 3368
rect 5034 3295 5214 3334
rect 5034 3261 5035 3295
rect 5035 3261 5069 3295
rect 5069 3261 5107 3295
rect 5107 3261 5141 3295
rect 5141 3261 5179 3295
rect 5179 3261 5213 3295
rect 5213 3261 5214 3295
rect 5034 3222 5214 3261
rect 5034 3188 5035 3222
rect 5035 3188 5069 3222
rect 5069 3188 5107 3222
rect 5107 3188 5141 3222
rect 5141 3188 5179 3222
rect 5179 3188 5213 3222
rect 5213 3188 5214 3222
rect 5034 3149 5214 3188
rect 5034 3115 5035 3149
rect 5035 3115 5069 3149
rect 5069 3115 5107 3149
rect 5107 3115 5141 3149
rect 5141 3115 5179 3149
rect 5179 3115 5213 3149
rect 5213 3115 5214 3149
rect 5034 3076 5214 3115
rect 5034 3042 5035 3076
rect 5035 3042 5069 3076
rect 5069 3042 5107 3076
rect 5107 3042 5141 3076
rect 5141 3042 5179 3076
rect 5179 3042 5213 3076
rect 5213 3042 5214 3076
rect 5034 3003 5214 3042
rect 5034 2969 5035 3003
rect 5035 2969 5069 3003
rect 5069 2969 5107 3003
rect 5107 2969 5141 3003
rect 5141 2969 5179 3003
rect 5179 2969 5213 3003
rect 5213 2969 5214 3003
rect 5034 2930 5214 2969
rect 5034 2896 5035 2930
rect 5035 2896 5069 2930
rect 5069 2896 5107 2930
rect 5107 2896 5141 2930
rect 5141 2896 5179 2930
rect 5179 2896 5213 2930
rect 5213 2896 5214 2930
rect 5034 2857 5214 2896
rect 5034 2823 5035 2857
rect 5035 2823 5069 2857
rect 5069 2823 5107 2857
rect 5107 2823 5141 2857
rect 5141 2823 5179 2857
rect 5179 2823 5213 2857
rect 5213 2823 5214 2857
rect 5034 2784 5214 2823
rect 5034 2750 5035 2784
rect 5035 2750 5069 2784
rect 5069 2750 5107 2784
rect 5107 2750 5141 2784
rect 5141 2750 5179 2784
rect 5179 2750 5213 2784
rect 5213 2750 5214 2784
rect 5034 2711 5214 2750
rect 5034 2677 5035 2711
rect 5035 2677 5069 2711
rect 5069 2677 5107 2711
rect 5107 2677 5141 2711
rect 5141 2677 5179 2711
rect 5179 2677 5213 2711
rect 5213 2677 5214 2711
rect 5034 2638 5214 2677
rect 5034 2604 5035 2638
rect 5035 2604 5069 2638
rect 5069 2604 5107 2638
rect 5107 2604 5141 2638
rect 5141 2604 5179 2638
rect 5179 2604 5213 2638
rect 5213 2604 5214 2638
rect 5034 2565 5214 2604
rect 5034 2531 5035 2565
rect 5035 2531 5069 2565
rect 5069 2531 5107 2565
rect 5107 2531 5141 2565
rect 5141 2531 5179 2565
rect 5179 2531 5213 2565
rect 5213 2531 5214 2565
rect 5034 2492 5214 2531
rect 5034 2458 5035 2492
rect 5035 2458 5069 2492
rect 5069 2458 5107 2492
rect 5107 2458 5141 2492
rect 5141 2458 5179 2492
rect 5179 2458 5213 2492
rect 5213 2458 5214 2492
rect 5034 2419 5214 2458
rect 5034 2385 5035 2419
rect 5035 2385 5069 2419
rect 5069 2385 5107 2419
rect 5107 2385 5141 2419
rect 5141 2385 5179 2419
rect 5179 2385 5213 2419
rect 5213 2385 5214 2419
rect 5034 2346 5214 2385
rect 5034 2312 5035 2346
rect 5035 2312 5069 2346
rect 5069 2312 5107 2346
rect 5107 2312 5141 2346
rect 5141 2312 5179 2346
rect 5179 2312 5213 2346
rect 5213 2312 5214 2346
rect 5034 2273 5214 2312
rect 5034 2239 5035 2273
rect 5035 2239 5069 2273
rect 5069 2239 5107 2273
rect 5107 2239 5141 2273
rect 5141 2239 5179 2273
rect 5179 2239 5213 2273
rect 5213 2239 5214 2273
rect 5034 2200 5214 2239
rect 5034 2166 5035 2200
rect 5035 2166 5069 2200
rect 5069 2166 5107 2200
rect 5107 2166 5141 2200
rect 5141 2166 5179 2200
rect 5179 2166 5213 2200
rect 5213 2166 5214 2200
rect 5034 2126 5214 2166
rect 5034 2092 5035 2126
rect 5035 2092 5069 2126
rect 5069 2092 5107 2126
rect 5107 2092 5141 2126
rect 5141 2092 5179 2126
rect 5179 2092 5213 2126
rect 5213 2092 5214 2126
rect 5034 2052 5214 2092
rect 5034 2018 5035 2052
rect 5035 2018 5069 2052
rect 5069 2018 5107 2052
rect 5107 2018 5141 2052
rect 5141 2018 5179 2052
rect 5179 2018 5213 2052
rect 5213 2018 5214 2052
rect 5034 1978 5214 2018
rect 5034 1944 5035 1978
rect 5035 1944 5069 1978
rect 5069 1944 5107 1978
rect 5107 1944 5141 1978
rect 5141 1944 5179 1978
rect 5179 1944 5213 1978
rect 5213 1944 5214 1978
rect 5034 1904 5214 1944
rect 5034 1870 5035 1904
rect 5035 1870 5069 1904
rect 5069 1870 5107 1904
rect 5107 1870 5141 1904
rect 5141 1870 5179 1904
rect 5179 1870 5213 1904
rect 5213 1870 5214 1904
rect 5034 1830 5214 1870
rect 5034 1796 5035 1830
rect 5035 1796 5069 1830
rect 5069 1796 5107 1830
rect 5107 1796 5141 1830
rect 5141 1796 5179 1830
rect 5179 1796 5213 1830
rect 5213 1796 5214 1830
rect 5034 1756 5214 1796
rect 5034 1722 5035 1756
rect 5035 1722 5069 1756
rect 5069 1722 5107 1756
rect 5107 1722 5141 1756
rect 5141 1722 5179 1756
rect 5179 1722 5213 1756
rect 5213 1722 5214 1756
rect 5034 1682 5214 1722
rect 5034 1648 5035 1682
rect 5035 1648 5069 1682
rect 5069 1648 5107 1682
rect 5107 1648 5141 1682
rect 5141 1648 5179 1682
rect 5179 1648 5213 1682
rect 5213 1648 5214 1682
rect 5034 1608 5214 1648
rect 5034 1574 5035 1608
rect 5035 1574 5069 1608
rect 5069 1574 5107 1608
rect 5107 1574 5141 1608
rect 5141 1574 5179 1608
rect 5179 1574 5213 1608
rect 5213 1574 5214 1608
rect 5034 1568 5214 1574
rect 5530 4092 5582 4124
rect 5594 4118 5646 4124
rect 5594 4092 5603 4118
rect 5603 4092 5637 4118
rect 5637 4092 5646 4118
rect 5658 4092 5710 4124
rect 5530 4072 5531 4092
rect 5531 4072 5582 4092
rect 5594 4072 5646 4092
rect 5658 4072 5709 4092
rect 5709 4072 5710 4092
rect 5530 4007 5531 4059
rect 5531 4007 5582 4059
rect 5594 4007 5646 4059
rect 5658 4007 5709 4059
rect 5709 4007 5710 4059
rect 5530 3942 5531 3994
rect 5531 3942 5582 3994
rect 5594 3942 5646 3994
rect 5658 3942 5709 3994
rect 5709 3942 5710 3994
rect 5530 3877 5531 3929
rect 5531 3877 5582 3929
rect 5594 3877 5646 3929
rect 5658 3877 5709 3929
rect 5709 3877 5710 3929
rect 5530 3812 5531 3864
rect 5531 3812 5582 3864
rect 5594 3812 5646 3864
rect 5658 3812 5709 3864
rect 5709 3812 5710 3864
rect 5530 3747 5531 3799
rect 5531 3747 5582 3799
rect 5594 3747 5646 3799
rect 5658 3747 5709 3799
rect 5709 3747 5710 3799
rect 5530 3682 5531 3734
rect 5531 3682 5582 3734
rect 5594 3682 5646 3734
rect 5658 3682 5709 3734
rect 5709 3682 5710 3734
rect 5530 3617 5531 3669
rect 5531 3617 5582 3669
rect 5594 3617 5646 3669
rect 5658 3617 5709 3669
rect 5709 3617 5710 3669
rect 5530 3194 5531 3604
rect 5531 3194 5709 3604
rect 5709 3194 5710 3604
rect 5530 3182 5710 3194
rect 5530 3148 5603 3182
rect 5603 3148 5637 3182
rect 5637 3148 5710 3182
rect 5530 3108 5710 3148
rect 5530 3074 5531 3108
rect 5531 3074 5565 3108
rect 5565 3074 5603 3108
rect 5603 3074 5637 3108
rect 5637 3074 5675 3108
rect 5675 3074 5709 3108
rect 5709 3074 5710 3108
rect 5530 3028 5710 3074
rect 5530 2994 5531 3028
rect 5531 2994 5565 3028
rect 5565 2994 5603 3028
rect 5603 2994 5637 3028
rect 5637 2994 5675 3028
rect 5675 2994 5709 3028
rect 5709 2994 5710 3028
rect 5530 2948 5710 2994
rect 5530 2914 5531 2948
rect 5531 2914 5565 2948
rect 5565 2914 5603 2948
rect 5603 2914 5637 2948
rect 5637 2914 5675 2948
rect 5675 2914 5709 2948
rect 5709 2914 5710 2948
rect 5530 2868 5710 2914
rect 5530 2834 5531 2868
rect 5531 2834 5565 2868
rect 5565 2834 5603 2868
rect 5603 2834 5637 2868
rect 5637 2834 5675 2868
rect 5675 2834 5709 2868
rect 5709 2834 5710 2868
rect 5530 2788 5710 2834
rect 5530 2754 5531 2788
rect 5531 2754 5565 2788
rect 5565 2754 5603 2788
rect 5603 2754 5637 2788
rect 5637 2754 5675 2788
rect 5675 2754 5709 2788
rect 5709 2754 5710 2788
rect 5530 2708 5710 2754
rect 5530 2674 5531 2708
rect 5531 2674 5565 2708
rect 5565 2674 5603 2708
rect 5603 2674 5637 2708
rect 5637 2674 5675 2708
rect 5675 2674 5709 2708
rect 5709 2674 5710 2708
rect 5530 2628 5710 2674
rect 5530 2594 5531 2628
rect 5531 2594 5565 2628
rect 5565 2594 5603 2628
rect 5603 2594 5637 2628
rect 5637 2594 5675 2628
rect 5675 2594 5709 2628
rect 5709 2594 5710 2628
rect 5530 2556 5710 2594
rect 5530 2522 5603 2556
rect 5603 2522 5637 2556
rect 5637 2522 5710 2556
rect 5530 2518 5710 2522
rect 5530 1620 5531 2518
rect 5531 1620 5709 2518
rect 5709 1620 5710 2518
rect 5530 1586 5603 1620
rect 5603 1586 5637 1620
rect 5637 1586 5710 1620
rect 5530 1568 5710 1586
rect 6026 4098 6078 4119
rect 6026 4067 6027 4098
rect 6027 4067 6061 4098
rect 6061 4067 6078 4098
rect 6090 4098 6142 4119
rect 6090 4067 6099 4098
rect 6099 4067 6133 4098
rect 6133 4067 6142 4098
rect 6154 4098 6206 4119
rect 6154 4067 6171 4098
rect 6171 4067 6205 4098
rect 6205 4067 6206 4098
rect 6026 4025 6078 4054
rect 6026 4002 6027 4025
rect 6027 4002 6061 4025
rect 6061 4002 6078 4025
rect 6090 4025 6142 4054
rect 6090 4002 6099 4025
rect 6099 4002 6133 4025
rect 6133 4002 6142 4025
rect 6154 4025 6206 4054
rect 6154 4002 6171 4025
rect 6171 4002 6205 4025
rect 6205 4002 6206 4025
rect 6026 3952 6078 3989
rect 6026 3937 6027 3952
rect 6027 3937 6061 3952
rect 6061 3937 6078 3952
rect 6090 3952 6142 3989
rect 6090 3937 6099 3952
rect 6099 3937 6133 3952
rect 6133 3937 6142 3952
rect 6154 3952 6206 3989
rect 6154 3937 6171 3952
rect 6171 3937 6205 3952
rect 6205 3937 6206 3952
rect 6026 3918 6027 3924
rect 6027 3918 6061 3924
rect 6061 3918 6099 3924
rect 6099 3918 6133 3924
rect 6133 3918 6171 3924
rect 6171 3918 6205 3924
rect 6205 3918 6206 3924
rect 6026 3879 6206 3918
rect 6026 3845 6027 3879
rect 6027 3845 6061 3879
rect 6061 3845 6099 3879
rect 6099 3845 6133 3879
rect 6133 3845 6171 3879
rect 6171 3845 6205 3879
rect 6205 3845 6206 3879
rect 6026 3806 6206 3845
rect 6026 3772 6027 3806
rect 6027 3772 6061 3806
rect 6061 3772 6099 3806
rect 6099 3772 6133 3806
rect 6133 3772 6171 3806
rect 6171 3772 6205 3806
rect 6205 3772 6206 3806
rect 6026 3733 6206 3772
rect 6026 3699 6027 3733
rect 6027 3699 6061 3733
rect 6061 3699 6099 3733
rect 6099 3699 6133 3733
rect 6133 3699 6171 3733
rect 6171 3699 6205 3733
rect 6205 3699 6206 3733
rect 6026 3660 6206 3699
rect 6026 3626 6027 3660
rect 6027 3626 6061 3660
rect 6061 3626 6099 3660
rect 6099 3626 6133 3660
rect 6133 3626 6171 3660
rect 6171 3626 6205 3660
rect 6205 3626 6206 3660
rect 6026 3587 6206 3626
rect 6026 3553 6027 3587
rect 6027 3553 6061 3587
rect 6061 3553 6099 3587
rect 6099 3553 6133 3587
rect 6133 3553 6171 3587
rect 6171 3553 6205 3587
rect 6205 3553 6206 3587
rect 6026 3514 6206 3553
rect 6026 3480 6027 3514
rect 6027 3480 6061 3514
rect 6061 3480 6099 3514
rect 6099 3480 6133 3514
rect 6133 3480 6171 3514
rect 6171 3480 6205 3514
rect 6205 3480 6206 3514
rect 6026 3441 6206 3480
rect 6026 3407 6027 3441
rect 6027 3407 6061 3441
rect 6061 3407 6099 3441
rect 6099 3407 6133 3441
rect 6133 3407 6171 3441
rect 6171 3407 6205 3441
rect 6205 3407 6206 3441
rect 6026 3368 6206 3407
rect 6026 3334 6027 3368
rect 6027 3334 6061 3368
rect 6061 3334 6099 3368
rect 6099 3334 6133 3368
rect 6133 3334 6171 3368
rect 6171 3334 6205 3368
rect 6205 3334 6206 3368
rect 6026 3295 6206 3334
rect 6026 3261 6027 3295
rect 6027 3261 6061 3295
rect 6061 3261 6099 3295
rect 6099 3261 6133 3295
rect 6133 3261 6171 3295
rect 6171 3261 6205 3295
rect 6205 3261 6206 3295
rect 6026 3222 6206 3261
rect 6026 3188 6027 3222
rect 6027 3188 6061 3222
rect 6061 3188 6099 3222
rect 6099 3188 6133 3222
rect 6133 3188 6171 3222
rect 6171 3188 6205 3222
rect 6205 3188 6206 3222
rect 6026 3149 6206 3188
rect 6026 3115 6027 3149
rect 6027 3115 6061 3149
rect 6061 3115 6099 3149
rect 6099 3115 6133 3149
rect 6133 3115 6171 3149
rect 6171 3115 6205 3149
rect 6205 3115 6206 3149
rect 6026 3076 6206 3115
rect 6026 3042 6027 3076
rect 6027 3042 6061 3076
rect 6061 3042 6099 3076
rect 6099 3042 6133 3076
rect 6133 3042 6171 3076
rect 6171 3042 6205 3076
rect 6205 3042 6206 3076
rect 6026 3003 6206 3042
rect 6026 2969 6027 3003
rect 6027 2969 6061 3003
rect 6061 2969 6099 3003
rect 6099 2969 6133 3003
rect 6133 2969 6171 3003
rect 6171 2969 6205 3003
rect 6205 2969 6206 3003
rect 6026 2930 6206 2969
rect 6026 2896 6027 2930
rect 6027 2896 6061 2930
rect 6061 2896 6099 2930
rect 6099 2896 6133 2930
rect 6133 2896 6171 2930
rect 6171 2896 6205 2930
rect 6205 2896 6206 2930
rect 6026 2857 6206 2896
rect 6026 2823 6027 2857
rect 6027 2823 6061 2857
rect 6061 2823 6099 2857
rect 6099 2823 6133 2857
rect 6133 2823 6171 2857
rect 6171 2823 6205 2857
rect 6205 2823 6206 2857
rect 6026 2784 6206 2823
rect 6026 2750 6027 2784
rect 6027 2750 6061 2784
rect 6061 2750 6099 2784
rect 6099 2750 6133 2784
rect 6133 2750 6171 2784
rect 6171 2750 6205 2784
rect 6205 2750 6206 2784
rect 6026 2711 6206 2750
rect 6026 2677 6027 2711
rect 6027 2677 6061 2711
rect 6061 2677 6099 2711
rect 6099 2677 6133 2711
rect 6133 2677 6171 2711
rect 6171 2677 6205 2711
rect 6205 2677 6206 2711
rect 6026 2638 6206 2677
rect 6026 2604 6027 2638
rect 6027 2604 6061 2638
rect 6061 2604 6099 2638
rect 6099 2604 6133 2638
rect 6133 2604 6171 2638
rect 6171 2604 6205 2638
rect 6205 2604 6206 2638
rect 6026 2565 6206 2604
rect 6026 2531 6027 2565
rect 6027 2531 6061 2565
rect 6061 2531 6099 2565
rect 6099 2531 6133 2565
rect 6133 2531 6171 2565
rect 6171 2531 6205 2565
rect 6205 2531 6206 2565
rect 6026 2492 6206 2531
rect 6026 2458 6027 2492
rect 6027 2458 6061 2492
rect 6061 2458 6099 2492
rect 6099 2458 6133 2492
rect 6133 2458 6171 2492
rect 6171 2458 6205 2492
rect 6205 2458 6206 2492
rect 6026 2419 6206 2458
rect 6026 2385 6027 2419
rect 6027 2385 6061 2419
rect 6061 2385 6099 2419
rect 6099 2385 6133 2419
rect 6133 2385 6171 2419
rect 6171 2385 6205 2419
rect 6205 2385 6206 2419
rect 6026 2346 6206 2385
rect 6026 2312 6027 2346
rect 6027 2312 6061 2346
rect 6061 2312 6099 2346
rect 6099 2312 6133 2346
rect 6133 2312 6171 2346
rect 6171 2312 6205 2346
rect 6205 2312 6206 2346
rect 6026 2273 6206 2312
rect 6026 2239 6027 2273
rect 6027 2239 6061 2273
rect 6061 2239 6099 2273
rect 6099 2239 6133 2273
rect 6133 2239 6171 2273
rect 6171 2239 6205 2273
rect 6205 2239 6206 2273
rect 6026 2200 6206 2239
rect 6026 2166 6027 2200
rect 6027 2166 6061 2200
rect 6061 2166 6099 2200
rect 6099 2166 6133 2200
rect 6133 2166 6171 2200
rect 6171 2166 6205 2200
rect 6205 2166 6206 2200
rect 6026 2126 6206 2166
rect 6026 2092 6027 2126
rect 6027 2092 6061 2126
rect 6061 2092 6099 2126
rect 6099 2092 6133 2126
rect 6133 2092 6171 2126
rect 6171 2092 6205 2126
rect 6205 2092 6206 2126
rect 6026 2052 6206 2092
rect 6026 2018 6027 2052
rect 6027 2018 6061 2052
rect 6061 2018 6099 2052
rect 6099 2018 6133 2052
rect 6133 2018 6171 2052
rect 6171 2018 6205 2052
rect 6205 2018 6206 2052
rect 6026 1978 6206 2018
rect 6026 1944 6027 1978
rect 6027 1944 6061 1978
rect 6061 1944 6099 1978
rect 6099 1944 6133 1978
rect 6133 1944 6171 1978
rect 6171 1944 6205 1978
rect 6205 1944 6206 1978
rect 6026 1904 6206 1944
rect 6026 1870 6027 1904
rect 6027 1870 6061 1904
rect 6061 1870 6099 1904
rect 6099 1870 6133 1904
rect 6133 1870 6171 1904
rect 6171 1870 6205 1904
rect 6205 1870 6206 1904
rect 6026 1830 6206 1870
rect 6026 1796 6027 1830
rect 6027 1796 6061 1830
rect 6061 1796 6099 1830
rect 6099 1796 6133 1830
rect 6133 1796 6171 1830
rect 6171 1796 6205 1830
rect 6205 1796 6206 1830
rect 6026 1756 6206 1796
rect 6026 1722 6027 1756
rect 6027 1722 6061 1756
rect 6061 1722 6099 1756
rect 6099 1722 6133 1756
rect 6133 1722 6171 1756
rect 6171 1722 6205 1756
rect 6205 1722 6206 1756
rect 6026 1682 6206 1722
rect 6026 1648 6027 1682
rect 6027 1648 6061 1682
rect 6061 1648 6099 1682
rect 6099 1648 6133 1682
rect 6133 1648 6171 1682
rect 6171 1648 6205 1682
rect 6205 1648 6206 1682
rect 6026 1608 6206 1648
rect 6026 1574 6027 1608
rect 6027 1574 6061 1608
rect 6061 1574 6099 1608
rect 6099 1574 6133 1608
rect 6133 1574 6171 1608
rect 6171 1574 6205 1608
rect 6205 1574 6206 1608
rect 6026 1568 6206 1574
rect 6522 4092 6574 4124
rect 6586 4118 6638 4124
rect 6586 4092 6595 4118
rect 6595 4092 6629 4118
rect 6629 4092 6638 4118
rect 6650 4092 6702 4124
rect 6522 4072 6523 4092
rect 6523 4072 6574 4092
rect 6586 4072 6638 4092
rect 6650 4072 6701 4092
rect 6701 4072 6702 4092
rect 6522 4007 6523 4059
rect 6523 4007 6574 4059
rect 6586 4007 6638 4059
rect 6650 4007 6701 4059
rect 6701 4007 6702 4059
rect 6522 3942 6523 3994
rect 6523 3942 6574 3994
rect 6586 3942 6638 3994
rect 6650 3942 6701 3994
rect 6701 3942 6702 3994
rect 6522 3877 6523 3929
rect 6523 3877 6574 3929
rect 6586 3877 6638 3929
rect 6650 3877 6701 3929
rect 6701 3877 6702 3929
rect 6522 3812 6523 3864
rect 6523 3812 6574 3864
rect 6586 3812 6638 3864
rect 6650 3812 6701 3864
rect 6701 3812 6702 3864
rect 6522 3747 6523 3799
rect 6523 3747 6574 3799
rect 6586 3747 6638 3799
rect 6650 3747 6701 3799
rect 6701 3747 6702 3799
rect 6522 3682 6523 3734
rect 6523 3682 6574 3734
rect 6586 3682 6638 3734
rect 6650 3682 6701 3734
rect 6701 3682 6702 3734
rect 6522 3617 6523 3669
rect 6523 3617 6574 3669
rect 6586 3617 6638 3669
rect 6650 3617 6701 3669
rect 6701 3617 6702 3669
rect 6522 3194 6523 3604
rect 6523 3194 6701 3604
rect 6701 3194 6702 3604
rect 6522 3182 6702 3194
rect 6522 3148 6595 3182
rect 6595 3148 6629 3182
rect 6629 3148 6702 3182
rect 6522 3108 6702 3148
rect 6522 3074 6523 3108
rect 6523 3074 6557 3108
rect 6557 3074 6595 3108
rect 6595 3074 6629 3108
rect 6629 3074 6667 3108
rect 6667 3074 6701 3108
rect 6701 3074 6702 3108
rect 6522 3028 6702 3074
rect 6522 2994 6523 3028
rect 6523 2994 6557 3028
rect 6557 2994 6595 3028
rect 6595 2994 6629 3028
rect 6629 2994 6667 3028
rect 6667 2994 6701 3028
rect 6701 2994 6702 3028
rect 6522 2948 6702 2994
rect 6522 2914 6523 2948
rect 6523 2914 6557 2948
rect 6557 2914 6595 2948
rect 6595 2914 6629 2948
rect 6629 2914 6667 2948
rect 6667 2914 6701 2948
rect 6701 2914 6702 2948
rect 6522 2868 6702 2914
rect 6522 2834 6523 2868
rect 6523 2834 6557 2868
rect 6557 2834 6595 2868
rect 6595 2834 6629 2868
rect 6629 2834 6667 2868
rect 6667 2834 6701 2868
rect 6701 2834 6702 2868
rect 6522 2788 6702 2834
rect 6522 2754 6523 2788
rect 6523 2754 6557 2788
rect 6557 2754 6595 2788
rect 6595 2754 6629 2788
rect 6629 2754 6667 2788
rect 6667 2754 6701 2788
rect 6701 2754 6702 2788
rect 6522 2708 6702 2754
rect 6522 2674 6523 2708
rect 6523 2674 6557 2708
rect 6557 2674 6595 2708
rect 6595 2674 6629 2708
rect 6629 2674 6667 2708
rect 6667 2674 6701 2708
rect 6701 2674 6702 2708
rect 6522 2628 6702 2674
rect 6522 2594 6523 2628
rect 6523 2594 6557 2628
rect 6557 2594 6595 2628
rect 6595 2594 6629 2628
rect 6629 2594 6667 2628
rect 6667 2594 6701 2628
rect 6701 2594 6702 2628
rect 6522 2556 6702 2594
rect 6522 2522 6595 2556
rect 6595 2522 6629 2556
rect 6629 2522 6702 2556
rect 6522 2518 6702 2522
rect 6522 1620 6523 2518
rect 6523 1620 6701 2518
rect 6701 1620 6702 2518
rect 6522 1586 6595 1620
rect 6595 1586 6629 1620
rect 6629 1586 6702 1620
rect 6522 1568 6702 1586
rect 7018 4098 7070 4119
rect 7018 4067 7019 4098
rect 7019 4067 7053 4098
rect 7053 4067 7070 4098
rect 7082 4098 7134 4119
rect 7082 4067 7091 4098
rect 7091 4067 7125 4098
rect 7125 4067 7134 4098
rect 7146 4098 7198 4119
rect 7146 4067 7163 4098
rect 7163 4067 7197 4098
rect 7197 4067 7198 4098
rect 7018 4025 7070 4054
rect 7018 4002 7019 4025
rect 7019 4002 7053 4025
rect 7053 4002 7070 4025
rect 7082 4025 7134 4054
rect 7082 4002 7091 4025
rect 7091 4002 7125 4025
rect 7125 4002 7134 4025
rect 7146 4025 7198 4054
rect 7146 4002 7163 4025
rect 7163 4002 7197 4025
rect 7197 4002 7198 4025
rect 7018 3952 7070 3989
rect 7018 3937 7019 3952
rect 7019 3937 7053 3952
rect 7053 3937 7070 3952
rect 7082 3952 7134 3989
rect 7082 3937 7091 3952
rect 7091 3937 7125 3952
rect 7125 3937 7134 3952
rect 7146 3952 7198 3989
rect 7146 3937 7163 3952
rect 7163 3937 7197 3952
rect 7197 3937 7198 3952
rect 7018 3918 7019 3924
rect 7019 3918 7053 3924
rect 7053 3918 7091 3924
rect 7091 3918 7125 3924
rect 7125 3918 7163 3924
rect 7163 3918 7197 3924
rect 7197 3918 7198 3924
rect 7018 3879 7198 3918
rect 7018 3845 7019 3879
rect 7019 3845 7053 3879
rect 7053 3845 7091 3879
rect 7091 3845 7125 3879
rect 7125 3845 7163 3879
rect 7163 3845 7197 3879
rect 7197 3845 7198 3879
rect 7018 3806 7198 3845
rect 7018 3772 7019 3806
rect 7019 3772 7053 3806
rect 7053 3772 7091 3806
rect 7091 3772 7125 3806
rect 7125 3772 7163 3806
rect 7163 3772 7197 3806
rect 7197 3772 7198 3806
rect 7018 3733 7198 3772
rect 7018 3699 7019 3733
rect 7019 3699 7053 3733
rect 7053 3699 7091 3733
rect 7091 3699 7125 3733
rect 7125 3699 7163 3733
rect 7163 3699 7197 3733
rect 7197 3699 7198 3733
rect 7018 3660 7198 3699
rect 7018 3626 7019 3660
rect 7019 3626 7053 3660
rect 7053 3626 7091 3660
rect 7091 3626 7125 3660
rect 7125 3626 7163 3660
rect 7163 3626 7197 3660
rect 7197 3626 7198 3660
rect 7018 3587 7198 3626
rect 7018 3553 7019 3587
rect 7019 3553 7053 3587
rect 7053 3553 7091 3587
rect 7091 3553 7125 3587
rect 7125 3553 7163 3587
rect 7163 3553 7197 3587
rect 7197 3553 7198 3587
rect 7018 3514 7198 3553
rect 7018 3480 7019 3514
rect 7019 3480 7053 3514
rect 7053 3480 7091 3514
rect 7091 3480 7125 3514
rect 7125 3480 7163 3514
rect 7163 3480 7197 3514
rect 7197 3480 7198 3514
rect 7018 3441 7198 3480
rect 7018 3407 7019 3441
rect 7019 3407 7053 3441
rect 7053 3407 7091 3441
rect 7091 3407 7125 3441
rect 7125 3407 7163 3441
rect 7163 3407 7197 3441
rect 7197 3407 7198 3441
rect 7018 3368 7198 3407
rect 7018 3334 7019 3368
rect 7019 3334 7053 3368
rect 7053 3334 7091 3368
rect 7091 3334 7125 3368
rect 7125 3334 7163 3368
rect 7163 3334 7197 3368
rect 7197 3334 7198 3368
rect 7018 3295 7198 3334
rect 7018 3261 7019 3295
rect 7019 3261 7053 3295
rect 7053 3261 7091 3295
rect 7091 3261 7125 3295
rect 7125 3261 7163 3295
rect 7163 3261 7197 3295
rect 7197 3261 7198 3295
rect 7018 3222 7198 3261
rect 7018 3188 7019 3222
rect 7019 3188 7053 3222
rect 7053 3188 7091 3222
rect 7091 3188 7125 3222
rect 7125 3188 7163 3222
rect 7163 3188 7197 3222
rect 7197 3188 7198 3222
rect 7018 3149 7198 3188
rect 7018 3115 7019 3149
rect 7019 3115 7053 3149
rect 7053 3115 7091 3149
rect 7091 3115 7125 3149
rect 7125 3115 7163 3149
rect 7163 3115 7197 3149
rect 7197 3115 7198 3149
rect 7018 3076 7198 3115
rect 7018 3042 7019 3076
rect 7019 3042 7053 3076
rect 7053 3042 7091 3076
rect 7091 3042 7125 3076
rect 7125 3042 7163 3076
rect 7163 3042 7197 3076
rect 7197 3042 7198 3076
rect 7018 3003 7198 3042
rect 7018 2969 7019 3003
rect 7019 2969 7053 3003
rect 7053 2969 7091 3003
rect 7091 2969 7125 3003
rect 7125 2969 7163 3003
rect 7163 2969 7197 3003
rect 7197 2969 7198 3003
rect 7018 2930 7198 2969
rect 7018 2896 7019 2930
rect 7019 2896 7053 2930
rect 7053 2896 7091 2930
rect 7091 2896 7125 2930
rect 7125 2896 7163 2930
rect 7163 2896 7197 2930
rect 7197 2896 7198 2930
rect 7018 2857 7198 2896
rect 7018 2823 7019 2857
rect 7019 2823 7053 2857
rect 7053 2823 7091 2857
rect 7091 2823 7125 2857
rect 7125 2823 7163 2857
rect 7163 2823 7197 2857
rect 7197 2823 7198 2857
rect 7018 2784 7198 2823
rect 7018 2750 7019 2784
rect 7019 2750 7053 2784
rect 7053 2750 7091 2784
rect 7091 2750 7125 2784
rect 7125 2750 7163 2784
rect 7163 2750 7197 2784
rect 7197 2750 7198 2784
rect 7018 2711 7198 2750
rect 7018 2677 7019 2711
rect 7019 2677 7053 2711
rect 7053 2677 7091 2711
rect 7091 2677 7125 2711
rect 7125 2677 7163 2711
rect 7163 2677 7197 2711
rect 7197 2677 7198 2711
rect 7018 2638 7198 2677
rect 7018 2604 7019 2638
rect 7019 2604 7053 2638
rect 7053 2604 7091 2638
rect 7091 2604 7125 2638
rect 7125 2604 7163 2638
rect 7163 2604 7197 2638
rect 7197 2604 7198 2638
rect 7018 2565 7198 2604
rect 7018 2531 7019 2565
rect 7019 2531 7053 2565
rect 7053 2531 7091 2565
rect 7091 2531 7125 2565
rect 7125 2531 7163 2565
rect 7163 2531 7197 2565
rect 7197 2531 7198 2565
rect 7018 2492 7198 2531
rect 7018 2458 7019 2492
rect 7019 2458 7053 2492
rect 7053 2458 7091 2492
rect 7091 2458 7125 2492
rect 7125 2458 7163 2492
rect 7163 2458 7197 2492
rect 7197 2458 7198 2492
rect 7018 2419 7198 2458
rect 7018 2385 7019 2419
rect 7019 2385 7053 2419
rect 7053 2385 7091 2419
rect 7091 2385 7125 2419
rect 7125 2385 7163 2419
rect 7163 2385 7197 2419
rect 7197 2385 7198 2419
rect 7018 2346 7198 2385
rect 7018 2312 7019 2346
rect 7019 2312 7053 2346
rect 7053 2312 7091 2346
rect 7091 2312 7125 2346
rect 7125 2312 7163 2346
rect 7163 2312 7197 2346
rect 7197 2312 7198 2346
rect 7018 2273 7198 2312
rect 7018 2239 7019 2273
rect 7019 2239 7053 2273
rect 7053 2239 7091 2273
rect 7091 2239 7125 2273
rect 7125 2239 7163 2273
rect 7163 2239 7197 2273
rect 7197 2239 7198 2273
rect 7018 2200 7198 2239
rect 7018 2166 7019 2200
rect 7019 2166 7053 2200
rect 7053 2166 7091 2200
rect 7091 2166 7125 2200
rect 7125 2166 7163 2200
rect 7163 2166 7197 2200
rect 7197 2166 7198 2200
rect 7018 2126 7198 2166
rect 7018 2092 7019 2126
rect 7019 2092 7053 2126
rect 7053 2092 7091 2126
rect 7091 2092 7125 2126
rect 7125 2092 7163 2126
rect 7163 2092 7197 2126
rect 7197 2092 7198 2126
rect 7018 2052 7198 2092
rect 7018 2018 7019 2052
rect 7019 2018 7053 2052
rect 7053 2018 7091 2052
rect 7091 2018 7125 2052
rect 7125 2018 7163 2052
rect 7163 2018 7197 2052
rect 7197 2018 7198 2052
rect 7018 1978 7198 2018
rect 7018 1944 7019 1978
rect 7019 1944 7053 1978
rect 7053 1944 7091 1978
rect 7091 1944 7125 1978
rect 7125 1944 7163 1978
rect 7163 1944 7197 1978
rect 7197 1944 7198 1978
rect 7018 1904 7198 1944
rect 7018 1870 7019 1904
rect 7019 1870 7053 1904
rect 7053 1870 7091 1904
rect 7091 1870 7125 1904
rect 7125 1870 7163 1904
rect 7163 1870 7197 1904
rect 7197 1870 7198 1904
rect 7018 1830 7198 1870
rect 7018 1796 7019 1830
rect 7019 1796 7053 1830
rect 7053 1796 7091 1830
rect 7091 1796 7125 1830
rect 7125 1796 7163 1830
rect 7163 1796 7197 1830
rect 7197 1796 7198 1830
rect 7018 1756 7198 1796
rect 7018 1722 7019 1756
rect 7019 1722 7053 1756
rect 7053 1722 7091 1756
rect 7091 1722 7125 1756
rect 7125 1722 7163 1756
rect 7163 1722 7197 1756
rect 7197 1722 7198 1756
rect 7018 1682 7198 1722
rect 7018 1648 7019 1682
rect 7019 1648 7053 1682
rect 7053 1648 7091 1682
rect 7091 1648 7125 1682
rect 7125 1648 7163 1682
rect 7163 1648 7197 1682
rect 7197 1648 7198 1682
rect 7018 1608 7198 1648
rect 7018 1574 7019 1608
rect 7019 1574 7053 1608
rect 7053 1574 7091 1608
rect 7091 1574 7125 1608
rect 7125 1574 7163 1608
rect 7163 1574 7197 1608
rect 7197 1574 7198 1608
rect 7018 1568 7198 1574
rect 7514 4092 7566 4124
rect 7578 4118 7630 4124
rect 7578 4092 7587 4118
rect 7587 4092 7621 4118
rect 7621 4092 7630 4118
rect 7642 4092 7694 4124
rect 7514 4072 7515 4092
rect 7515 4072 7566 4092
rect 7578 4072 7630 4092
rect 7642 4072 7693 4092
rect 7693 4072 7694 4092
rect 7514 4007 7515 4059
rect 7515 4007 7566 4059
rect 7578 4007 7630 4059
rect 7642 4007 7693 4059
rect 7693 4007 7694 4059
rect 7514 3942 7515 3994
rect 7515 3942 7566 3994
rect 7578 3942 7630 3994
rect 7642 3942 7693 3994
rect 7693 3942 7694 3994
rect 7514 3877 7515 3929
rect 7515 3877 7566 3929
rect 7578 3877 7630 3929
rect 7642 3877 7693 3929
rect 7693 3877 7694 3929
rect 7514 3812 7515 3864
rect 7515 3812 7566 3864
rect 7578 3812 7630 3864
rect 7642 3812 7693 3864
rect 7693 3812 7694 3864
rect 7514 3747 7515 3799
rect 7515 3747 7566 3799
rect 7578 3747 7630 3799
rect 7642 3747 7693 3799
rect 7693 3747 7694 3799
rect 7514 3682 7515 3734
rect 7515 3682 7566 3734
rect 7578 3682 7630 3734
rect 7642 3682 7693 3734
rect 7693 3682 7694 3734
rect 7514 3617 7515 3669
rect 7515 3617 7566 3669
rect 7578 3617 7630 3669
rect 7642 3617 7693 3669
rect 7693 3617 7694 3669
rect 7514 3194 7515 3604
rect 7515 3194 7693 3604
rect 7693 3194 7694 3604
rect 7514 3182 7694 3194
rect 7514 3148 7587 3182
rect 7587 3148 7621 3182
rect 7621 3148 7694 3182
rect 7514 3108 7694 3148
rect 7514 3074 7515 3108
rect 7515 3074 7549 3108
rect 7549 3074 7587 3108
rect 7587 3074 7621 3108
rect 7621 3074 7659 3108
rect 7659 3074 7693 3108
rect 7693 3074 7694 3108
rect 7514 3028 7694 3074
rect 7514 2994 7515 3028
rect 7515 2994 7549 3028
rect 7549 2994 7587 3028
rect 7587 2994 7621 3028
rect 7621 2994 7659 3028
rect 7659 2994 7693 3028
rect 7693 2994 7694 3028
rect 7514 2948 7694 2994
rect 7514 2914 7515 2948
rect 7515 2914 7549 2948
rect 7549 2914 7587 2948
rect 7587 2914 7621 2948
rect 7621 2914 7659 2948
rect 7659 2914 7693 2948
rect 7693 2914 7694 2948
rect 7514 2868 7694 2914
rect 7514 2834 7515 2868
rect 7515 2834 7549 2868
rect 7549 2834 7587 2868
rect 7587 2834 7621 2868
rect 7621 2834 7659 2868
rect 7659 2834 7693 2868
rect 7693 2834 7694 2868
rect 7514 2788 7694 2834
rect 7514 2754 7515 2788
rect 7515 2754 7549 2788
rect 7549 2754 7587 2788
rect 7587 2754 7621 2788
rect 7621 2754 7659 2788
rect 7659 2754 7693 2788
rect 7693 2754 7694 2788
rect 7514 2708 7694 2754
rect 7514 2674 7515 2708
rect 7515 2674 7549 2708
rect 7549 2674 7587 2708
rect 7587 2674 7621 2708
rect 7621 2674 7659 2708
rect 7659 2674 7693 2708
rect 7693 2674 7694 2708
rect 7514 2628 7694 2674
rect 7514 2594 7515 2628
rect 7515 2594 7549 2628
rect 7549 2594 7587 2628
rect 7587 2594 7621 2628
rect 7621 2594 7659 2628
rect 7659 2594 7693 2628
rect 7693 2594 7694 2628
rect 7514 2556 7694 2594
rect 7514 2522 7587 2556
rect 7587 2522 7621 2556
rect 7621 2522 7694 2556
rect 7514 2518 7694 2522
rect 7514 1620 7515 2518
rect 7515 1620 7693 2518
rect 7693 1620 7694 2518
rect 7514 1586 7587 1620
rect 7587 1586 7621 1620
rect 7621 1586 7694 1620
rect 7514 1568 7694 1586
rect 8010 4098 8062 4119
rect 8010 4067 8011 4098
rect 8011 4067 8045 4098
rect 8045 4067 8062 4098
rect 8074 4098 8126 4119
rect 8074 4067 8083 4098
rect 8083 4067 8117 4098
rect 8117 4067 8126 4098
rect 8138 4098 8190 4119
rect 8138 4067 8155 4098
rect 8155 4067 8189 4098
rect 8189 4067 8190 4098
rect 8010 4025 8062 4054
rect 8010 4002 8011 4025
rect 8011 4002 8045 4025
rect 8045 4002 8062 4025
rect 8074 4025 8126 4054
rect 8074 4002 8083 4025
rect 8083 4002 8117 4025
rect 8117 4002 8126 4025
rect 8138 4025 8190 4054
rect 8138 4002 8155 4025
rect 8155 4002 8189 4025
rect 8189 4002 8190 4025
rect 8010 3952 8062 3989
rect 8010 3937 8011 3952
rect 8011 3937 8045 3952
rect 8045 3937 8062 3952
rect 8074 3952 8126 3989
rect 8074 3937 8083 3952
rect 8083 3937 8117 3952
rect 8117 3937 8126 3952
rect 8138 3952 8190 3989
rect 8138 3937 8155 3952
rect 8155 3937 8189 3952
rect 8189 3937 8190 3952
rect 8010 3918 8011 3924
rect 8011 3918 8045 3924
rect 8045 3918 8083 3924
rect 8083 3918 8117 3924
rect 8117 3918 8155 3924
rect 8155 3918 8189 3924
rect 8189 3918 8190 3924
rect 8010 3879 8190 3918
rect 8010 3845 8011 3879
rect 8011 3845 8045 3879
rect 8045 3845 8083 3879
rect 8083 3845 8117 3879
rect 8117 3845 8155 3879
rect 8155 3845 8189 3879
rect 8189 3845 8190 3879
rect 8010 3806 8190 3845
rect 8010 3772 8011 3806
rect 8011 3772 8045 3806
rect 8045 3772 8083 3806
rect 8083 3772 8117 3806
rect 8117 3772 8155 3806
rect 8155 3772 8189 3806
rect 8189 3772 8190 3806
rect 8010 3733 8190 3772
rect 8010 3699 8011 3733
rect 8011 3699 8045 3733
rect 8045 3699 8083 3733
rect 8083 3699 8117 3733
rect 8117 3699 8155 3733
rect 8155 3699 8189 3733
rect 8189 3699 8190 3733
rect 8010 3660 8190 3699
rect 8010 3626 8011 3660
rect 8011 3626 8045 3660
rect 8045 3626 8083 3660
rect 8083 3626 8117 3660
rect 8117 3626 8155 3660
rect 8155 3626 8189 3660
rect 8189 3626 8190 3660
rect 8010 3587 8190 3626
rect 8010 3553 8011 3587
rect 8011 3553 8045 3587
rect 8045 3553 8083 3587
rect 8083 3553 8117 3587
rect 8117 3553 8155 3587
rect 8155 3553 8189 3587
rect 8189 3553 8190 3587
rect 8010 3514 8190 3553
rect 8010 3480 8011 3514
rect 8011 3480 8045 3514
rect 8045 3480 8083 3514
rect 8083 3480 8117 3514
rect 8117 3480 8155 3514
rect 8155 3480 8189 3514
rect 8189 3480 8190 3514
rect 8010 3441 8190 3480
rect 8010 3407 8011 3441
rect 8011 3407 8045 3441
rect 8045 3407 8083 3441
rect 8083 3407 8117 3441
rect 8117 3407 8155 3441
rect 8155 3407 8189 3441
rect 8189 3407 8190 3441
rect 8010 3368 8190 3407
rect 8010 3334 8011 3368
rect 8011 3334 8045 3368
rect 8045 3334 8083 3368
rect 8083 3334 8117 3368
rect 8117 3334 8155 3368
rect 8155 3334 8189 3368
rect 8189 3334 8190 3368
rect 8010 3295 8190 3334
rect 8010 3261 8011 3295
rect 8011 3261 8045 3295
rect 8045 3261 8083 3295
rect 8083 3261 8117 3295
rect 8117 3261 8155 3295
rect 8155 3261 8189 3295
rect 8189 3261 8190 3295
rect 8010 3222 8190 3261
rect 8010 3188 8011 3222
rect 8011 3188 8045 3222
rect 8045 3188 8083 3222
rect 8083 3188 8117 3222
rect 8117 3188 8155 3222
rect 8155 3188 8189 3222
rect 8189 3188 8190 3222
rect 8010 3149 8190 3188
rect 8010 3115 8011 3149
rect 8011 3115 8045 3149
rect 8045 3115 8083 3149
rect 8083 3115 8117 3149
rect 8117 3115 8155 3149
rect 8155 3115 8189 3149
rect 8189 3115 8190 3149
rect 8010 3076 8190 3115
rect 8010 3042 8011 3076
rect 8011 3042 8045 3076
rect 8045 3042 8083 3076
rect 8083 3042 8117 3076
rect 8117 3042 8155 3076
rect 8155 3042 8189 3076
rect 8189 3042 8190 3076
rect 8010 3003 8190 3042
rect 8010 2969 8011 3003
rect 8011 2969 8045 3003
rect 8045 2969 8083 3003
rect 8083 2969 8117 3003
rect 8117 2969 8155 3003
rect 8155 2969 8189 3003
rect 8189 2969 8190 3003
rect 8010 2930 8190 2969
rect 8010 2896 8011 2930
rect 8011 2896 8045 2930
rect 8045 2896 8083 2930
rect 8083 2896 8117 2930
rect 8117 2896 8155 2930
rect 8155 2896 8189 2930
rect 8189 2896 8190 2930
rect 8010 2857 8190 2896
rect 8010 2823 8011 2857
rect 8011 2823 8045 2857
rect 8045 2823 8083 2857
rect 8083 2823 8117 2857
rect 8117 2823 8155 2857
rect 8155 2823 8189 2857
rect 8189 2823 8190 2857
rect 8010 2784 8190 2823
rect 8010 2750 8011 2784
rect 8011 2750 8045 2784
rect 8045 2750 8083 2784
rect 8083 2750 8117 2784
rect 8117 2750 8155 2784
rect 8155 2750 8189 2784
rect 8189 2750 8190 2784
rect 8010 2711 8190 2750
rect 8010 2677 8011 2711
rect 8011 2677 8045 2711
rect 8045 2677 8083 2711
rect 8083 2677 8117 2711
rect 8117 2677 8155 2711
rect 8155 2677 8189 2711
rect 8189 2677 8190 2711
rect 8010 2638 8190 2677
rect 8010 2604 8011 2638
rect 8011 2604 8045 2638
rect 8045 2604 8083 2638
rect 8083 2604 8117 2638
rect 8117 2604 8155 2638
rect 8155 2604 8189 2638
rect 8189 2604 8190 2638
rect 8010 2565 8190 2604
rect 8010 2531 8011 2565
rect 8011 2531 8045 2565
rect 8045 2531 8083 2565
rect 8083 2531 8117 2565
rect 8117 2531 8155 2565
rect 8155 2531 8189 2565
rect 8189 2531 8190 2565
rect 8010 2492 8190 2531
rect 8010 2458 8011 2492
rect 8011 2458 8045 2492
rect 8045 2458 8083 2492
rect 8083 2458 8117 2492
rect 8117 2458 8155 2492
rect 8155 2458 8189 2492
rect 8189 2458 8190 2492
rect 8010 2419 8190 2458
rect 8010 2385 8011 2419
rect 8011 2385 8045 2419
rect 8045 2385 8083 2419
rect 8083 2385 8117 2419
rect 8117 2385 8155 2419
rect 8155 2385 8189 2419
rect 8189 2385 8190 2419
rect 8010 2346 8190 2385
rect 8010 2312 8011 2346
rect 8011 2312 8045 2346
rect 8045 2312 8083 2346
rect 8083 2312 8117 2346
rect 8117 2312 8155 2346
rect 8155 2312 8189 2346
rect 8189 2312 8190 2346
rect 8010 2273 8190 2312
rect 8010 2239 8011 2273
rect 8011 2239 8045 2273
rect 8045 2239 8083 2273
rect 8083 2239 8117 2273
rect 8117 2239 8155 2273
rect 8155 2239 8189 2273
rect 8189 2239 8190 2273
rect 8010 2200 8190 2239
rect 8010 2166 8011 2200
rect 8011 2166 8045 2200
rect 8045 2166 8083 2200
rect 8083 2166 8117 2200
rect 8117 2166 8155 2200
rect 8155 2166 8189 2200
rect 8189 2166 8190 2200
rect 8010 2126 8190 2166
rect 8010 2092 8011 2126
rect 8011 2092 8045 2126
rect 8045 2092 8083 2126
rect 8083 2092 8117 2126
rect 8117 2092 8155 2126
rect 8155 2092 8189 2126
rect 8189 2092 8190 2126
rect 8010 2052 8190 2092
rect 8010 2018 8011 2052
rect 8011 2018 8045 2052
rect 8045 2018 8083 2052
rect 8083 2018 8117 2052
rect 8117 2018 8155 2052
rect 8155 2018 8189 2052
rect 8189 2018 8190 2052
rect 8010 1978 8190 2018
rect 8010 1944 8011 1978
rect 8011 1944 8045 1978
rect 8045 1944 8083 1978
rect 8083 1944 8117 1978
rect 8117 1944 8155 1978
rect 8155 1944 8189 1978
rect 8189 1944 8190 1978
rect 8010 1904 8190 1944
rect 8010 1870 8011 1904
rect 8011 1870 8045 1904
rect 8045 1870 8083 1904
rect 8083 1870 8117 1904
rect 8117 1870 8155 1904
rect 8155 1870 8189 1904
rect 8189 1870 8190 1904
rect 8010 1830 8190 1870
rect 8010 1796 8011 1830
rect 8011 1796 8045 1830
rect 8045 1796 8083 1830
rect 8083 1796 8117 1830
rect 8117 1796 8155 1830
rect 8155 1796 8189 1830
rect 8189 1796 8190 1830
rect 8010 1756 8190 1796
rect 8010 1722 8011 1756
rect 8011 1722 8045 1756
rect 8045 1722 8083 1756
rect 8083 1722 8117 1756
rect 8117 1722 8155 1756
rect 8155 1722 8189 1756
rect 8189 1722 8190 1756
rect 8010 1682 8190 1722
rect 8010 1648 8011 1682
rect 8011 1648 8045 1682
rect 8045 1648 8083 1682
rect 8083 1648 8117 1682
rect 8117 1648 8155 1682
rect 8155 1648 8189 1682
rect 8189 1648 8190 1682
rect 8010 1608 8190 1648
rect 8010 1574 8011 1608
rect 8011 1574 8045 1608
rect 8045 1574 8083 1608
rect 8083 1574 8117 1608
rect 8117 1574 8155 1608
rect 8155 1574 8189 1608
rect 8189 1574 8190 1608
rect 8010 1568 8190 1574
rect 8506 4092 8558 4124
rect 8570 4118 8622 4124
rect 8570 4092 8579 4118
rect 8579 4092 8613 4118
rect 8613 4092 8622 4118
rect 8634 4092 8686 4124
rect 8506 4072 8507 4092
rect 8507 4072 8558 4092
rect 8570 4072 8622 4092
rect 8634 4072 8685 4092
rect 8685 4072 8686 4092
rect 8506 4007 8507 4059
rect 8507 4007 8558 4059
rect 8570 4007 8622 4059
rect 8634 4007 8685 4059
rect 8685 4007 8686 4059
rect 8506 3942 8507 3994
rect 8507 3942 8558 3994
rect 8570 3942 8622 3994
rect 8634 3942 8685 3994
rect 8685 3942 8686 3994
rect 8506 3877 8507 3929
rect 8507 3877 8558 3929
rect 8570 3877 8622 3929
rect 8634 3877 8685 3929
rect 8685 3877 8686 3929
rect 8506 3812 8507 3864
rect 8507 3812 8558 3864
rect 8570 3812 8622 3864
rect 8634 3812 8685 3864
rect 8685 3812 8686 3864
rect 8506 3747 8507 3799
rect 8507 3747 8558 3799
rect 8570 3747 8622 3799
rect 8634 3747 8685 3799
rect 8685 3747 8686 3799
rect 8506 3682 8507 3734
rect 8507 3682 8558 3734
rect 8570 3682 8622 3734
rect 8634 3682 8685 3734
rect 8685 3682 8686 3734
rect 8506 3617 8507 3669
rect 8507 3617 8558 3669
rect 8570 3617 8622 3669
rect 8634 3617 8685 3669
rect 8685 3617 8686 3669
rect 8506 3194 8507 3604
rect 8507 3194 8685 3604
rect 8685 3194 8686 3604
rect 8506 3182 8686 3194
rect 8506 3148 8579 3182
rect 8579 3148 8613 3182
rect 8613 3148 8686 3182
rect 8506 3108 8686 3148
rect 8506 3074 8507 3108
rect 8507 3074 8541 3108
rect 8541 3074 8579 3108
rect 8579 3074 8613 3108
rect 8613 3074 8651 3108
rect 8651 3074 8685 3108
rect 8685 3074 8686 3108
rect 8506 3028 8686 3074
rect 8506 2994 8507 3028
rect 8507 2994 8541 3028
rect 8541 2994 8579 3028
rect 8579 2994 8613 3028
rect 8613 2994 8651 3028
rect 8651 2994 8685 3028
rect 8685 2994 8686 3028
rect 8506 2948 8686 2994
rect 8506 2914 8507 2948
rect 8507 2914 8541 2948
rect 8541 2914 8579 2948
rect 8579 2914 8613 2948
rect 8613 2914 8651 2948
rect 8651 2914 8685 2948
rect 8685 2914 8686 2948
rect 8506 2868 8686 2914
rect 8506 2834 8507 2868
rect 8507 2834 8541 2868
rect 8541 2834 8579 2868
rect 8579 2834 8613 2868
rect 8613 2834 8651 2868
rect 8651 2834 8685 2868
rect 8685 2834 8686 2868
rect 8506 2788 8686 2834
rect 8506 2754 8507 2788
rect 8507 2754 8541 2788
rect 8541 2754 8579 2788
rect 8579 2754 8613 2788
rect 8613 2754 8651 2788
rect 8651 2754 8685 2788
rect 8685 2754 8686 2788
rect 8506 2708 8686 2754
rect 8506 2674 8507 2708
rect 8507 2674 8541 2708
rect 8541 2674 8579 2708
rect 8579 2674 8613 2708
rect 8613 2674 8651 2708
rect 8651 2674 8685 2708
rect 8685 2674 8686 2708
rect 8506 2628 8686 2674
rect 8506 2594 8507 2628
rect 8507 2594 8541 2628
rect 8541 2594 8579 2628
rect 8579 2594 8613 2628
rect 8613 2594 8651 2628
rect 8651 2594 8685 2628
rect 8685 2594 8686 2628
rect 8506 2556 8686 2594
rect 8506 2522 8579 2556
rect 8579 2522 8613 2556
rect 8613 2522 8686 2556
rect 8506 2518 8686 2522
rect 8506 1620 8507 2518
rect 8507 1620 8685 2518
rect 8685 1620 8686 2518
rect 8506 1586 8579 1620
rect 8579 1586 8613 1620
rect 8613 1586 8686 1620
rect 8506 1568 8686 1586
rect 9002 4098 9054 4119
rect 9002 4067 9003 4098
rect 9003 4067 9037 4098
rect 9037 4067 9054 4098
rect 9066 4098 9118 4119
rect 9066 4067 9075 4098
rect 9075 4067 9109 4098
rect 9109 4067 9118 4098
rect 9130 4098 9182 4119
rect 9130 4067 9147 4098
rect 9147 4067 9181 4098
rect 9181 4067 9182 4098
rect 9002 4025 9054 4054
rect 9002 4002 9003 4025
rect 9003 4002 9037 4025
rect 9037 4002 9054 4025
rect 9066 4025 9118 4054
rect 9066 4002 9075 4025
rect 9075 4002 9109 4025
rect 9109 4002 9118 4025
rect 9130 4025 9182 4054
rect 9130 4002 9147 4025
rect 9147 4002 9181 4025
rect 9181 4002 9182 4025
rect 9002 3952 9054 3989
rect 9002 3937 9003 3952
rect 9003 3937 9037 3952
rect 9037 3937 9054 3952
rect 9066 3952 9118 3989
rect 9066 3937 9075 3952
rect 9075 3937 9109 3952
rect 9109 3937 9118 3952
rect 9130 3952 9182 3989
rect 9130 3937 9147 3952
rect 9147 3937 9181 3952
rect 9181 3937 9182 3952
rect 9002 3918 9003 3924
rect 9003 3918 9037 3924
rect 9037 3918 9075 3924
rect 9075 3918 9109 3924
rect 9109 3918 9147 3924
rect 9147 3918 9181 3924
rect 9181 3918 9182 3924
rect 9002 3879 9182 3918
rect 9002 3845 9003 3879
rect 9003 3845 9037 3879
rect 9037 3845 9075 3879
rect 9075 3845 9109 3879
rect 9109 3845 9147 3879
rect 9147 3845 9181 3879
rect 9181 3845 9182 3879
rect 9002 3806 9182 3845
rect 9002 3772 9003 3806
rect 9003 3772 9037 3806
rect 9037 3772 9075 3806
rect 9075 3772 9109 3806
rect 9109 3772 9147 3806
rect 9147 3772 9181 3806
rect 9181 3772 9182 3806
rect 9002 3733 9182 3772
rect 9002 3699 9003 3733
rect 9003 3699 9037 3733
rect 9037 3699 9075 3733
rect 9075 3699 9109 3733
rect 9109 3699 9147 3733
rect 9147 3699 9181 3733
rect 9181 3699 9182 3733
rect 9002 3660 9182 3699
rect 9002 3626 9003 3660
rect 9003 3626 9037 3660
rect 9037 3626 9075 3660
rect 9075 3626 9109 3660
rect 9109 3626 9147 3660
rect 9147 3626 9181 3660
rect 9181 3626 9182 3660
rect 9002 3587 9182 3626
rect 9002 3553 9003 3587
rect 9003 3553 9037 3587
rect 9037 3553 9075 3587
rect 9075 3553 9109 3587
rect 9109 3553 9147 3587
rect 9147 3553 9181 3587
rect 9181 3553 9182 3587
rect 9002 3514 9182 3553
rect 9002 3480 9003 3514
rect 9003 3480 9037 3514
rect 9037 3480 9075 3514
rect 9075 3480 9109 3514
rect 9109 3480 9147 3514
rect 9147 3480 9181 3514
rect 9181 3480 9182 3514
rect 9002 3441 9182 3480
rect 9002 3407 9003 3441
rect 9003 3407 9037 3441
rect 9037 3407 9075 3441
rect 9075 3407 9109 3441
rect 9109 3407 9147 3441
rect 9147 3407 9181 3441
rect 9181 3407 9182 3441
rect 9002 3368 9182 3407
rect 9002 3334 9003 3368
rect 9003 3334 9037 3368
rect 9037 3334 9075 3368
rect 9075 3334 9109 3368
rect 9109 3334 9147 3368
rect 9147 3334 9181 3368
rect 9181 3334 9182 3368
rect 9002 3295 9182 3334
rect 9002 3261 9003 3295
rect 9003 3261 9037 3295
rect 9037 3261 9075 3295
rect 9075 3261 9109 3295
rect 9109 3261 9147 3295
rect 9147 3261 9181 3295
rect 9181 3261 9182 3295
rect 9002 3222 9182 3261
rect 9002 3188 9003 3222
rect 9003 3188 9037 3222
rect 9037 3188 9075 3222
rect 9075 3188 9109 3222
rect 9109 3188 9147 3222
rect 9147 3188 9181 3222
rect 9181 3188 9182 3222
rect 9002 3149 9182 3188
rect 9002 3115 9003 3149
rect 9003 3115 9037 3149
rect 9037 3115 9075 3149
rect 9075 3115 9109 3149
rect 9109 3115 9147 3149
rect 9147 3115 9181 3149
rect 9181 3115 9182 3149
rect 9002 3076 9182 3115
rect 9002 3042 9003 3076
rect 9003 3042 9037 3076
rect 9037 3042 9075 3076
rect 9075 3042 9109 3076
rect 9109 3042 9147 3076
rect 9147 3042 9181 3076
rect 9181 3042 9182 3076
rect 9002 3003 9182 3042
rect 9002 2969 9003 3003
rect 9003 2969 9037 3003
rect 9037 2969 9075 3003
rect 9075 2969 9109 3003
rect 9109 2969 9147 3003
rect 9147 2969 9181 3003
rect 9181 2969 9182 3003
rect 9002 2930 9182 2969
rect 9002 2896 9003 2930
rect 9003 2896 9037 2930
rect 9037 2896 9075 2930
rect 9075 2896 9109 2930
rect 9109 2896 9147 2930
rect 9147 2896 9181 2930
rect 9181 2896 9182 2930
rect 9002 2857 9182 2896
rect 9002 2823 9003 2857
rect 9003 2823 9037 2857
rect 9037 2823 9075 2857
rect 9075 2823 9109 2857
rect 9109 2823 9147 2857
rect 9147 2823 9181 2857
rect 9181 2823 9182 2857
rect 9002 2784 9182 2823
rect 9002 2750 9003 2784
rect 9003 2750 9037 2784
rect 9037 2750 9075 2784
rect 9075 2750 9109 2784
rect 9109 2750 9147 2784
rect 9147 2750 9181 2784
rect 9181 2750 9182 2784
rect 9002 2711 9182 2750
rect 9002 2677 9003 2711
rect 9003 2677 9037 2711
rect 9037 2677 9075 2711
rect 9075 2677 9109 2711
rect 9109 2677 9147 2711
rect 9147 2677 9181 2711
rect 9181 2677 9182 2711
rect 9002 2638 9182 2677
rect 9002 2604 9003 2638
rect 9003 2604 9037 2638
rect 9037 2604 9075 2638
rect 9075 2604 9109 2638
rect 9109 2604 9147 2638
rect 9147 2604 9181 2638
rect 9181 2604 9182 2638
rect 9002 2565 9182 2604
rect 9002 2531 9003 2565
rect 9003 2531 9037 2565
rect 9037 2531 9075 2565
rect 9075 2531 9109 2565
rect 9109 2531 9147 2565
rect 9147 2531 9181 2565
rect 9181 2531 9182 2565
rect 9002 2492 9182 2531
rect 9002 2458 9003 2492
rect 9003 2458 9037 2492
rect 9037 2458 9075 2492
rect 9075 2458 9109 2492
rect 9109 2458 9147 2492
rect 9147 2458 9181 2492
rect 9181 2458 9182 2492
rect 9002 2419 9182 2458
rect 9002 2385 9003 2419
rect 9003 2385 9037 2419
rect 9037 2385 9075 2419
rect 9075 2385 9109 2419
rect 9109 2385 9147 2419
rect 9147 2385 9181 2419
rect 9181 2385 9182 2419
rect 9002 2346 9182 2385
rect 9002 2312 9003 2346
rect 9003 2312 9037 2346
rect 9037 2312 9075 2346
rect 9075 2312 9109 2346
rect 9109 2312 9147 2346
rect 9147 2312 9181 2346
rect 9181 2312 9182 2346
rect 9002 2273 9182 2312
rect 9002 2239 9003 2273
rect 9003 2239 9037 2273
rect 9037 2239 9075 2273
rect 9075 2239 9109 2273
rect 9109 2239 9147 2273
rect 9147 2239 9181 2273
rect 9181 2239 9182 2273
rect 9002 2200 9182 2239
rect 9002 2166 9003 2200
rect 9003 2166 9037 2200
rect 9037 2166 9075 2200
rect 9075 2166 9109 2200
rect 9109 2166 9147 2200
rect 9147 2166 9181 2200
rect 9181 2166 9182 2200
rect 9002 2126 9182 2166
rect 9002 2092 9003 2126
rect 9003 2092 9037 2126
rect 9037 2092 9075 2126
rect 9075 2092 9109 2126
rect 9109 2092 9147 2126
rect 9147 2092 9181 2126
rect 9181 2092 9182 2126
rect 9002 2052 9182 2092
rect 9002 2018 9003 2052
rect 9003 2018 9037 2052
rect 9037 2018 9075 2052
rect 9075 2018 9109 2052
rect 9109 2018 9147 2052
rect 9147 2018 9181 2052
rect 9181 2018 9182 2052
rect 9002 1978 9182 2018
rect 9002 1944 9003 1978
rect 9003 1944 9037 1978
rect 9037 1944 9075 1978
rect 9075 1944 9109 1978
rect 9109 1944 9147 1978
rect 9147 1944 9181 1978
rect 9181 1944 9182 1978
rect 9002 1904 9182 1944
rect 9002 1870 9003 1904
rect 9003 1870 9037 1904
rect 9037 1870 9075 1904
rect 9075 1870 9109 1904
rect 9109 1870 9147 1904
rect 9147 1870 9181 1904
rect 9181 1870 9182 1904
rect 9002 1830 9182 1870
rect 9002 1796 9003 1830
rect 9003 1796 9037 1830
rect 9037 1796 9075 1830
rect 9075 1796 9109 1830
rect 9109 1796 9147 1830
rect 9147 1796 9181 1830
rect 9181 1796 9182 1830
rect 9002 1756 9182 1796
rect 9002 1722 9003 1756
rect 9003 1722 9037 1756
rect 9037 1722 9075 1756
rect 9075 1722 9109 1756
rect 9109 1722 9147 1756
rect 9147 1722 9181 1756
rect 9181 1722 9182 1756
rect 9002 1682 9182 1722
rect 9002 1648 9003 1682
rect 9003 1648 9037 1682
rect 9037 1648 9075 1682
rect 9075 1648 9109 1682
rect 9109 1648 9147 1682
rect 9147 1648 9181 1682
rect 9181 1648 9182 1682
rect 9002 1608 9182 1648
rect 9002 1574 9003 1608
rect 9003 1574 9037 1608
rect 9037 1574 9075 1608
rect 9075 1574 9109 1608
rect 9109 1574 9147 1608
rect 9147 1574 9181 1608
rect 9181 1574 9182 1608
rect 9002 1568 9182 1574
rect 9498 4092 9550 4124
rect 9562 4118 9614 4124
rect 9562 4092 9571 4118
rect 9571 4092 9605 4118
rect 9605 4092 9614 4118
rect 9626 4092 9678 4124
rect 9498 4072 9499 4092
rect 9499 4072 9550 4092
rect 9562 4072 9614 4092
rect 9626 4072 9677 4092
rect 9677 4072 9678 4092
rect 9498 4007 9499 4059
rect 9499 4007 9550 4059
rect 9562 4007 9614 4059
rect 9626 4007 9677 4059
rect 9677 4007 9678 4059
rect 9498 3942 9499 3994
rect 9499 3942 9550 3994
rect 9562 3942 9614 3994
rect 9626 3942 9677 3994
rect 9677 3942 9678 3994
rect 9498 3877 9499 3929
rect 9499 3877 9550 3929
rect 9562 3877 9614 3929
rect 9626 3877 9677 3929
rect 9677 3877 9678 3929
rect 9498 3812 9499 3864
rect 9499 3812 9550 3864
rect 9562 3812 9614 3864
rect 9626 3812 9677 3864
rect 9677 3812 9678 3864
rect 9498 3747 9499 3799
rect 9499 3747 9550 3799
rect 9562 3747 9614 3799
rect 9626 3747 9677 3799
rect 9677 3747 9678 3799
rect 9498 3682 9499 3734
rect 9499 3682 9550 3734
rect 9562 3682 9614 3734
rect 9626 3682 9677 3734
rect 9677 3682 9678 3734
rect 9498 3617 9499 3669
rect 9499 3617 9550 3669
rect 9562 3617 9614 3669
rect 9626 3617 9677 3669
rect 9677 3617 9678 3669
rect 9498 3194 9499 3604
rect 9499 3194 9677 3604
rect 9677 3194 9678 3604
rect 9498 3182 9678 3194
rect 9498 3148 9571 3182
rect 9571 3148 9605 3182
rect 9605 3148 9678 3182
rect 9498 3108 9678 3148
rect 9498 3074 9499 3108
rect 9499 3074 9533 3108
rect 9533 3074 9571 3108
rect 9571 3074 9605 3108
rect 9605 3074 9643 3108
rect 9643 3074 9677 3108
rect 9677 3074 9678 3108
rect 9498 3028 9678 3074
rect 9498 2994 9499 3028
rect 9499 2994 9533 3028
rect 9533 2994 9571 3028
rect 9571 2994 9605 3028
rect 9605 2994 9643 3028
rect 9643 2994 9677 3028
rect 9677 2994 9678 3028
rect 9498 2948 9678 2994
rect 9498 2914 9499 2948
rect 9499 2914 9533 2948
rect 9533 2914 9571 2948
rect 9571 2914 9605 2948
rect 9605 2914 9643 2948
rect 9643 2914 9677 2948
rect 9677 2914 9678 2948
rect 9498 2868 9678 2914
rect 9498 2834 9499 2868
rect 9499 2834 9533 2868
rect 9533 2834 9571 2868
rect 9571 2834 9605 2868
rect 9605 2834 9643 2868
rect 9643 2834 9677 2868
rect 9677 2834 9678 2868
rect 9498 2788 9678 2834
rect 9498 2754 9499 2788
rect 9499 2754 9533 2788
rect 9533 2754 9571 2788
rect 9571 2754 9605 2788
rect 9605 2754 9643 2788
rect 9643 2754 9677 2788
rect 9677 2754 9678 2788
rect 9498 2708 9678 2754
rect 9498 2674 9499 2708
rect 9499 2674 9533 2708
rect 9533 2674 9571 2708
rect 9571 2674 9605 2708
rect 9605 2674 9643 2708
rect 9643 2674 9677 2708
rect 9677 2674 9678 2708
rect 9498 2628 9678 2674
rect 9498 2594 9499 2628
rect 9499 2594 9533 2628
rect 9533 2594 9571 2628
rect 9571 2594 9605 2628
rect 9605 2594 9643 2628
rect 9643 2594 9677 2628
rect 9677 2594 9678 2628
rect 9498 2556 9678 2594
rect 9498 2522 9571 2556
rect 9571 2522 9605 2556
rect 9605 2522 9678 2556
rect 9498 2518 9678 2522
rect 9498 1620 9499 2518
rect 9499 1620 9677 2518
rect 9677 1620 9678 2518
rect 9498 1586 9571 1620
rect 9571 1586 9605 1620
rect 9605 1586 9678 1620
rect 9498 1568 9678 1586
rect 9994 4098 10046 4119
rect 9994 4067 9995 4098
rect 9995 4067 10029 4098
rect 10029 4067 10046 4098
rect 10058 4098 10110 4119
rect 10058 4067 10067 4098
rect 10067 4067 10101 4098
rect 10101 4067 10110 4098
rect 10122 4098 10174 4119
rect 10122 4067 10139 4098
rect 10139 4067 10173 4098
rect 10173 4067 10174 4098
rect 9994 4025 10046 4054
rect 9994 4002 9995 4025
rect 9995 4002 10029 4025
rect 10029 4002 10046 4025
rect 10058 4025 10110 4054
rect 10058 4002 10067 4025
rect 10067 4002 10101 4025
rect 10101 4002 10110 4025
rect 10122 4025 10174 4054
rect 10122 4002 10139 4025
rect 10139 4002 10173 4025
rect 10173 4002 10174 4025
rect 9994 3952 10046 3989
rect 9994 3937 9995 3952
rect 9995 3937 10029 3952
rect 10029 3937 10046 3952
rect 10058 3952 10110 3989
rect 10058 3937 10067 3952
rect 10067 3937 10101 3952
rect 10101 3937 10110 3952
rect 10122 3952 10174 3989
rect 10122 3937 10139 3952
rect 10139 3937 10173 3952
rect 10173 3937 10174 3952
rect 9994 3918 9995 3924
rect 9995 3918 10029 3924
rect 10029 3918 10067 3924
rect 10067 3918 10101 3924
rect 10101 3918 10139 3924
rect 10139 3918 10173 3924
rect 10173 3918 10174 3924
rect 9994 3879 10174 3918
rect 9994 3845 9995 3879
rect 9995 3845 10029 3879
rect 10029 3845 10067 3879
rect 10067 3845 10101 3879
rect 10101 3845 10139 3879
rect 10139 3845 10173 3879
rect 10173 3845 10174 3879
rect 9994 3806 10174 3845
rect 9994 3772 9995 3806
rect 9995 3772 10029 3806
rect 10029 3772 10067 3806
rect 10067 3772 10101 3806
rect 10101 3772 10139 3806
rect 10139 3772 10173 3806
rect 10173 3772 10174 3806
rect 9994 3733 10174 3772
rect 9994 3699 9995 3733
rect 9995 3699 10029 3733
rect 10029 3699 10067 3733
rect 10067 3699 10101 3733
rect 10101 3699 10139 3733
rect 10139 3699 10173 3733
rect 10173 3699 10174 3733
rect 9994 3660 10174 3699
rect 9994 3626 9995 3660
rect 9995 3626 10029 3660
rect 10029 3626 10067 3660
rect 10067 3626 10101 3660
rect 10101 3626 10139 3660
rect 10139 3626 10173 3660
rect 10173 3626 10174 3660
rect 9994 3587 10174 3626
rect 9994 3553 9995 3587
rect 9995 3553 10029 3587
rect 10029 3553 10067 3587
rect 10067 3553 10101 3587
rect 10101 3553 10139 3587
rect 10139 3553 10173 3587
rect 10173 3553 10174 3587
rect 9994 3514 10174 3553
rect 9994 3480 9995 3514
rect 9995 3480 10029 3514
rect 10029 3480 10067 3514
rect 10067 3480 10101 3514
rect 10101 3480 10139 3514
rect 10139 3480 10173 3514
rect 10173 3480 10174 3514
rect 9994 3441 10174 3480
rect 9994 3407 9995 3441
rect 9995 3407 10029 3441
rect 10029 3407 10067 3441
rect 10067 3407 10101 3441
rect 10101 3407 10139 3441
rect 10139 3407 10173 3441
rect 10173 3407 10174 3441
rect 9994 3368 10174 3407
rect 9994 3334 9995 3368
rect 9995 3334 10029 3368
rect 10029 3334 10067 3368
rect 10067 3334 10101 3368
rect 10101 3334 10139 3368
rect 10139 3334 10173 3368
rect 10173 3334 10174 3368
rect 9994 3295 10174 3334
rect 9994 3261 9995 3295
rect 9995 3261 10029 3295
rect 10029 3261 10067 3295
rect 10067 3261 10101 3295
rect 10101 3261 10139 3295
rect 10139 3261 10173 3295
rect 10173 3261 10174 3295
rect 9994 3222 10174 3261
rect 9994 3188 9995 3222
rect 9995 3188 10029 3222
rect 10029 3188 10067 3222
rect 10067 3188 10101 3222
rect 10101 3188 10139 3222
rect 10139 3188 10173 3222
rect 10173 3188 10174 3222
rect 9994 3149 10174 3188
rect 9994 3115 9995 3149
rect 9995 3115 10029 3149
rect 10029 3115 10067 3149
rect 10067 3115 10101 3149
rect 10101 3115 10139 3149
rect 10139 3115 10173 3149
rect 10173 3115 10174 3149
rect 9994 3076 10174 3115
rect 9994 3042 9995 3076
rect 9995 3042 10029 3076
rect 10029 3042 10067 3076
rect 10067 3042 10101 3076
rect 10101 3042 10139 3076
rect 10139 3042 10173 3076
rect 10173 3042 10174 3076
rect 9994 3003 10174 3042
rect 9994 2969 9995 3003
rect 9995 2969 10029 3003
rect 10029 2969 10067 3003
rect 10067 2969 10101 3003
rect 10101 2969 10139 3003
rect 10139 2969 10173 3003
rect 10173 2969 10174 3003
rect 9994 2930 10174 2969
rect 9994 2896 9995 2930
rect 9995 2896 10029 2930
rect 10029 2896 10067 2930
rect 10067 2896 10101 2930
rect 10101 2896 10139 2930
rect 10139 2896 10173 2930
rect 10173 2896 10174 2930
rect 9994 2857 10174 2896
rect 9994 2823 9995 2857
rect 9995 2823 10029 2857
rect 10029 2823 10067 2857
rect 10067 2823 10101 2857
rect 10101 2823 10139 2857
rect 10139 2823 10173 2857
rect 10173 2823 10174 2857
rect 9994 2784 10174 2823
rect 9994 2750 9995 2784
rect 9995 2750 10029 2784
rect 10029 2750 10067 2784
rect 10067 2750 10101 2784
rect 10101 2750 10139 2784
rect 10139 2750 10173 2784
rect 10173 2750 10174 2784
rect 9994 2711 10174 2750
rect 9994 2677 9995 2711
rect 9995 2677 10029 2711
rect 10029 2677 10067 2711
rect 10067 2677 10101 2711
rect 10101 2677 10139 2711
rect 10139 2677 10173 2711
rect 10173 2677 10174 2711
rect 9994 2638 10174 2677
rect 9994 2604 9995 2638
rect 9995 2604 10029 2638
rect 10029 2604 10067 2638
rect 10067 2604 10101 2638
rect 10101 2604 10139 2638
rect 10139 2604 10173 2638
rect 10173 2604 10174 2638
rect 9994 2565 10174 2604
rect 9994 2531 9995 2565
rect 9995 2531 10029 2565
rect 10029 2531 10067 2565
rect 10067 2531 10101 2565
rect 10101 2531 10139 2565
rect 10139 2531 10173 2565
rect 10173 2531 10174 2565
rect 9994 2492 10174 2531
rect 9994 2458 9995 2492
rect 9995 2458 10029 2492
rect 10029 2458 10067 2492
rect 10067 2458 10101 2492
rect 10101 2458 10139 2492
rect 10139 2458 10173 2492
rect 10173 2458 10174 2492
rect 9994 2419 10174 2458
rect 9994 2385 9995 2419
rect 9995 2385 10029 2419
rect 10029 2385 10067 2419
rect 10067 2385 10101 2419
rect 10101 2385 10139 2419
rect 10139 2385 10173 2419
rect 10173 2385 10174 2419
rect 9994 2346 10174 2385
rect 9994 2312 9995 2346
rect 9995 2312 10029 2346
rect 10029 2312 10067 2346
rect 10067 2312 10101 2346
rect 10101 2312 10139 2346
rect 10139 2312 10173 2346
rect 10173 2312 10174 2346
rect 9994 2273 10174 2312
rect 9994 2239 9995 2273
rect 9995 2239 10029 2273
rect 10029 2239 10067 2273
rect 10067 2239 10101 2273
rect 10101 2239 10139 2273
rect 10139 2239 10173 2273
rect 10173 2239 10174 2273
rect 9994 2200 10174 2239
rect 9994 2166 9995 2200
rect 9995 2166 10029 2200
rect 10029 2166 10067 2200
rect 10067 2166 10101 2200
rect 10101 2166 10139 2200
rect 10139 2166 10173 2200
rect 10173 2166 10174 2200
rect 9994 2126 10174 2166
rect 9994 2092 9995 2126
rect 9995 2092 10029 2126
rect 10029 2092 10067 2126
rect 10067 2092 10101 2126
rect 10101 2092 10139 2126
rect 10139 2092 10173 2126
rect 10173 2092 10174 2126
rect 9994 2052 10174 2092
rect 9994 2018 9995 2052
rect 9995 2018 10029 2052
rect 10029 2018 10067 2052
rect 10067 2018 10101 2052
rect 10101 2018 10139 2052
rect 10139 2018 10173 2052
rect 10173 2018 10174 2052
rect 9994 1978 10174 2018
rect 9994 1944 9995 1978
rect 9995 1944 10029 1978
rect 10029 1944 10067 1978
rect 10067 1944 10101 1978
rect 10101 1944 10139 1978
rect 10139 1944 10173 1978
rect 10173 1944 10174 1978
rect 9994 1904 10174 1944
rect 9994 1870 9995 1904
rect 9995 1870 10029 1904
rect 10029 1870 10067 1904
rect 10067 1870 10101 1904
rect 10101 1870 10139 1904
rect 10139 1870 10173 1904
rect 10173 1870 10174 1904
rect 9994 1830 10174 1870
rect 9994 1796 9995 1830
rect 9995 1796 10029 1830
rect 10029 1796 10067 1830
rect 10067 1796 10101 1830
rect 10101 1796 10139 1830
rect 10139 1796 10173 1830
rect 10173 1796 10174 1830
rect 9994 1756 10174 1796
rect 9994 1722 9995 1756
rect 9995 1722 10029 1756
rect 10029 1722 10067 1756
rect 10067 1722 10101 1756
rect 10101 1722 10139 1756
rect 10139 1722 10173 1756
rect 10173 1722 10174 1756
rect 9994 1682 10174 1722
rect 9994 1648 9995 1682
rect 9995 1648 10029 1682
rect 10029 1648 10067 1682
rect 10067 1648 10101 1682
rect 10101 1648 10139 1682
rect 10139 1648 10173 1682
rect 10173 1648 10174 1682
rect 9994 1608 10174 1648
rect 9994 1574 9995 1608
rect 9995 1574 10029 1608
rect 10029 1574 10067 1608
rect 10067 1574 10101 1608
rect 10101 1574 10139 1608
rect 10139 1574 10173 1608
rect 10173 1574 10174 1608
rect 9994 1568 10174 1574
rect 10490 4092 10542 4124
rect 10554 4118 10606 4124
rect 10554 4092 10563 4118
rect 10563 4092 10597 4118
rect 10597 4092 10606 4118
rect 10618 4092 10670 4124
rect 10490 4072 10491 4092
rect 10491 4072 10542 4092
rect 10554 4072 10606 4092
rect 10618 4072 10669 4092
rect 10669 4072 10670 4092
rect 10490 4007 10491 4059
rect 10491 4007 10542 4059
rect 10554 4007 10606 4059
rect 10618 4007 10669 4059
rect 10669 4007 10670 4059
rect 10490 3942 10491 3994
rect 10491 3942 10542 3994
rect 10554 3942 10606 3994
rect 10618 3942 10669 3994
rect 10669 3942 10670 3994
rect 10490 3877 10491 3929
rect 10491 3877 10542 3929
rect 10554 3877 10606 3929
rect 10618 3877 10669 3929
rect 10669 3877 10670 3929
rect 10490 3812 10491 3864
rect 10491 3812 10542 3864
rect 10554 3812 10606 3864
rect 10618 3812 10669 3864
rect 10669 3812 10670 3864
rect 10490 3747 10491 3799
rect 10491 3747 10542 3799
rect 10554 3747 10606 3799
rect 10618 3747 10669 3799
rect 10669 3747 10670 3799
rect 10490 3682 10491 3734
rect 10491 3682 10542 3734
rect 10554 3682 10606 3734
rect 10618 3682 10669 3734
rect 10669 3682 10670 3734
rect 10490 3617 10491 3669
rect 10491 3617 10542 3669
rect 10554 3617 10606 3669
rect 10618 3617 10669 3669
rect 10669 3617 10670 3669
rect 10490 3194 10491 3604
rect 10491 3194 10669 3604
rect 10669 3194 10670 3604
rect 10490 3182 10670 3194
rect 10490 3148 10563 3182
rect 10563 3148 10597 3182
rect 10597 3148 10670 3182
rect 10490 3108 10670 3148
rect 10490 3074 10491 3108
rect 10491 3074 10525 3108
rect 10525 3074 10563 3108
rect 10563 3074 10597 3108
rect 10597 3074 10635 3108
rect 10635 3074 10669 3108
rect 10669 3074 10670 3108
rect 10490 3028 10670 3074
rect 10490 2994 10491 3028
rect 10491 2994 10525 3028
rect 10525 2994 10563 3028
rect 10563 2994 10597 3028
rect 10597 2994 10635 3028
rect 10635 2994 10669 3028
rect 10669 2994 10670 3028
rect 10490 2948 10670 2994
rect 10490 2914 10491 2948
rect 10491 2914 10525 2948
rect 10525 2914 10563 2948
rect 10563 2914 10597 2948
rect 10597 2914 10635 2948
rect 10635 2914 10669 2948
rect 10669 2914 10670 2948
rect 10490 2868 10670 2914
rect 10490 2834 10491 2868
rect 10491 2834 10525 2868
rect 10525 2834 10563 2868
rect 10563 2834 10597 2868
rect 10597 2834 10635 2868
rect 10635 2834 10669 2868
rect 10669 2834 10670 2868
rect 10490 2788 10670 2834
rect 10490 2754 10491 2788
rect 10491 2754 10525 2788
rect 10525 2754 10563 2788
rect 10563 2754 10597 2788
rect 10597 2754 10635 2788
rect 10635 2754 10669 2788
rect 10669 2754 10670 2788
rect 10490 2708 10670 2754
rect 10490 2674 10491 2708
rect 10491 2674 10525 2708
rect 10525 2674 10563 2708
rect 10563 2674 10597 2708
rect 10597 2674 10635 2708
rect 10635 2674 10669 2708
rect 10669 2674 10670 2708
rect 10490 2628 10670 2674
rect 10490 2594 10491 2628
rect 10491 2594 10525 2628
rect 10525 2594 10563 2628
rect 10563 2594 10597 2628
rect 10597 2594 10635 2628
rect 10635 2594 10669 2628
rect 10669 2594 10670 2628
rect 10490 2556 10670 2594
rect 10490 2522 10563 2556
rect 10563 2522 10597 2556
rect 10597 2522 10670 2556
rect 10490 2518 10670 2522
rect 10490 1620 10491 2518
rect 10491 1620 10669 2518
rect 10669 1620 10670 2518
rect 10490 1586 10563 1620
rect 10563 1586 10597 1620
rect 10597 1586 10670 1620
rect 10490 1568 10670 1586
rect 10986 4098 11038 4119
rect 10986 4067 10987 4098
rect 10987 4067 11021 4098
rect 11021 4067 11038 4098
rect 11050 4098 11102 4119
rect 11050 4067 11059 4098
rect 11059 4067 11093 4098
rect 11093 4067 11102 4098
rect 11114 4098 11166 4119
rect 11114 4067 11131 4098
rect 11131 4067 11165 4098
rect 11165 4067 11166 4098
rect 10986 4025 11038 4054
rect 10986 4002 10987 4025
rect 10987 4002 11021 4025
rect 11021 4002 11038 4025
rect 11050 4025 11102 4054
rect 11050 4002 11059 4025
rect 11059 4002 11093 4025
rect 11093 4002 11102 4025
rect 11114 4025 11166 4054
rect 11114 4002 11131 4025
rect 11131 4002 11165 4025
rect 11165 4002 11166 4025
rect 10986 3952 11038 3989
rect 10986 3937 10987 3952
rect 10987 3937 11021 3952
rect 11021 3937 11038 3952
rect 11050 3952 11102 3989
rect 11050 3937 11059 3952
rect 11059 3937 11093 3952
rect 11093 3937 11102 3952
rect 11114 3952 11166 3989
rect 11114 3937 11131 3952
rect 11131 3937 11165 3952
rect 11165 3937 11166 3952
rect 10986 3918 10987 3924
rect 10987 3918 11021 3924
rect 11021 3918 11059 3924
rect 11059 3918 11093 3924
rect 11093 3918 11131 3924
rect 11131 3918 11165 3924
rect 11165 3918 11166 3924
rect 10986 3879 11166 3918
rect 10986 3845 10987 3879
rect 10987 3845 11021 3879
rect 11021 3845 11059 3879
rect 11059 3845 11093 3879
rect 11093 3845 11131 3879
rect 11131 3845 11165 3879
rect 11165 3845 11166 3879
rect 10986 3806 11166 3845
rect 10986 3772 10987 3806
rect 10987 3772 11021 3806
rect 11021 3772 11059 3806
rect 11059 3772 11093 3806
rect 11093 3772 11131 3806
rect 11131 3772 11165 3806
rect 11165 3772 11166 3806
rect 10986 3733 11166 3772
rect 10986 3699 10987 3733
rect 10987 3699 11021 3733
rect 11021 3699 11059 3733
rect 11059 3699 11093 3733
rect 11093 3699 11131 3733
rect 11131 3699 11165 3733
rect 11165 3699 11166 3733
rect 10986 3660 11166 3699
rect 10986 3626 10987 3660
rect 10987 3626 11021 3660
rect 11021 3626 11059 3660
rect 11059 3626 11093 3660
rect 11093 3626 11131 3660
rect 11131 3626 11165 3660
rect 11165 3626 11166 3660
rect 10986 3587 11166 3626
rect 10986 3553 10987 3587
rect 10987 3553 11021 3587
rect 11021 3553 11059 3587
rect 11059 3553 11093 3587
rect 11093 3553 11131 3587
rect 11131 3553 11165 3587
rect 11165 3553 11166 3587
rect 10986 3514 11166 3553
rect 10986 3480 10987 3514
rect 10987 3480 11021 3514
rect 11021 3480 11059 3514
rect 11059 3480 11093 3514
rect 11093 3480 11131 3514
rect 11131 3480 11165 3514
rect 11165 3480 11166 3514
rect 10986 3441 11166 3480
rect 10986 3407 10987 3441
rect 10987 3407 11021 3441
rect 11021 3407 11059 3441
rect 11059 3407 11093 3441
rect 11093 3407 11131 3441
rect 11131 3407 11165 3441
rect 11165 3407 11166 3441
rect 10986 3368 11166 3407
rect 10986 3334 10987 3368
rect 10987 3334 11021 3368
rect 11021 3334 11059 3368
rect 11059 3334 11093 3368
rect 11093 3334 11131 3368
rect 11131 3334 11165 3368
rect 11165 3334 11166 3368
rect 10986 3295 11166 3334
rect 10986 3261 10987 3295
rect 10987 3261 11021 3295
rect 11021 3261 11059 3295
rect 11059 3261 11093 3295
rect 11093 3261 11131 3295
rect 11131 3261 11165 3295
rect 11165 3261 11166 3295
rect 10986 3222 11166 3261
rect 10986 3188 10987 3222
rect 10987 3188 11021 3222
rect 11021 3188 11059 3222
rect 11059 3188 11093 3222
rect 11093 3188 11131 3222
rect 11131 3188 11165 3222
rect 11165 3188 11166 3222
rect 10986 3149 11166 3188
rect 10986 3115 10987 3149
rect 10987 3115 11021 3149
rect 11021 3115 11059 3149
rect 11059 3115 11093 3149
rect 11093 3115 11131 3149
rect 11131 3115 11165 3149
rect 11165 3115 11166 3149
rect 10986 3076 11166 3115
rect 10986 3042 10987 3076
rect 10987 3042 11021 3076
rect 11021 3042 11059 3076
rect 11059 3042 11093 3076
rect 11093 3042 11131 3076
rect 11131 3042 11165 3076
rect 11165 3042 11166 3076
rect 10986 3003 11166 3042
rect 10986 2969 10987 3003
rect 10987 2969 11021 3003
rect 11021 2969 11059 3003
rect 11059 2969 11093 3003
rect 11093 2969 11131 3003
rect 11131 2969 11165 3003
rect 11165 2969 11166 3003
rect 10986 2930 11166 2969
rect 10986 2896 10987 2930
rect 10987 2896 11021 2930
rect 11021 2896 11059 2930
rect 11059 2896 11093 2930
rect 11093 2896 11131 2930
rect 11131 2896 11165 2930
rect 11165 2896 11166 2930
rect 10986 2857 11166 2896
rect 10986 2823 10987 2857
rect 10987 2823 11021 2857
rect 11021 2823 11059 2857
rect 11059 2823 11093 2857
rect 11093 2823 11131 2857
rect 11131 2823 11165 2857
rect 11165 2823 11166 2857
rect 10986 2784 11166 2823
rect 10986 2750 10987 2784
rect 10987 2750 11021 2784
rect 11021 2750 11059 2784
rect 11059 2750 11093 2784
rect 11093 2750 11131 2784
rect 11131 2750 11165 2784
rect 11165 2750 11166 2784
rect 10986 2711 11166 2750
rect 10986 2677 10987 2711
rect 10987 2677 11021 2711
rect 11021 2677 11059 2711
rect 11059 2677 11093 2711
rect 11093 2677 11131 2711
rect 11131 2677 11165 2711
rect 11165 2677 11166 2711
rect 10986 2638 11166 2677
rect 10986 2604 10987 2638
rect 10987 2604 11021 2638
rect 11021 2604 11059 2638
rect 11059 2604 11093 2638
rect 11093 2604 11131 2638
rect 11131 2604 11165 2638
rect 11165 2604 11166 2638
rect 10986 2565 11166 2604
rect 10986 2531 10987 2565
rect 10987 2531 11021 2565
rect 11021 2531 11059 2565
rect 11059 2531 11093 2565
rect 11093 2531 11131 2565
rect 11131 2531 11165 2565
rect 11165 2531 11166 2565
rect 10986 2492 11166 2531
rect 10986 2458 10987 2492
rect 10987 2458 11021 2492
rect 11021 2458 11059 2492
rect 11059 2458 11093 2492
rect 11093 2458 11131 2492
rect 11131 2458 11165 2492
rect 11165 2458 11166 2492
rect 10986 2419 11166 2458
rect 10986 2385 10987 2419
rect 10987 2385 11021 2419
rect 11021 2385 11059 2419
rect 11059 2385 11093 2419
rect 11093 2385 11131 2419
rect 11131 2385 11165 2419
rect 11165 2385 11166 2419
rect 10986 2346 11166 2385
rect 10986 2312 10987 2346
rect 10987 2312 11021 2346
rect 11021 2312 11059 2346
rect 11059 2312 11093 2346
rect 11093 2312 11131 2346
rect 11131 2312 11165 2346
rect 11165 2312 11166 2346
rect 10986 2273 11166 2312
rect 10986 2239 10987 2273
rect 10987 2239 11021 2273
rect 11021 2239 11059 2273
rect 11059 2239 11093 2273
rect 11093 2239 11131 2273
rect 11131 2239 11165 2273
rect 11165 2239 11166 2273
rect 10986 2200 11166 2239
rect 10986 2166 10987 2200
rect 10987 2166 11021 2200
rect 11021 2166 11059 2200
rect 11059 2166 11093 2200
rect 11093 2166 11131 2200
rect 11131 2166 11165 2200
rect 11165 2166 11166 2200
rect 10986 2126 11166 2166
rect 10986 2092 10987 2126
rect 10987 2092 11021 2126
rect 11021 2092 11059 2126
rect 11059 2092 11093 2126
rect 11093 2092 11131 2126
rect 11131 2092 11165 2126
rect 11165 2092 11166 2126
rect 10986 2052 11166 2092
rect 10986 2018 10987 2052
rect 10987 2018 11021 2052
rect 11021 2018 11059 2052
rect 11059 2018 11093 2052
rect 11093 2018 11131 2052
rect 11131 2018 11165 2052
rect 11165 2018 11166 2052
rect 10986 1978 11166 2018
rect 10986 1944 10987 1978
rect 10987 1944 11021 1978
rect 11021 1944 11059 1978
rect 11059 1944 11093 1978
rect 11093 1944 11131 1978
rect 11131 1944 11165 1978
rect 11165 1944 11166 1978
rect 10986 1904 11166 1944
rect 10986 1870 10987 1904
rect 10987 1870 11021 1904
rect 11021 1870 11059 1904
rect 11059 1870 11093 1904
rect 11093 1870 11131 1904
rect 11131 1870 11165 1904
rect 11165 1870 11166 1904
rect 10986 1830 11166 1870
rect 10986 1796 10987 1830
rect 10987 1796 11021 1830
rect 11021 1796 11059 1830
rect 11059 1796 11093 1830
rect 11093 1796 11131 1830
rect 11131 1796 11165 1830
rect 11165 1796 11166 1830
rect 10986 1756 11166 1796
rect 10986 1722 10987 1756
rect 10987 1722 11021 1756
rect 11021 1722 11059 1756
rect 11059 1722 11093 1756
rect 11093 1722 11131 1756
rect 11131 1722 11165 1756
rect 11165 1722 11166 1756
rect 10986 1682 11166 1722
rect 10986 1648 10987 1682
rect 10987 1648 11021 1682
rect 11021 1648 11059 1682
rect 11059 1648 11093 1682
rect 11093 1648 11131 1682
rect 11131 1648 11165 1682
rect 11165 1648 11166 1682
rect 10986 1608 11166 1648
rect 10986 1574 10987 1608
rect 10987 1574 11021 1608
rect 11021 1574 11059 1608
rect 11059 1574 11093 1608
rect 11093 1574 11131 1608
rect 11131 1574 11165 1608
rect 11165 1574 11166 1608
rect 10986 1568 11166 1574
rect 11482 4092 11534 4124
rect 11546 4118 11598 4124
rect 11546 4092 11555 4118
rect 11555 4092 11589 4118
rect 11589 4092 11598 4118
rect 11610 4092 11662 4124
rect 11482 4072 11483 4092
rect 11483 4072 11534 4092
rect 11546 4072 11598 4092
rect 11610 4072 11661 4092
rect 11661 4072 11662 4092
rect 11482 4007 11483 4059
rect 11483 4007 11534 4059
rect 11546 4007 11598 4059
rect 11610 4007 11661 4059
rect 11661 4007 11662 4059
rect 11482 3942 11483 3994
rect 11483 3942 11534 3994
rect 11546 3942 11598 3994
rect 11610 3942 11661 3994
rect 11661 3942 11662 3994
rect 11482 3877 11483 3929
rect 11483 3877 11534 3929
rect 11546 3877 11598 3929
rect 11610 3877 11661 3929
rect 11661 3877 11662 3929
rect 11482 3812 11483 3864
rect 11483 3812 11534 3864
rect 11546 3812 11598 3864
rect 11610 3812 11661 3864
rect 11661 3812 11662 3864
rect 11482 3747 11483 3799
rect 11483 3747 11534 3799
rect 11546 3747 11598 3799
rect 11610 3747 11661 3799
rect 11661 3747 11662 3799
rect 11482 3682 11483 3734
rect 11483 3682 11534 3734
rect 11546 3682 11598 3734
rect 11610 3682 11661 3734
rect 11661 3682 11662 3734
rect 11482 3617 11483 3669
rect 11483 3617 11534 3669
rect 11546 3617 11598 3669
rect 11610 3617 11661 3669
rect 11661 3617 11662 3669
rect 11482 3194 11483 3604
rect 11483 3194 11661 3604
rect 11661 3194 11662 3604
rect 11482 3182 11662 3194
rect 11482 3148 11555 3182
rect 11555 3148 11589 3182
rect 11589 3148 11662 3182
rect 11482 3108 11662 3148
rect 11482 3074 11483 3108
rect 11483 3074 11517 3108
rect 11517 3074 11555 3108
rect 11555 3074 11589 3108
rect 11589 3074 11627 3108
rect 11627 3074 11661 3108
rect 11661 3074 11662 3108
rect 11482 3028 11662 3074
rect 11482 2994 11483 3028
rect 11483 2994 11517 3028
rect 11517 2994 11555 3028
rect 11555 2994 11589 3028
rect 11589 2994 11627 3028
rect 11627 2994 11661 3028
rect 11661 2994 11662 3028
rect 11482 2948 11662 2994
rect 11482 2914 11483 2948
rect 11483 2914 11517 2948
rect 11517 2914 11555 2948
rect 11555 2914 11589 2948
rect 11589 2914 11627 2948
rect 11627 2914 11661 2948
rect 11661 2914 11662 2948
rect 11482 2868 11662 2914
rect 11482 2834 11483 2868
rect 11483 2834 11517 2868
rect 11517 2834 11555 2868
rect 11555 2834 11589 2868
rect 11589 2834 11627 2868
rect 11627 2834 11661 2868
rect 11661 2834 11662 2868
rect 11482 2788 11662 2834
rect 11482 2754 11483 2788
rect 11483 2754 11517 2788
rect 11517 2754 11555 2788
rect 11555 2754 11589 2788
rect 11589 2754 11627 2788
rect 11627 2754 11661 2788
rect 11661 2754 11662 2788
rect 11482 2708 11662 2754
rect 11482 2674 11483 2708
rect 11483 2674 11517 2708
rect 11517 2674 11555 2708
rect 11555 2674 11589 2708
rect 11589 2674 11627 2708
rect 11627 2674 11661 2708
rect 11661 2674 11662 2708
rect 11482 2628 11662 2674
rect 11482 2594 11483 2628
rect 11483 2594 11517 2628
rect 11517 2594 11555 2628
rect 11555 2594 11589 2628
rect 11589 2594 11627 2628
rect 11627 2594 11661 2628
rect 11661 2594 11662 2628
rect 11482 2556 11662 2594
rect 11482 2522 11555 2556
rect 11555 2522 11589 2556
rect 11589 2522 11662 2556
rect 11482 2518 11662 2522
rect 11482 1620 11483 2518
rect 11483 1620 11661 2518
rect 11661 1620 11662 2518
rect 11482 1586 11555 1620
rect 11555 1586 11589 1620
rect 11589 1586 11662 1620
rect 11482 1568 11662 1586
rect 11978 4098 12030 4119
rect 11978 4067 11979 4098
rect 11979 4067 12013 4098
rect 12013 4067 12030 4098
rect 12042 4098 12094 4119
rect 12042 4067 12051 4098
rect 12051 4067 12085 4098
rect 12085 4067 12094 4098
rect 12106 4098 12158 4119
rect 12106 4067 12123 4098
rect 12123 4067 12157 4098
rect 12157 4067 12158 4098
rect 11978 4025 12030 4054
rect 11978 4002 11979 4025
rect 11979 4002 12013 4025
rect 12013 4002 12030 4025
rect 12042 4025 12094 4054
rect 12042 4002 12051 4025
rect 12051 4002 12085 4025
rect 12085 4002 12094 4025
rect 12106 4025 12158 4054
rect 12106 4002 12123 4025
rect 12123 4002 12157 4025
rect 12157 4002 12158 4025
rect 11978 3952 12030 3989
rect 11978 3937 11979 3952
rect 11979 3937 12013 3952
rect 12013 3937 12030 3952
rect 12042 3952 12094 3989
rect 12042 3937 12051 3952
rect 12051 3937 12085 3952
rect 12085 3937 12094 3952
rect 12106 3952 12158 3989
rect 12106 3937 12123 3952
rect 12123 3937 12157 3952
rect 12157 3937 12158 3952
rect 11978 3918 11979 3924
rect 11979 3918 12013 3924
rect 12013 3918 12051 3924
rect 12051 3918 12085 3924
rect 12085 3918 12123 3924
rect 12123 3918 12157 3924
rect 12157 3918 12158 3924
rect 11978 3879 12158 3918
rect 11978 3845 11979 3879
rect 11979 3845 12013 3879
rect 12013 3845 12051 3879
rect 12051 3845 12085 3879
rect 12085 3845 12123 3879
rect 12123 3845 12157 3879
rect 12157 3845 12158 3879
rect 11978 3806 12158 3845
rect 11978 3772 11979 3806
rect 11979 3772 12013 3806
rect 12013 3772 12051 3806
rect 12051 3772 12085 3806
rect 12085 3772 12123 3806
rect 12123 3772 12157 3806
rect 12157 3772 12158 3806
rect 11978 3733 12158 3772
rect 11978 3699 11979 3733
rect 11979 3699 12013 3733
rect 12013 3699 12051 3733
rect 12051 3699 12085 3733
rect 12085 3699 12123 3733
rect 12123 3699 12157 3733
rect 12157 3699 12158 3733
rect 11978 3660 12158 3699
rect 11978 3626 11979 3660
rect 11979 3626 12013 3660
rect 12013 3626 12051 3660
rect 12051 3626 12085 3660
rect 12085 3626 12123 3660
rect 12123 3626 12157 3660
rect 12157 3626 12158 3660
rect 11978 3587 12158 3626
rect 11978 3553 11979 3587
rect 11979 3553 12013 3587
rect 12013 3553 12051 3587
rect 12051 3553 12085 3587
rect 12085 3553 12123 3587
rect 12123 3553 12157 3587
rect 12157 3553 12158 3587
rect 11978 3514 12158 3553
rect 11978 3480 11979 3514
rect 11979 3480 12013 3514
rect 12013 3480 12051 3514
rect 12051 3480 12085 3514
rect 12085 3480 12123 3514
rect 12123 3480 12157 3514
rect 12157 3480 12158 3514
rect 11978 3441 12158 3480
rect 11978 3407 11979 3441
rect 11979 3407 12013 3441
rect 12013 3407 12051 3441
rect 12051 3407 12085 3441
rect 12085 3407 12123 3441
rect 12123 3407 12157 3441
rect 12157 3407 12158 3441
rect 11978 3368 12158 3407
rect 11978 3334 11979 3368
rect 11979 3334 12013 3368
rect 12013 3334 12051 3368
rect 12051 3334 12085 3368
rect 12085 3334 12123 3368
rect 12123 3334 12157 3368
rect 12157 3334 12158 3368
rect 11978 3295 12158 3334
rect 11978 3261 11979 3295
rect 11979 3261 12013 3295
rect 12013 3261 12051 3295
rect 12051 3261 12085 3295
rect 12085 3261 12123 3295
rect 12123 3261 12157 3295
rect 12157 3261 12158 3295
rect 11978 3222 12158 3261
rect 11978 3188 11979 3222
rect 11979 3188 12013 3222
rect 12013 3188 12051 3222
rect 12051 3188 12085 3222
rect 12085 3188 12123 3222
rect 12123 3188 12157 3222
rect 12157 3188 12158 3222
rect 11978 3149 12158 3188
rect 11978 3115 11979 3149
rect 11979 3115 12013 3149
rect 12013 3115 12051 3149
rect 12051 3115 12085 3149
rect 12085 3115 12123 3149
rect 12123 3115 12157 3149
rect 12157 3115 12158 3149
rect 11978 3076 12158 3115
rect 11978 3042 11979 3076
rect 11979 3042 12013 3076
rect 12013 3042 12051 3076
rect 12051 3042 12085 3076
rect 12085 3042 12123 3076
rect 12123 3042 12157 3076
rect 12157 3042 12158 3076
rect 11978 3003 12158 3042
rect 11978 2969 11979 3003
rect 11979 2969 12013 3003
rect 12013 2969 12051 3003
rect 12051 2969 12085 3003
rect 12085 2969 12123 3003
rect 12123 2969 12157 3003
rect 12157 2969 12158 3003
rect 11978 2930 12158 2969
rect 11978 2896 11979 2930
rect 11979 2896 12013 2930
rect 12013 2896 12051 2930
rect 12051 2896 12085 2930
rect 12085 2896 12123 2930
rect 12123 2896 12157 2930
rect 12157 2896 12158 2930
rect 11978 2857 12158 2896
rect 11978 2823 11979 2857
rect 11979 2823 12013 2857
rect 12013 2823 12051 2857
rect 12051 2823 12085 2857
rect 12085 2823 12123 2857
rect 12123 2823 12157 2857
rect 12157 2823 12158 2857
rect 11978 2784 12158 2823
rect 11978 2750 11979 2784
rect 11979 2750 12013 2784
rect 12013 2750 12051 2784
rect 12051 2750 12085 2784
rect 12085 2750 12123 2784
rect 12123 2750 12157 2784
rect 12157 2750 12158 2784
rect 11978 2711 12158 2750
rect 11978 2677 11979 2711
rect 11979 2677 12013 2711
rect 12013 2677 12051 2711
rect 12051 2677 12085 2711
rect 12085 2677 12123 2711
rect 12123 2677 12157 2711
rect 12157 2677 12158 2711
rect 11978 2638 12158 2677
rect 11978 2604 11979 2638
rect 11979 2604 12013 2638
rect 12013 2604 12051 2638
rect 12051 2604 12085 2638
rect 12085 2604 12123 2638
rect 12123 2604 12157 2638
rect 12157 2604 12158 2638
rect 11978 2565 12158 2604
rect 11978 2531 11979 2565
rect 11979 2531 12013 2565
rect 12013 2531 12051 2565
rect 12051 2531 12085 2565
rect 12085 2531 12123 2565
rect 12123 2531 12157 2565
rect 12157 2531 12158 2565
rect 11978 2492 12158 2531
rect 11978 2458 11979 2492
rect 11979 2458 12013 2492
rect 12013 2458 12051 2492
rect 12051 2458 12085 2492
rect 12085 2458 12123 2492
rect 12123 2458 12157 2492
rect 12157 2458 12158 2492
rect 11978 2419 12158 2458
rect 11978 2385 11979 2419
rect 11979 2385 12013 2419
rect 12013 2385 12051 2419
rect 12051 2385 12085 2419
rect 12085 2385 12123 2419
rect 12123 2385 12157 2419
rect 12157 2385 12158 2419
rect 11978 2346 12158 2385
rect 11978 2312 11979 2346
rect 11979 2312 12013 2346
rect 12013 2312 12051 2346
rect 12051 2312 12085 2346
rect 12085 2312 12123 2346
rect 12123 2312 12157 2346
rect 12157 2312 12158 2346
rect 11978 2273 12158 2312
rect 11978 2239 11979 2273
rect 11979 2239 12013 2273
rect 12013 2239 12051 2273
rect 12051 2239 12085 2273
rect 12085 2239 12123 2273
rect 12123 2239 12157 2273
rect 12157 2239 12158 2273
rect 11978 2200 12158 2239
rect 11978 2166 11979 2200
rect 11979 2166 12013 2200
rect 12013 2166 12051 2200
rect 12051 2166 12085 2200
rect 12085 2166 12123 2200
rect 12123 2166 12157 2200
rect 12157 2166 12158 2200
rect 11978 2126 12158 2166
rect 11978 2092 11979 2126
rect 11979 2092 12013 2126
rect 12013 2092 12051 2126
rect 12051 2092 12085 2126
rect 12085 2092 12123 2126
rect 12123 2092 12157 2126
rect 12157 2092 12158 2126
rect 11978 2052 12158 2092
rect 11978 2018 11979 2052
rect 11979 2018 12013 2052
rect 12013 2018 12051 2052
rect 12051 2018 12085 2052
rect 12085 2018 12123 2052
rect 12123 2018 12157 2052
rect 12157 2018 12158 2052
rect 11978 1978 12158 2018
rect 11978 1944 11979 1978
rect 11979 1944 12013 1978
rect 12013 1944 12051 1978
rect 12051 1944 12085 1978
rect 12085 1944 12123 1978
rect 12123 1944 12157 1978
rect 12157 1944 12158 1978
rect 11978 1904 12158 1944
rect 11978 1870 11979 1904
rect 11979 1870 12013 1904
rect 12013 1870 12051 1904
rect 12051 1870 12085 1904
rect 12085 1870 12123 1904
rect 12123 1870 12157 1904
rect 12157 1870 12158 1904
rect 11978 1830 12158 1870
rect 11978 1796 11979 1830
rect 11979 1796 12013 1830
rect 12013 1796 12051 1830
rect 12051 1796 12085 1830
rect 12085 1796 12123 1830
rect 12123 1796 12157 1830
rect 12157 1796 12158 1830
rect 11978 1756 12158 1796
rect 11978 1722 11979 1756
rect 11979 1722 12013 1756
rect 12013 1722 12051 1756
rect 12051 1722 12085 1756
rect 12085 1722 12123 1756
rect 12123 1722 12157 1756
rect 12157 1722 12158 1756
rect 11978 1682 12158 1722
rect 11978 1648 11979 1682
rect 11979 1648 12013 1682
rect 12013 1648 12051 1682
rect 12051 1648 12085 1682
rect 12085 1648 12123 1682
rect 12123 1648 12157 1682
rect 12157 1648 12158 1682
rect 11978 1608 12158 1648
rect 11978 1574 11979 1608
rect 11979 1574 12013 1608
rect 12013 1574 12051 1608
rect 12051 1574 12085 1608
rect 12085 1574 12123 1608
rect 12123 1574 12157 1608
rect 12157 1574 12158 1608
rect 11978 1568 12158 1574
rect 12474 4092 12526 4124
rect 12538 4118 12590 4124
rect 12538 4092 12547 4118
rect 12547 4092 12581 4118
rect 12581 4092 12590 4118
rect 12602 4092 12654 4124
rect 12474 4072 12475 4092
rect 12475 4072 12526 4092
rect 12538 4072 12590 4092
rect 12602 4072 12653 4092
rect 12653 4072 12654 4092
rect 12474 4007 12475 4059
rect 12475 4007 12526 4059
rect 12538 4007 12590 4059
rect 12602 4007 12653 4059
rect 12653 4007 12654 4059
rect 12474 3942 12475 3994
rect 12475 3942 12526 3994
rect 12538 3942 12590 3994
rect 12602 3942 12653 3994
rect 12653 3942 12654 3994
rect 12474 3877 12475 3929
rect 12475 3877 12526 3929
rect 12538 3877 12590 3929
rect 12602 3877 12653 3929
rect 12653 3877 12654 3929
rect 12474 3812 12475 3864
rect 12475 3812 12526 3864
rect 12538 3812 12590 3864
rect 12602 3812 12653 3864
rect 12653 3812 12654 3864
rect 12474 3747 12475 3799
rect 12475 3747 12526 3799
rect 12538 3747 12590 3799
rect 12602 3747 12653 3799
rect 12653 3747 12654 3799
rect 12474 3682 12475 3734
rect 12475 3682 12526 3734
rect 12538 3682 12590 3734
rect 12602 3682 12653 3734
rect 12653 3682 12654 3734
rect 12474 3617 12475 3669
rect 12475 3617 12526 3669
rect 12538 3617 12590 3669
rect 12602 3617 12653 3669
rect 12653 3617 12654 3669
rect 12474 3194 12475 3604
rect 12475 3194 12653 3604
rect 12653 3194 12654 3604
rect 12474 3182 12654 3194
rect 12474 3148 12547 3182
rect 12547 3148 12581 3182
rect 12581 3148 12654 3182
rect 12474 3108 12654 3148
rect 12474 3074 12475 3108
rect 12475 3074 12509 3108
rect 12509 3074 12547 3108
rect 12547 3074 12581 3108
rect 12581 3074 12619 3108
rect 12619 3074 12653 3108
rect 12653 3074 12654 3108
rect 12474 3028 12654 3074
rect 12474 2994 12475 3028
rect 12475 2994 12509 3028
rect 12509 2994 12547 3028
rect 12547 2994 12581 3028
rect 12581 2994 12619 3028
rect 12619 2994 12653 3028
rect 12653 2994 12654 3028
rect 12474 2948 12654 2994
rect 12474 2914 12475 2948
rect 12475 2914 12509 2948
rect 12509 2914 12547 2948
rect 12547 2914 12581 2948
rect 12581 2914 12619 2948
rect 12619 2914 12653 2948
rect 12653 2914 12654 2948
rect 12474 2868 12654 2914
rect 12474 2834 12475 2868
rect 12475 2834 12509 2868
rect 12509 2834 12547 2868
rect 12547 2834 12581 2868
rect 12581 2834 12619 2868
rect 12619 2834 12653 2868
rect 12653 2834 12654 2868
rect 12474 2788 12654 2834
rect 12474 2754 12475 2788
rect 12475 2754 12509 2788
rect 12509 2754 12547 2788
rect 12547 2754 12581 2788
rect 12581 2754 12619 2788
rect 12619 2754 12653 2788
rect 12653 2754 12654 2788
rect 12474 2708 12654 2754
rect 12474 2674 12475 2708
rect 12475 2674 12509 2708
rect 12509 2674 12547 2708
rect 12547 2674 12581 2708
rect 12581 2674 12619 2708
rect 12619 2674 12653 2708
rect 12653 2674 12654 2708
rect 12474 2628 12654 2674
rect 12474 2594 12475 2628
rect 12475 2594 12509 2628
rect 12509 2594 12547 2628
rect 12547 2594 12581 2628
rect 12581 2594 12619 2628
rect 12619 2594 12653 2628
rect 12653 2594 12654 2628
rect 12474 2556 12654 2594
rect 12474 2522 12547 2556
rect 12547 2522 12581 2556
rect 12581 2522 12654 2556
rect 12474 2518 12654 2522
rect 12474 1620 12475 2518
rect 12475 1620 12653 2518
rect 12653 1620 12654 2518
rect 12474 1586 12547 1620
rect 12547 1586 12581 1620
rect 12581 1586 12654 1620
rect 12474 1568 12654 1586
rect 12970 4098 13022 4119
rect 12970 4067 12971 4098
rect 12971 4067 13005 4098
rect 13005 4067 13022 4098
rect 13034 4098 13086 4119
rect 13034 4067 13043 4098
rect 13043 4067 13077 4098
rect 13077 4067 13086 4098
rect 13098 4098 13150 4119
rect 13098 4067 13115 4098
rect 13115 4067 13149 4098
rect 13149 4067 13150 4098
rect 12970 4025 13022 4054
rect 12970 4002 12971 4025
rect 12971 4002 13005 4025
rect 13005 4002 13022 4025
rect 13034 4025 13086 4054
rect 13034 4002 13043 4025
rect 13043 4002 13077 4025
rect 13077 4002 13086 4025
rect 13098 4025 13150 4054
rect 13098 4002 13115 4025
rect 13115 4002 13149 4025
rect 13149 4002 13150 4025
rect 12970 3952 13022 3989
rect 12970 3937 12971 3952
rect 12971 3937 13005 3952
rect 13005 3937 13022 3952
rect 13034 3952 13086 3989
rect 13034 3937 13043 3952
rect 13043 3937 13077 3952
rect 13077 3937 13086 3952
rect 13098 3952 13150 3989
rect 13098 3937 13115 3952
rect 13115 3937 13149 3952
rect 13149 3937 13150 3952
rect 12970 3918 12971 3924
rect 12971 3918 13005 3924
rect 13005 3918 13043 3924
rect 13043 3918 13077 3924
rect 13077 3918 13115 3924
rect 13115 3918 13149 3924
rect 13149 3918 13150 3924
rect 12970 3879 13150 3918
rect 12970 3845 12971 3879
rect 12971 3845 13005 3879
rect 13005 3845 13043 3879
rect 13043 3845 13077 3879
rect 13077 3845 13115 3879
rect 13115 3845 13149 3879
rect 13149 3845 13150 3879
rect 12970 3806 13150 3845
rect 12970 3772 12971 3806
rect 12971 3772 13005 3806
rect 13005 3772 13043 3806
rect 13043 3772 13077 3806
rect 13077 3772 13115 3806
rect 13115 3772 13149 3806
rect 13149 3772 13150 3806
rect 12970 3733 13150 3772
rect 12970 3699 12971 3733
rect 12971 3699 13005 3733
rect 13005 3699 13043 3733
rect 13043 3699 13077 3733
rect 13077 3699 13115 3733
rect 13115 3699 13149 3733
rect 13149 3699 13150 3733
rect 12970 3660 13150 3699
rect 12970 3626 12971 3660
rect 12971 3626 13005 3660
rect 13005 3626 13043 3660
rect 13043 3626 13077 3660
rect 13077 3626 13115 3660
rect 13115 3626 13149 3660
rect 13149 3626 13150 3660
rect 12970 3587 13150 3626
rect 12970 3553 12971 3587
rect 12971 3553 13005 3587
rect 13005 3553 13043 3587
rect 13043 3553 13077 3587
rect 13077 3553 13115 3587
rect 13115 3553 13149 3587
rect 13149 3553 13150 3587
rect 12970 3514 13150 3553
rect 12970 3480 12971 3514
rect 12971 3480 13005 3514
rect 13005 3480 13043 3514
rect 13043 3480 13077 3514
rect 13077 3480 13115 3514
rect 13115 3480 13149 3514
rect 13149 3480 13150 3514
rect 12970 3441 13150 3480
rect 12970 3407 12971 3441
rect 12971 3407 13005 3441
rect 13005 3407 13043 3441
rect 13043 3407 13077 3441
rect 13077 3407 13115 3441
rect 13115 3407 13149 3441
rect 13149 3407 13150 3441
rect 12970 3368 13150 3407
rect 12970 3334 12971 3368
rect 12971 3334 13005 3368
rect 13005 3334 13043 3368
rect 13043 3334 13077 3368
rect 13077 3334 13115 3368
rect 13115 3334 13149 3368
rect 13149 3334 13150 3368
rect 12970 3295 13150 3334
rect 12970 3261 12971 3295
rect 12971 3261 13005 3295
rect 13005 3261 13043 3295
rect 13043 3261 13077 3295
rect 13077 3261 13115 3295
rect 13115 3261 13149 3295
rect 13149 3261 13150 3295
rect 12970 3222 13150 3261
rect 12970 3188 12971 3222
rect 12971 3188 13005 3222
rect 13005 3188 13043 3222
rect 13043 3188 13077 3222
rect 13077 3188 13115 3222
rect 13115 3188 13149 3222
rect 13149 3188 13150 3222
rect 12970 3149 13150 3188
rect 12970 3115 12971 3149
rect 12971 3115 13005 3149
rect 13005 3115 13043 3149
rect 13043 3115 13077 3149
rect 13077 3115 13115 3149
rect 13115 3115 13149 3149
rect 13149 3115 13150 3149
rect 12970 3076 13150 3115
rect 12970 3042 12971 3076
rect 12971 3042 13005 3076
rect 13005 3042 13043 3076
rect 13043 3042 13077 3076
rect 13077 3042 13115 3076
rect 13115 3042 13149 3076
rect 13149 3042 13150 3076
rect 12970 3003 13150 3042
rect 12970 2969 12971 3003
rect 12971 2969 13005 3003
rect 13005 2969 13043 3003
rect 13043 2969 13077 3003
rect 13077 2969 13115 3003
rect 13115 2969 13149 3003
rect 13149 2969 13150 3003
rect 12970 2930 13150 2969
rect 12970 2896 12971 2930
rect 12971 2896 13005 2930
rect 13005 2896 13043 2930
rect 13043 2896 13077 2930
rect 13077 2896 13115 2930
rect 13115 2896 13149 2930
rect 13149 2896 13150 2930
rect 12970 2857 13150 2896
rect 12970 2823 12971 2857
rect 12971 2823 13005 2857
rect 13005 2823 13043 2857
rect 13043 2823 13077 2857
rect 13077 2823 13115 2857
rect 13115 2823 13149 2857
rect 13149 2823 13150 2857
rect 12970 2784 13150 2823
rect 12970 2750 12971 2784
rect 12971 2750 13005 2784
rect 13005 2750 13043 2784
rect 13043 2750 13077 2784
rect 13077 2750 13115 2784
rect 13115 2750 13149 2784
rect 13149 2750 13150 2784
rect 12970 2711 13150 2750
rect 12970 2677 12971 2711
rect 12971 2677 13005 2711
rect 13005 2677 13043 2711
rect 13043 2677 13077 2711
rect 13077 2677 13115 2711
rect 13115 2677 13149 2711
rect 13149 2677 13150 2711
rect 12970 2638 13150 2677
rect 12970 2604 12971 2638
rect 12971 2604 13005 2638
rect 13005 2604 13043 2638
rect 13043 2604 13077 2638
rect 13077 2604 13115 2638
rect 13115 2604 13149 2638
rect 13149 2604 13150 2638
rect 12970 2565 13150 2604
rect 12970 2531 12971 2565
rect 12971 2531 13005 2565
rect 13005 2531 13043 2565
rect 13043 2531 13077 2565
rect 13077 2531 13115 2565
rect 13115 2531 13149 2565
rect 13149 2531 13150 2565
rect 12970 2492 13150 2531
rect 12970 2458 12971 2492
rect 12971 2458 13005 2492
rect 13005 2458 13043 2492
rect 13043 2458 13077 2492
rect 13077 2458 13115 2492
rect 13115 2458 13149 2492
rect 13149 2458 13150 2492
rect 12970 2419 13150 2458
rect 12970 2385 12971 2419
rect 12971 2385 13005 2419
rect 13005 2385 13043 2419
rect 13043 2385 13077 2419
rect 13077 2385 13115 2419
rect 13115 2385 13149 2419
rect 13149 2385 13150 2419
rect 12970 2346 13150 2385
rect 12970 2312 12971 2346
rect 12971 2312 13005 2346
rect 13005 2312 13043 2346
rect 13043 2312 13077 2346
rect 13077 2312 13115 2346
rect 13115 2312 13149 2346
rect 13149 2312 13150 2346
rect 12970 2273 13150 2312
rect 12970 2239 12971 2273
rect 12971 2239 13005 2273
rect 13005 2239 13043 2273
rect 13043 2239 13077 2273
rect 13077 2239 13115 2273
rect 13115 2239 13149 2273
rect 13149 2239 13150 2273
rect 12970 2200 13150 2239
rect 12970 2166 12971 2200
rect 12971 2166 13005 2200
rect 13005 2166 13043 2200
rect 13043 2166 13077 2200
rect 13077 2166 13115 2200
rect 13115 2166 13149 2200
rect 13149 2166 13150 2200
rect 12970 2126 13150 2166
rect 12970 2092 12971 2126
rect 12971 2092 13005 2126
rect 13005 2092 13043 2126
rect 13043 2092 13077 2126
rect 13077 2092 13115 2126
rect 13115 2092 13149 2126
rect 13149 2092 13150 2126
rect 12970 2052 13150 2092
rect 12970 2018 12971 2052
rect 12971 2018 13005 2052
rect 13005 2018 13043 2052
rect 13043 2018 13077 2052
rect 13077 2018 13115 2052
rect 13115 2018 13149 2052
rect 13149 2018 13150 2052
rect 12970 1978 13150 2018
rect 12970 1944 12971 1978
rect 12971 1944 13005 1978
rect 13005 1944 13043 1978
rect 13043 1944 13077 1978
rect 13077 1944 13115 1978
rect 13115 1944 13149 1978
rect 13149 1944 13150 1978
rect 12970 1904 13150 1944
rect 12970 1870 12971 1904
rect 12971 1870 13005 1904
rect 13005 1870 13043 1904
rect 13043 1870 13077 1904
rect 13077 1870 13115 1904
rect 13115 1870 13149 1904
rect 13149 1870 13150 1904
rect 12970 1830 13150 1870
rect 12970 1796 12971 1830
rect 12971 1796 13005 1830
rect 13005 1796 13043 1830
rect 13043 1796 13077 1830
rect 13077 1796 13115 1830
rect 13115 1796 13149 1830
rect 13149 1796 13150 1830
rect 12970 1756 13150 1796
rect 12970 1722 12971 1756
rect 12971 1722 13005 1756
rect 13005 1722 13043 1756
rect 13043 1722 13077 1756
rect 13077 1722 13115 1756
rect 13115 1722 13149 1756
rect 13149 1722 13150 1756
rect 12970 1682 13150 1722
rect 12970 1648 12971 1682
rect 12971 1648 13005 1682
rect 13005 1648 13043 1682
rect 13043 1648 13077 1682
rect 13077 1648 13115 1682
rect 13115 1648 13149 1682
rect 13149 1648 13150 1682
rect 12970 1608 13150 1648
rect 12970 1574 12971 1608
rect 12971 1574 13005 1608
rect 13005 1574 13043 1608
rect 13043 1574 13077 1608
rect 13077 1574 13115 1608
rect 13115 1574 13149 1608
rect 13149 1574 13150 1608
rect 12970 1568 13150 1574
rect 13466 4092 13518 4124
rect 13530 4118 13582 4124
rect 13530 4092 13539 4118
rect 13539 4092 13573 4118
rect 13573 4092 13582 4118
rect 13594 4092 13646 4124
rect 13466 4072 13467 4092
rect 13467 4072 13518 4092
rect 13530 4072 13582 4092
rect 13594 4072 13645 4092
rect 13645 4072 13646 4092
rect 13466 4007 13467 4059
rect 13467 4007 13518 4059
rect 13530 4007 13582 4059
rect 13594 4007 13645 4059
rect 13645 4007 13646 4059
rect 13466 3942 13467 3994
rect 13467 3942 13518 3994
rect 13530 3942 13582 3994
rect 13594 3942 13645 3994
rect 13645 3942 13646 3994
rect 13466 3877 13467 3929
rect 13467 3877 13518 3929
rect 13530 3877 13582 3929
rect 13594 3877 13645 3929
rect 13645 3877 13646 3929
rect 13466 3812 13467 3864
rect 13467 3812 13518 3864
rect 13530 3812 13582 3864
rect 13594 3812 13645 3864
rect 13645 3812 13646 3864
rect 13466 3747 13467 3799
rect 13467 3747 13518 3799
rect 13530 3747 13582 3799
rect 13594 3747 13645 3799
rect 13645 3747 13646 3799
rect 13466 3682 13467 3734
rect 13467 3682 13518 3734
rect 13530 3682 13582 3734
rect 13594 3682 13645 3734
rect 13645 3682 13646 3734
rect 13466 3617 13467 3669
rect 13467 3617 13518 3669
rect 13530 3617 13582 3669
rect 13594 3617 13645 3669
rect 13645 3617 13646 3669
rect 13466 3194 13467 3604
rect 13467 3194 13645 3604
rect 13645 3194 13646 3604
rect 13466 3182 13646 3194
rect 13466 3148 13539 3182
rect 13539 3148 13573 3182
rect 13573 3148 13646 3182
rect 13466 3108 13646 3148
rect 13466 3074 13467 3108
rect 13467 3074 13501 3108
rect 13501 3074 13539 3108
rect 13539 3074 13573 3108
rect 13573 3074 13611 3108
rect 13611 3074 13645 3108
rect 13645 3074 13646 3108
rect 13466 3028 13646 3074
rect 13466 2994 13467 3028
rect 13467 2994 13501 3028
rect 13501 2994 13539 3028
rect 13539 2994 13573 3028
rect 13573 2994 13611 3028
rect 13611 2994 13645 3028
rect 13645 2994 13646 3028
rect 13466 2948 13646 2994
rect 13466 2914 13467 2948
rect 13467 2914 13501 2948
rect 13501 2914 13539 2948
rect 13539 2914 13573 2948
rect 13573 2914 13611 2948
rect 13611 2914 13645 2948
rect 13645 2914 13646 2948
rect 13466 2868 13646 2914
rect 13466 2834 13467 2868
rect 13467 2834 13501 2868
rect 13501 2834 13539 2868
rect 13539 2834 13573 2868
rect 13573 2834 13611 2868
rect 13611 2834 13645 2868
rect 13645 2834 13646 2868
rect 13466 2788 13646 2834
rect 13466 2754 13467 2788
rect 13467 2754 13501 2788
rect 13501 2754 13539 2788
rect 13539 2754 13573 2788
rect 13573 2754 13611 2788
rect 13611 2754 13645 2788
rect 13645 2754 13646 2788
rect 13466 2708 13646 2754
rect 13466 2674 13467 2708
rect 13467 2674 13501 2708
rect 13501 2674 13539 2708
rect 13539 2674 13573 2708
rect 13573 2674 13611 2708
rect 13611 2674 13645 2708
rect 13645 2674 13646 2708
rect 13466 2628 13646 2674
rect 13466 2594 13467 2628
rect 13467 2594 13501 2628
rect 13501 2594 13539 2628
rect 13539 2594 13573 2628
rect 13573 2594 13611 2628
rect 13611 2594 13645 2628
rect 13645 2594 13646 2628
rect 13466 2556 13646 2594
rect 13466 2522 13539 2556
rect 13539 2522 13573 2556
rect 13573 2522 13646 2556
rect 13466 2518 13646 2522
rect 13466 1620 13467 2518
rect 13467 1620 13645 2518
rect 13645 1620 13646 2518
rect 13466 1586 13539 1620
rect 13539 1586 13573 1620
rect 13573 1586 13646 1620
rect 13466 1568 13646 1586
rect 13991 4098 14043 4124
rect 13991 4072 13997 4098
rect 13997 4072 14035 4098
rect 14035 4072 14043 4098
rect 14083 4072 14135 4124
rect 13991 4024 14043 4060
rect 13991 4008 13997 4024
rect 13997 4008 14035 4024
rect 14035 4008 14043 4024
rect 14083 4008 14135 4060
rect 13991 3990 13997 3996
rect 13997 3990 14035 3996
rect 14035 3990 14043 3996
rect 13991 3950 14043 3990
rect 13991 3944 13997 3950
rect 13997 3944 14035 3950
rect 14035 3944 14043 3950
rect 14083 3944 14135 3996
rect 13991 3916 13997 3932
rect 13997 3916 14035 3932
rect 14035 3916 14043 3932
rect 13991 3880 14043 3916
rect 14083 3880 14135 3932
rect 13991 3842 13997 3868
rect 13997 3842 14035 3868
rect 14035 3842 14043 3868
rect 13991 3816 14043 3842
rect 14083 3816 14135 3868
rect 13991 3802 14043 3804
rect 13991 3768 13997 3802
rect 13997 3768 14035 3802
rect 14035 3768 14043 3802
rect 13991 3752 14043 3768
rect 14083 3752 14135 3804
rect 13991 3728 14043 3740
rect 13991 3694 13997 3728
rect 13997 3694 14035 3728
rect 14035 3694 14043 3728
rect 13991 3688 14043 3694
rect 14083 3688 14135 3740
rect 13991 3654 14043 3676
rect 13991 3624 13997 3654
rect 13997 3624 14035 3654
rect 14035 3624 14043 3654
rect 14083 3624 14135 3676
rect 13991 3580 14043 3612
rect 13991 3560 13997 3580
rect 13997 3560 14035 3580
rect 14035 3560 14043 3580
rect 14083 3560 14135 3612
rect 13991 3546 13997 3548
rect 13997 3546 14035 3548
rect 14035 3546 14043 3548
rect 13991 3506 14043 3546
rect 13991 3496 13997 3506
rect 13997 3496 14035 3506
rect 14035 3496 14043 3506
rect 14083 3496 14135 3548
rect 13991 3472 13997 3484
rect 13997 3472 14035 3484
rect 14035 3472 14043 3484
rect 13991 3432 14043 3472
rect 14083 3432 14135 3484
rect 13991 3398 13997 3420
rect 13997 3398 14035 3420
rect 14035 3398 14043 3420
rect 13991 3368 14043 3398
rect 14083 3368 14135 3420
rect 13991 3324 13997 3356
rect 13997 3324 14035 3356
rect 14035 3324 14043 3356
rect 13991 3304 14043 3324
rect 14083 3304 14135 3356
rect 13991 3284 14043 3292
rect 13991 3250 13997 3284
rect 13997 3250 14035 3284
rect 14035 3250 14043 3284
rect 13991 3240 14043 3250
rect 14083 3240 14135 3292
rect 13991 3210 14043 3228
rect 13991 3176 13997 3210
rect 13997 3176 14035 3210
rect 14035 3176 14043 3210
rect 14083 3176 14135 3228
rect 13991 3136 14043 3164
rect 13991 3112 13997 3136
rect 13997 3112 14035 3136
rect 14035 3112 14043 3136
rect 14083 3112 14135 3164
rect 13991 3062 14043 3100
rect 13991 3048 13997 3062
rect 13997 3048 14035 3062
rect 14035 3048 14043 3062
rect 14083 3048 14135 3100
rect 13991 3028 13997 3036
rect 13997 3028 14035 3036
rect 14035 3028 14043 3036
rect 13991 2988 14043 3028
rect 13991 2984 13997 2988
rect 13997 2984 14035 2988
rect 14035 2984 14043 2988
rect 14083 2984 14135 3036
rect 13991 2954 13997 2972
rect 13997 2954 14035 2972
rect 14035 2954 14043 2972
rect 13991 2920 14043 2954
rect 14083 2920 14135 2972
rect 13991 2880 13997 2908
rect 13997 2880 14035 2908
rect 14035 2880 14043 2908
rect 13991 2856 14043 2880
rect 14083 2856 14135 2908
rect 13991 2840 14043 2844
rect 13991 2806 13997 2840
rect 13997 2806 14035 2840
rect 14035 2806 14043 2840
rect 13991 2792 14043 2806
rect 14083 2792 14135 2844
rect 13991 2766 14043 2780
rect 13991 2732 13997 2766
rect 13997 2732 14035 2766
rect 14035 2732 14043 2766
rect 13991 2728 14043 2732
rect 14083 2728 14135 2780
rect 13991 2692 14043 2716
rect 13991 2664 13997 2692
rect 13997 2664 14035 2692
rect 14035 2664 14043 2692
rect 14083 2664 14135 2716
rect 13991 2618 14043 2652
rect 13991 2600 13997 2618
rect 13997 2600 14035 2618
rect 14035 2600 14043 2618
rect 14083 2600 14135 2652
rect 13991 2584 13997 2588
rect 13997 2584 14035 2588
rect 14035 2584 14043 2588
rect 13991 2544 14043 2584
rect 13991 2536 13997 2544
rect 13997 2536 14035 2544
rect 14035 2536 14043 2544
rect 14083 2536 14135 2588
rect 13991 2510 13997 2524
rect 13997 2510 14035 2524
rect 14035 2510 14043 2524
rect 13991 2472 14043 2510
rect 14083 2472 14135 2524
rect 13991 2436 13997 2460
rect 13997 2436 14035 2460
rect 14035 2436 14043 2460
rect 13991 2408 14043 2436
rect 14083 2408 14135 2460
rect 13991 2362 13997 2396
rect 13997 2362 14035 2396
rect 14035 2362 14043 2396
rect 13991 2344 14043 2362
rect 14083 2344 14135 2396
rect 13991 2322 14043 2332
rect 13991 2288 13997 2322
rect 13997 2288 14035 2322
rect 14035 2288 14043 2322
rect 13991 2280 14043 2288
rect 14083 2280 14135 2332
rect 13991 2248 14043 2268
rect 13991 2216 13997 2248
rect 13997 2216 14035 2248
rect 14035 2216 14043 2248
rect 14083 2216 14135 2268
rect 13991 2174 14043 2204
rect 13991 2152 13997 2174
rect 13997 2152 14035 2174
rect 14035 2152 14043 2174
rect 14083 2152 14135 2204
rect 13991 2100 14043 2140
rect 13991 2088 13997 2100
rect 13997 2088 14035 2100
rect 14035 2088 14043 2100
rect 14083 2088 14135 2140
rect 13991 2066 13997 2075
rect 13997 2066 14035 2075
rect 14035 2066 14043 2075
rect 13991 2026 14043 2066
rect 13991 2023 13997 2026
rect 13997 2023 14035 2026
rect 14035 2023 14043 2026
rect 14083 2023 14135 2075
rect 13991 1992 13997 2010
rect 13997 1992 14035 2010
rect 14035 1992 14043 2010
rect 13991 1958 14043 1992
rect 14083 1958 14135 2010
rect 13991 1918 13997 1945
rect 13997 1918 14035 1945
rect 14035 1918 14043 1945
rect 13991 1893 14043 1918
rect 14083 1893 14135 1945
rect 13991 1878 14043 1880
rect 13991 1844 13997 1878
rect 13997 1844 14035 1878
rect 14035 1844 14043 1878
rect 13991 1828 14043 1844
rect 14083 1828 14135 1880
rect 13991 1804 14043 1815
rect 13991 1770 13997 1804
rect 13997 1770 14035 1804
rect 14035 1770 14043 1804
rect 13991 1763 14043 1770
rect 14083 1763 14135 1815
rect 13991 1730 14043 1750
rect 13991 1698 13997 1730
rect 13997 1698 14035 1730
rect 14035 1698 14043 1730
rect 14083 1698 14135 1750
rect 13991 1656 14043 1685
rect 13991 1633 13997 1656
rect 13997 1633 14035 1656
rect 14035 1633 14043 1656
rect 14083 1633 14135 1685
rect 13991 1582 14043 1620
rect 13991 1568 13997 1582
rect 13997 1568 14035 1582
rect 14035 1568 14043 1582
rect 14083 1568 14135 1620
rect 14350 4106 14356 4124
rect 14356 4106 14390 4124
rect 14390 4106 14402 4124
rect 14350 4072 14402 4106
rect 14422 4072 14428 4124
rect 14428 4072 14474 4124
rect 14494 4072 14546 4124
rect 14566 4072 14606 4124
rect 14606 4072 14618 4124
rect 14350 4033 14356 4059
rect 14356 4033 14390 4059
rect 14390 4033 14402 4059
rect 14350 4007 14402 4033
rect 14422 4007 14428 4059
rect 14428 4007 14474 4059
rect 14494 4007 14546 4059
rect 14566 4007 14606 4059
rect 14606 4007 14618 4059
rect 14350 3960 14356 3994
rect 14356 3960 14390 3994
rect 14390 3960 14402 3994
rect 14350 3942 14402 3960
rect 14422 3960 14428 3994
rect 14428 3960 14474 3994
rect 14494 3960 14546 3994
rect 14566 3960 14606 3994
rect 14606 3960 14618 3994
rect 14422 3952 14474 3960
rect 14422 3942 14428 3952
rect 14428 3942 14462 3952
rect 14462 3942 14474 3952
rect 14494 3942 14546 3960
rect 14566 3942 14618 3960
rect 14350 3921 14402 3929
rect 14350 3887 14356 3921
rect 14356 3887 14390 3921
rect 14390 3887 14402 3921
rect 14350 3877 14402 3887
rect 14422 3918 14428 3929
rect 14428 3918 14462 3929
rect 14462 3918 14474 3929
rect 14422 3880 14474 3918
rect 14422 3877 14428 3880
rect 14428 3877 14462 3880
rect 14462 3877 14474 3880
rect 14494 3921 14546 3929
rect 14494 3887 14500 3921
rect 14500 3887 14534 3921
rect 14534 3887 14546 3921
rect 14494 3877 14546 3887
rect 14566 3921 14618 3929
rect 14566 3887 14572 3921
rect 14572 3887 14606 3921
rect 14606 3887 14618 3921
rect 14566 3877 14618 3887
rect 14350 3848 14402 3864
rect 14350 3814 14356 3848
rect 14356 3814 14390 3848
rect 14390 3814 14402 3848
rect 14350 3812 14402 3814
rect 14422 3846 14428 3864
rect 14428 3846 14462 3864
rect 14462 3846 14474 3864
rect 14422 3812 14474 3846
rect 14494 3848 14546 3864
rect 14494 3814 14500 3848
rect 14500 3814 14534 3848
rect 14534 3814 14546 3848
rect 14494 3812 14546 3814
rect 14566 3848 14618 3864
rect 14566 3814 14572 3848
rect 14572 3814 14606 3848
rect 14606 3814 14618 3848
rect 14566 3812 14618 3814
rect 14350 3775 14402 3799
rect 14350 3747 14356 3775
rect 14356 3747 14390 3775
rect 14390 3747 14402 3775
rect 14422 3774 14428 3799
rect 14428 3774 14462 3799
rect 14462 3774 14474 3799
rect 14422 3747 14474 3774
rect 14494 3775 14546 3799
rect 14494 3747 14500 3775
rect 14500 3747 14534 3775
rect 14534 3747 14546 3775
rect 14566 3775 14618 3799
rect 14566 3747 14572 3775
rect 14572 3747 14606 3775
rect 14606 3747 14618 3775
rect 14350 3702 14402 3734
rect 14350 3682 14356 3702
rect 14356 3682 14390 3702
rect 14390 3682 14402 3702
rect 14422 3702 14428 3734
rect 14428 3702 14462 3734
rect 14462 3702 14474 3734
rect 14422 3682 14474 3702
rect 14494 3702 14546 3734
rect 14494 3682 14500 3702
rect 14500 3682 14534 3702
rect 14534 3682 14546 3702
rect 14566 3702 14618 3734
rect 14566 3682 14572 3702
rect 14572 3682 14606 3702
rect 14606 3682 14618 3702
rect 14350 3668 14356 3669
rect 14356 3668 14390 3669
rect 14390 3668 14402 3669
rect 14350 3629 14402 3668
rect 14350 3617 14356 3629
rect 14356 3617 14390 3629
rect 14390 3617 14402 3629
rect 14422 3664 14474 3669
rect 14422 3630 14428 3664
rect 14428 3630 14462 3664
rect 14462 3630 14474 3664
rect 14422 3617 14474 3630
rect 14494 3668 14500 3669
rect 14500 3668 14534 3669
rect 14534 3668 14546 3669
rect 14494 3629 14546 3668
rect 14494 3617 14500 3629
rect 14500 3617 14534 3629
rect 14534 3617 14546 3629
rect 14566 3668 14572 3669
rect 14572 3668 14606 3669
rect 14606 3668 14618 3669
rect 14566 3629 14618 3668
rect 14566 3617 14572 3629
rect 14572 3617 14606 3629
rect 14606 3617 14618 3629
rect 14350 3595 14356 3604
rect 14356 3595 14390 3604
rect 14390 3595 14402 3604
rect 14350 3556 14402 3595
rect 14350 3552 14356 3556
rect 14356 3552 14390 3556
rect 14390 3552 14402 3556
rect 14422 3592 14474 3604
rect 14422 3558 14428 3592
rect 14428 3558 14462 3592
rect 14462 3558 14474 3592
rect 14422 3552 14474 3558
rect 14494 3595 14500 3604
rect 14500 3595 14534 3604
rect 14534 3595 14546 3604
rect 14494 3556 14546 3595
rect 14494 3552 14500 3556
rect 14500 3552 14534 3556
rect 14534 3552 14546 3556
rect 14566 3595 14572 3604
rect 14572 3595 14606 3604
rect 14606 3595 14618 3604
rect 14566 3556 14618 3595
rect 14566 3552 14572 3556
rect 14572 3552 14606 3556
rect 14606 3552 14618 3556
rect 14350 3522 14356 3540
rect 14356 3522 14390 3540
rect 14390 3522 14402 3540
rect 14350 3488 14402 3522
rect 14422 3520 14474 3540
rect 14422 3488 14428 3520
rect 14428 3488 14462 3520
rect 14462 3488 14474 3520
rect 14494 3522 14500 3540
rect 14500 3522 14534 3540
rect 14534 3522 14546 3540
rect 14494 3488 14546 3522
rect 14566 3522 14572 3540
rect 14572 3522 14606 3540
rect 14606 3522 14618 3540
rect 14566 3488 14618 3522
rect 14350 3449 14356 3476
rect 14356 3449 14390 3476
rect 14390 3449 14402 3476
rect 14350 3424 14402 3449
rect 14422 3448 14474 3476
rect 14422 3424 14428 3448
rect 14428 3424 14462 3448
rect 14462 3424 14474 3448
rect 14494 3449 14500 3476
rect 14500 3449 14534 3476
rect 14534 3449 14546 3476
rect 14494 3424 14546 3449
rect 14566 3449 14572 3476
rect 14572 3449 14606 3476
rect 14606 3449 14618 3476
rect 14566 3424 14618 3449
rect 14350 3410 14402 3412
rect 14350 3376 14356 3410
rect 14356 3376 14390 3410
rect 14390 3376 14402 3410
rect 14350 3360 14402 3376
rect 14422 3376 14474 3412
rect 14422 3360 14428 3376
rect 14428 3360 14462 3376
rect 14462 3360 14474 3376
rect 14494 3410 14546 3412
rect 14494 3376 14500 3410
rect 14500 3376 14534 3410
rect 14534 3376 14546 3410
rect 14494 3360 14546 3376
rect 14566 3410 14618 3412
rect 14566 3376 14572 3410
rect 14572 3376 14606 3410
rect 14606 3376 14618 3410
rect 14566 3360 14618 3376
rect 14350 3337 14402 3348
rect 14350 3303 14356 3337
rect 14356 3303 14390 3337
rect 14390 3303 14402 3337
rect 14350 3296 14402 3303
rect 14422 3342 14428 3348
rect 14428 3342 14462 3348
rect 14462 3342 14474 3348
rect 14422 3304 14474 3342
rect 14422 3296 14428 3304
rect 14428 3296 14462 3304
rect 14462 3296 14474 3304
rect 14494 3337 14546 3348
rect 14494 3303 14500 3337
rect 14500 3303 14534 3337
rect 14534 3303 14546 3337
rect 14494 3296 14546 3303
rect 14566 3337 14618 3348
rect 14566 3303 14572 3337
rect 14572 3303 14606 3337
rect 14606 3303 14618 3337
rect 14566 3296 14618 3303
rect 14350 3264 14402 3284
rect 14350 3232 14356 3264
rect 14356 3232 14390 3264
rect 14390 3232 14402 3264
rect 14422 3270 14428 3284
rect 14428 3270 14462 3284
rect 14462 3270 14474 3284
rect 14422 3232 14474 3270
rect 14494 3264 14546 3284
rect 14494 3232 14500 3264
rect 14500 3232 14534 3264
rect 14534 3232 14546 3264
rect 14566 3264 14618 3284
rect 14566 3232 14572 3264
rect 14572 3232 14606 3264
rect 14606 3232 14618 3264
rect 14350 3191 14402 3220
rect 14350 3168 14356 3191
rect 14356 3168 14390 3191
rect 14390 3168 14402 3191
rect 14422 3198 14428 3220
rect 14428 3198 14462 3220
rect 14462 3198 14474 3220
rect 14422 3168 14474 3198
rect 14494 3191 14546 3220
rect 14494 3168 14500 3191
rect 14500 3168 14534 3191
rect 14534 3168 14546 3191
rect 14566 3191 14618 3220
rect 14566 3168 14572 3191
rect 14572 3168 14606 3191
rect 14606 3168 14618 3191
rect 14350 3118 14402 3156
rect 14350 3104 14356 3118
rect 14356 3104 14390 3118
rect 14390 3104 14402 3118
rect 14422 3126 14428 3156
rect 14428 3126 14462 3156
rect 14462 3126 14474 3156
rect 14422 3104 14474 3126
rect 14494 3118 14546 3156
rect 14494 3104 14500 3118
rect 14500 3104 14534 3118
rect 14534 3104 14546 3118
rect 14566 3118 14618 3156
rect 14566 3104 14572 3118
rect 14572 3104 14606 3118
rect 14606 3104 14618 3118
rect 14350 3084 14356 3092
rect 14356 3084 14390 3092
rect 14390 3084 14402 3092
rect 14350 3045 14402 3084
rect 14350 3040 14356 3045
rect 14356 3040 14390 3045
rect 14390 3040 14402 3045
rect 14422 3088 14474 3092
rect 14422 3054 14428 3088
rect 14428 3054 14462 3088
rect 14462 3054 14474 3088
rect 14422 3040 14474 3054
rect 14494 3084 14500 3092
rect 14500 3084 14534 3092
rect 14534 3084 14546 3092
rect 14494 3045 14546 3084
rect 14494 3040 14500 3045
rect 14500 3040 14534 3045
rect 14534 3040 14546 3045
rect 14566 3084 14572 3092
rect 14572 3084 14606 3092
rect 14606 3084 14618 3092
rect 14566 3045 14618 3084
rect 14566 3040 14572 3045
rect 14572 3040 14606 3045
rect 14606 3040 14618 3045
rect 14350 3011 14356 3028
rect 14356 3011 14390 3028
rect 14390 3011 14402 3028
rect 14350 2976 14402 3011
rect 14422 3016 14474 3028
rect 14422 2982 14428 3016
rect 14428 2982 14462 3016
rect 14462 2982 14474 3016
rect 14422 2976 14474 2982
rect 14494 3011 14500 3028
rect 14500 3011 14534 3028
rect 14534 3011 14546 3028
rect 14494 2976 14546 3011
rect 14566 3011 14572 3028
rect 14572 3011 14606 3028
rect 14606 3011 14618 3028
rect 14566 2976 14618 3011
rect 14350 2938 14356 2964
rect 14356 2938 14390 2964
rect 14390 2938 14402 2964
rect 14350 2912 14402 2938
rect 14422 2944 14474 2964
rect 14422 2912 14428 2944
rect 14428 2912 14462 2944
rect 14462 2912 14474 2944
rect 14494 2938 14500 2964
rect 14500 2938 14534 2964
rect 14534 2938 14546 2964
rect 14494 2912 14546 2938
rect 14566 2938 14572 2964
rect 14572 2938 14606 2964
rect 14606 2938 14618 2964
rect 14566 2912 14618 2938
rect 14350 2899 14402 2900
rect 14350 2865 14356 2899
rect 14356 2865 14390 2899
rect 14390 2865 14402 2899
rect 14350 2848 14402 2865
rect 14422 2872 14474 2900
rect 14422 2848 14428 2872
rect 14428 2848 14462 2872
rect 14462 2848 14474 2872
rect 14494 2899 14546 2900
rect 14494 2865 14500 2899
rect 14500 2865 14534 2899
rect 14534 2865 14546 2899
rect 14494 2848 14546 2865
rect 14566 2899 14618 2900
rect 14566 2865 14572 2899
rect 14572 2865 14606 2899
rect 14606 2865 14618 2899
rect 14566 2848 14618 2865
rect 14350 2826 14402 2836
rect 14350 2792 14356 2826
rect 14356 2792 14390 2826
rect 14390 2792 14402 2826
rect 14350 2784 14402 2792
rect 14422 2800 14474 2836
rect 14422 2784 14428 2800
rect 14428 2784 14462 2800
rect 14462 2784 14474 2800
rect 14494 2826 14546 2836
rect 14494 2792 14500 2826
rect 14500 2792 14534 2826
rect 14534 2792 14546 2826
rect 14494 2784 14546 2792
rect 14566 2826 14618 2836
rect 14566 2792 14572 2826
rect 14572 2792 14606 2826
rect 14606 2792 14618 2826
rect 14566 2784 14618 2792
rect 14350 2753 14402 2772
rect 14350 2720 14356 2753
rect 14356 2720 14390 2753
rect 14390 2720 14402 2753
rect 14422 2766 14428 2772
rect 14428 2766 14462 2772
rect 14462 2766 14474 2772
rect 14422 2728 14474 2766
rect 14422 2720 14428 2728
rect 14428 2720 14462 2728
rect 14462 2720 14474 2728
rect 14494 2753 14546 2772
rect 14494 2720 14500 2753
rect 14500 2720 14534 2753
rect 14534 2720 14546 2753
rect 14566 2753 14618 2772
rect 14566 2720 14572 2753
rect 14572 2720 14606 2753
rect 14606 2720 14618 2753
rect 14350 2680 14402 2708
rect 14350 2656 14356 2680
rect 14356 2656 14390 2680
rect 14390 2656 14402 2680
rect 14422 2694 14428 2708
rect 14428 2694 14462 2708
rect 14462 2694 14474 2708
rect 14422 2656 14474 2694
rect 14494 2680 14546 2708
rect 14494 2656 14500 2680
rect 14500 2656 14534 2680
rect 14534 2656 14546 2680
rect 14566 2680 14618 2708
rect 14566 2656 14572 2680
rect 14572 2656 14606 2680
rect 14606 2656 14618 2680
rect 14350 2607 14402 2644
rect 14350 2592 14356 2607
rect 14356 2592 14390 2607
rect 14390 2592 14402 2607
rect 14422 2622 14428 2644
rect 14428 2622 14462 2644
rect 14462 2622 14474 2644
rect 14422 2592 14474 2622
rect 14494 2607 14546 2644
rect 14494 2592 14500 2607
rect 14500 2592 14534 2607
rect 14534 2592 14546 2607
rect 14566 2607 14618 2644
rect 14566 2592 14572 2607
rect 14572 2592 14606 2607
rect 14606 2592 14618 2607
rect 14350 2573 14356 2580
rect 14356 2573 14390 2580
rect 14390 2573 14402 2580
rect 14350 2534 14402 2573
rect 14350 2528 14356 2534
rect 14356 2528 14390 2534
rect 14390 2528 14402 2534
rect 14422 2550 14428 2580
rect 14428 2550 14462 2580
rect 14462 2550 14474 2580
rect 14422 2528 14474 2550
rect 14494 2573 14500 2580
rect 14500 2573 14534 2580
rect 14534 2573 14546 2580
rect 14494 2534 14546 2573
rect 14494 2528 14500 2534
rect 14500 2528 14534 2534
rect 14534 2528 14546 2534
rect 14566 2573 14572 2580
rect 14572 2573 14606 2580
rect 14606 2573 14618 2580
rect 14566 2534 14618 2573
rect 14566 2528 14572 2534
rect 14572 2528 14606 2534
rect 14606 2528 14618 2534
rect 14350 2500 14356 2516
rect 14356 2500 14390 2516
rect 14390 2500 14402 2516
rect 14350 2464 14402 2500
rect 14422 2512 14474 2516
rect 14422 2478 14428 2512
rect 14428 2478 14462 2512
rect 14462 2478 14474 2512
rect 14422 2464 14474 2478
rect 14494 2500 14500 2516
rect 14500 2500 14534 2516
rect 14534 2500 14546 2516
rect 14494 2464 14546 2500
rect 14566 2500 14572 2516
rect 14572 2500 14606 2516
rect 14606 2500 14618 2516
rect 14566 2464 14618 2500
rect 14350 2427 14356 2452
rect 14356 2427 14390 2452
rect 14390 2427 14402 2452
rect 14350 2400 14402 2427
rect 14422 2440 14474 2452
rect 14422 2406 14428 2440
rect 14428 2406 14462 2440
rect 14462 2406 14474 2440
rect 14422 2400 14474 2406
rect 14494 2427 14500 2452
rect 14500 2427 14534 2452
rect 14534 2427 14546 2452
rect 14494 2400 14546 2427
rect 14566 2427 14572 2452
rect 14572 2427 14606 2452
rect 14606 2427 14618 2452
rect 14566 2400 14618 2427
rect 14350 2354 14356 2388
rect 14356 2354 14390 2388
rect 14390 2354 14402 2388
rect 14350 2336 14402 2354
rect 14422 2368 14474 2388
rect 14422 2336 14428 2368
rect 14428 2336 14462 2368
rect 14462 2336 14474 2368
rect 14494 2354 14500 2388
rect 14500 2354 14534 2388
rect 14534 2354 14546 2388
rect 14494 2336 14546 2354
rect 14566 2354 14572 2388
rect 14572 2354 14606 2388
rect 14606 2354 14618 2388
rect 14566 2336 14618 2354
rect 14350 2315 14402 2324
rect 14350 2281 14356 2315
rect 14356 2281 14390 2315
rect 14390 2281 14402 2315
rect 14350 2272 14402 2281
rect 14422 2296 14474 2324
rect 14422 2272 14428 2296
rect 14428 2272 14462 2296
rect 14462 2272 14474 2296
rect 14494 2315 14546 2324
rect 14494 2281 14500 2315
rect 14500 2281 14534 2315
rect 14534 2281 14546 2315
rect 14494 2272 14546 2281
rect 14566 2315 14618 2324
rect 14566 2281 14572 2315
rect 14572 2281 14606 2315
rect 14606 2281 14618 2315
rect 14566 2272 14618 2281
rect 14350 2242 14402 2260
rect 14350 2208 14356 2242
rect 14356 2208 14390 2242
rect 14390 2208 14402 2242
rect 14422 2224 14474 2260
rect 14422 2208 14428 2224
rect 14428 2208 14462 2224
rect 14462 2208 14474 2224
rect 14494 2242 14546 2260
rect 14494 2208 14500 2242
rect 14500 2208 14534 2242
rect 14534 2208 14546 2242
rect 14566 2242 14618 2260
rect 14566 2208 14572 2242
rect 14572 2208 14606 2242
rect 14606 2208 14618 2242
rect 14350 2169 14402 2196
rect 14350 2144 14356 2169
rect 14356 2144 14390 2169
rect 14390 2144 14402 2169
rect 14422 2190 14428 2196
rect 14428 2190 14462 2196
rect 14462 2190 14474 2196
rect 14422 2152 14474 2190
rect 14422 2144 14428 2152
rect 14428 2144 14462 2152
rect 14462 2144 14474 2152
rect 14494 2169 14546 2196
rect 14494 2144 14500 2169
rect 14500 2144 14534 2169
rect 14534 2144 14546 2169
rect 14566 2169 14618 2196
rect 14566 2144 14572 2169
rect 14572 2144 14606 2169
rect 14606 2144 14618 2169
rect 14350 2096 14402 2132
rect 14350 2080 14356 2096
rect 14356 2080 14390 2096
rect 14390 2080 14402 2096
rect 14422 2118 14428 2132
rect 14428 2118 14462 2132
rect 14462 2118 14474 2132
rect 14422 2080 14474 2118
rect 14494 2096 14546 2132
rect 14494 2080 14500 2096
rect 14500 2080 14534 2096
rect 14534 2080 14546 2096
rect 14566 2096 14618 2132
rect 14566 2080 14572 2096
rect 14572 2080 14606 2096
rect 14606 2080 14618 2096
rect 14350 2062 14356 2068
rect 14356 2062 14390 2068
rect 14390 2062 14402 2068
rect 14350 2023 14402 2062
rect 14350 2016 14356 2023
rect 14356 2016 14390 2023
rect 14390 2016 14402 2023
rect 14422 2046 14428 2068
rect 14428 2046 14462 2068
rect 14462 2046 14474 2068
rect 14422 2016 14474 2046
rect 14494 2062 14500 2068
rect 14500 2062 14534 2068
rect 14534 2062 14546 2068
rect 14494 2023 14546 2062
rect 14494 2016 14500 2023
rect 14500 2016 14534 2023
rect 14534 2016 14546 2023
rect 14566 2062 14572 2068
rect 14572 2062 14606 2068
rect 14606 2062 14618 2068
rect 14566 2023 14618 2062
rect 14566 2016 14572 2023
rect 14572 2016 14606 2023
rect 14606 2016 14618 2023
rect 14350 1989 14356 2004
rect 14356 1989 14390 2004
rect 14390 1989 14402 2004
rect 14350 1952 14402 1989
rect 14422 1974 14428 2004
rect 14428 1974 14462 2004
rect 14462 1974 14474 2004
rect 14422 1952 14474 1974
rect 14494 1989 14500 2004
rect 14500 1989 14534 2004
rect 14534 1989 14546 2004
rect 14494 1952 14546 1989
rect 14566 1989 14572 2004
rect 14572 1989 14606 2004
rect 14606 1989 14618 2004
rect 14566 1952 14618 1989
rect 14350 1916 14356 1940
rect 14356 1916 14390 1940
rect 14390 1916 14402 1940
rect 14350 1888 14402 1916
rect 14422 1936 14474 1940
rect 14422 1902 14428 1936
rect 14428 1902 14462 1936
rect 14462 1902 14474 1936
rect 14422 1888 14474 1902
rect 14494 1916 14500 1940
rect 14500 1916 14534 1940
rect 14534 1916 14546 1940
rect 14494 1888 14546 1916
rect 14566 1916 14572 1940
rect 14572 1916 14606 1940
rect 14606 1916 14618 1940
rect 14566 1888 14618 1916
rect 14350 1843 14356 1876
rect 14356 1843 14390 1876
rect 14390 1843 14402 1876
rect 14350 1824 14402 1843
rect 14422 1864 14474 1876
rect 14422 1830 14428 1864
rect 14428 1830 14462 1864
rect 14462 1830 14474 1864
rect 14422 1824 14474 1830
rect 14494 1843 14500 1876
rect 14500 1843 14534 1876
rect 14534 1843 14546 1876
rect 14494 1824 14546 1843
rect 14566 1843 14572 1876
rect 14572 1843 14606 1876
rect 14606 1843 14618 1876
rect 14566 1824 14618 1843
rect 14350 1804 14402 1812
rect 14350 1770 14356 1804
rect 14356 1770 14390 1804
rect 14390 1770 14402 1804
rect 14350 1760 14402 1770
rect 14422 1792 14474 1812
rect 14422 1760 14428 1792
rect 14428 1760 14462 1792
rect 14462 1760 14474 1792
rect 14494 1804 14546 1812
rect 14494 1770 14500 1804
rect 14500 1770 14534 1804
rect 14534 1770 14546 1804
rect 14494 1760 14546 1770
rect 14566 1804 14618 1812
rect 14566 1770 14572 1804
rect 14572 1770 14606 1804
rect 14606 1770 14618 1804
rect 14566 1760 14618 1770
rect 14350 1731 14402 1748
rect 14350 1697 14356 1731
rect 14356 1697 14390 1731
rect 14390 1697 14402 1731
rect 14350 1696 14402 1697
rect 14422 1720 14474 1748
rect 14422 1696 14428 1720
rect 14428 1696 14462 1720
rect 14462 1696 14474 1720
rect 14494 1731 14546 1748
rect 14494 1697 14500 1731
rect 14500 1697 14534 1731
rect 14534 1697 14546 1731
rect 14494 1696 14546 1697
rect 14566 1731 14618 1748
rect 14566 1697 14572 1731
rect 14572 1697 14606 1731
rect 14606 1697 14618 1731
rect 14566 1696 14618 1697
rect 14350 1657 14402 1684
rect 14350 1632 14356 1657
rect 14356 1632 14390 1657
rect 14390 1632 14402 1657
rect 14422 1648 14474 1684
rect 14422 1632 14428 1648
rect 14428 1632 14462 1648
rect 14462 1632 14474 1648
rect 14494 1658 14546 1684
rect 14494 1632 14500 1658
rect 14500 1632 14534 1658
rect 14534 1632 14546 1658
rect 14566 1658 14618 1684
rect 14566 1632 14572 1658
rect 14572 1632 14606 1658
rect 14606 1632 14618 1658
rect 14350 1583 14402 1620
rect 14350 1568 14356 1583
rect 14356 1568 14390 1583
rect 14390 1568 14402 1583
rect 14422 1614 14428 1620
rect 14428 1614 14462 1620
rect 14462 1614 14474 1620
rect 14422 1576 14474 1614
rect 14422 1568 14428 1576
rect 14428 1568 14462 1576
rect 14462 1568 14474 1576
rect 14494 1585 14546 1620
rect 14494 1568 14500 1585
rect 14500 1568 14534 1585
rect 14534 1568 14546 1585
rect 14566 1585 14618 1620
rect 14566 1568 14572 1585
rect 14572 1568 14606 1585
rect 14606 1568 14618 1585
rect 518 1513 570 1530
rect 518 1479 529 1513
rect 529 1479 563 1513
rect 563 1479 570 1513
rect 518 1478 570 1479
rect 590 1513 642 1530
rect 590 1479 601 1513
rect 601 1479 635 1513
rect 635 1479 642 1513
rect 590 1478 642 1479
rect 662 1478 674 1530
rect 674 1478 714 1530
rect 734 1478 780 1530
rect 780 1478 786 1530
rect 518 1440 570 1465
rect 518 1413 529 1440
rect 529 1413 563 1440
rect 563 1413 570 1440
rect 590 1440 642 1465
rect 590 1413 601 1440
rect 601 1413 635 1440
rect 635 1413 642 1440
rect 662 1413 674 1465
rect 674 1413 714 1465
rect 734 1413 780 1465
rect 780 1413 786 1465
rect 518 1367 570 1400
rect 518 1348 529 1367
rect 529 1348 563 1367
rect 563 1348 570 1367
rect 590 1367 642 1400
rect 590 1348 601 1367
rect 601 1348 635 1367
rect 635 1348 642 1367
rect 662 1348 674 1400
rect 674 1348 714 1400
rect 734 1348 780 1400
rect 780 1348 786 1400
rect 518 1333 529 1335
rect 529 1333 563 1335
rect 563 1333 570 1335
rect 518 1294 570 1333
rect 518 1283 529 1294
rect 529 1283 563 1294
rect 563 1283 570 1294
rect 590 1333 601 1335
rect 601 1333 635 1335
rect 635 1333 642 1335
rect 590 1294 642 1333
rect 590 1283 601 1294
rect 601 1283 635 1294
rect 635 1283 642 1294
rect 662 1283 674 1335
rect 674 1283 714 1335
rect 734 1283 780 1335
rect 780 1283 786 1335
rect 518 1260 529 1270
rect 529 1260 563 1270
rect 563 1260 570 1270
rect 518 1221 570 1260
rect 518 1218 529 1221
rect 529 1218 563 1221
rect 563 1218 570 1221
rect 590 1260 601 1270
rect 601 1260 635 1270
rect 635 1260 642 1270
rect 590 1221 642 1260
rect 590 1218 601 1221
rect 601 1218 635 1221
rect 635 1218 642 1221
rect 662 1218 674 1270
rect 674 1218 714 1270
rect 734 1218 780 1270
rect 780 1218 786 1270
rect 518 1187 529 1205
rect 529 1187 563 1205
rect 563 1187 570 1205
rect 518 1153 570 1187
rect 590 1187 601 1205
rect 601 1187 635 1205
rect 635 1187 642 1205
rect 590 1153 642 1187
rect 662 1153 674 1205
rect 674 1153 714 1205
rect 734 1153 780 1205
rect 780 1153 786 1205
rect 518 1114 529 1140
rect 529 1114 563 1140
rect 563 1114 570 1140
rect 518 1088 570 1114
rect 590 1114 601 1140
rect 601 1114 635 1140
rect 635 1114 642 1140
rect 590 1088 642 1114
rect 662 1088 674 1140
rect 674 1088 714 1140
rect 734 1088 780 1140
rect 780 1088 786 1140
rect 518 1041 529 1075
rect 529 1041 563 1075
rect 563 1041 570 1075
rect 518 1023 570 1041
rect 590 1041 601 1075
rect 601 1041 635 1075
rect 635 1041 642 1075
rect 590 1023 642 1041
rect 662 1023 674 1075
rect 674 1023 714 1075
rect 734 1023 780 1075
rect 780 1023 786 1075
rect 518 1002 570 1010
rect 518 968 529 1002
rect 529 968 563 1002
rect 563 968 570 1002
rect 518 958 570 968
rect 590 1002 642 1010
rect 590 968 601 1002
rect 601 968 635 1002
rect 635 968 642 1002
rect 590 958 642 968
rect 662 958 674 1010
rect 674 958 714 1010
rect 734 958 780 1010
rect 780 958 786 1010
rect 518 929 570 945
rect 518 895 529 929
rect 529 895 563 929
rect 563 895 570 929
rect 518 893 570 895
rect 590 929 642 945
rect 590 895 601 929
rect 601 895 635 929
rect 635 895 642 929
rect 590 893 642 895
rect 662 894 674 945
rect 674 894 714 945
rect 734 894 780 945
rect 662 893 714 894
rect 734 893 746 894
rect 746 893 780 894
rect 780 893 786 945
rect 518 828 570 880
rect 590 828 642 880
rect 662 828 714 880
rect 734 828 786 880
<< metal2 >>
rect 518 4456 786 4462
rect 570 4404 590 4456
rect 642 4404 662 4456
rect 714 4404 734 4456
rect 518 4390 786 4404
rect 570 4338 590 4390
rect 642 4338 662 4390
rect 714 4338 734 4390
rect 518 4325 786 4338
rect 570 4273 590 4325
rect 642 4273 662 4325
rect 714 4273 734 4325
rect 518 4260 786 4273
rect 570 4208 590 4260
rect 642 4208 662 4260
rect 714 4208 734 4260
rect 518 4195 786 4208
rect 570 4143 590 4195
rect 642 4143 662 4195
rect 714 4143 734 4195
rect 518 4130 786 4143
rect 570 4078 590 4130
rect 642 4078 662 4130
rect 714 4078 734 4130
rect 518 4065 786 4078
rect 570 4013 590 4065
rect 642 4013 662 4065
rect 714 4013 734 4065
rect 518 4000 786 4013
rect 570 3948 590 4000
rect 642 3948 662 4000
rect 714 3948 734 4000
rect 518 3935 786 3948
rect 570 3883 590 3935
rect 642 3883 662 3935
rect 714 3883 734 3935
rect 518 3870 786 3883
rect 570 3818 590 3870
rect 642 3818 662 3870
rect 714 3818 734 3870
rect 518 3805 786 3818
rect 570 3753 590 3805
rect 642 3753 662 3805
rect 714 3753 734 3805
rect 518 3740 786 3753
rect 570 3688 590 3740
rect 642 3688 662 3740
rect 714 3688 734 3740
rect 518 3675 786 3688
rect 570 3623 590 3675
rect 642 3623 662 3675
rect 714 3623 734 3675
rect 518 3610 786 3623
rect 570 3558 590 3610
rect 642 3558 662 3610
rect 714 3558 734 3610
rect 518 3545 786 3558
rect 570 3493 590 3545
rect 642 3493 662 3545
rect 714 3493 734 3545
rect 518 3480 786 3493
rect 570 3428 590 3480
rect 642 3428 662 3480
rect 714 3428 734 3480
rect 518 3415 786 3428
rect 570 3363 590 3415
rect 642 3363 662 3415
rect 714 3363 734 3415
rect 518 3350 786 3363
rect 570 3298 590 3350
rect 642 3298 662 3350
rect 714 3298 734 3350
rect 518 3285 786 3298
rect 570 3233 590 3285
rect 642 3233 662 3285
rect 714 3233 734 3285
rect 518 3220 786 3233
rect 570 3168 590 3220
rect 642 3168 662 3220
rect 714 3168 734 3220
rect 518 3155 786 3168
rect 570 3103 590 3155
rect 642 3103 662 3155
rect 714 3103 734 3155
rect 518 3090 786 3103
rect 570 3038 590 3090
rect 642 3038 662 3090
rect 714 3038 734 3090
rect 518 3025 786 3038
rect 570 2973 590 3025
rect 642 2973 662 3025
rect 714 2973 734 3025
rect 518 2960 786 2973
rect 570 2908 590 2960
rect 642 2908 662 2960
rect 714 2908 734 2960
rect 518 2895 786 2908
rect 570 2843 590 2895
rect 642 2843 662 2895
rect 714 2843 734 2895
rect 518 2830 786 2843
rect 570 2778 590 2830
rect 642 2778 662 2830
rect 714 2778 734 2830
rect 518 2765 786 2778
rect 570 2713 590 2765
rect 642 2713 662 2765
rect 714 2713 734 2765
rect 518 2700 786 2713
rect 570 2648 590 2700
rect 642 2648 662 2700
rect 714 2648 734 2700
rect 518 2635 786 2648
rect 570 2583 590 2635
rect 642 2583 662 2635
rect 714 2583 734 2635
rect 518 2570 786 2583
rect 570 2518 590 2570
rect 642 2518 662 2570
rect 714 2518 734 2570
rect 518 2505 786 2518
rect 570 2453 590 2505
rect 642 2453 662 2505
rect 714 2453 734 2505
rect 518 2440 786 2453
rect 570 2388 590 2440
rect 642 2388 662 2440
rect 714 2388 734 2440
rect 518 2375 786 2388
rect 570 2323 590 2375
rect 642 2323 662 2375
rect 714 2323 734 2375
rect 518 2310 786 2323
rect 570 2258 590 2310
rect 642 2258 662 2310
rect 714 2258 734 2310
rect 518 2245 786 2258
rect 570 2193 590 2245
rect 642 2193 662 2245
rect 714 2193 734 2245
rect 518 2180 786 2193
rect 570 2128 590 2180
rect 642 2128 662 2180
rect 714 2128 734 2180
rect 518 2115 786 2128
rect 570 2063 590 2115
rect 642 2063 662 2115
rect 714 2063 734 2115
rect 518 2050 786 2063
rect 570 1998 590 2050
rect 642 1998 662 2050
rect 714 1998 734 2050
rect 518 1985 786 1998
rect 570 1933 590 1985
rect 642 1933 662 1985
rect 714 1933 734 1985
rect 518 1920 786 1933
rect 570 1868 590 1920
rect 642 1868 662 1920
rect 714 1868 734 1920
rect 518 1855 786 1868
rect 570 1803 590 1855
rect 642 1803 662 1855
rect 714 1803 734 1855
rect 518 1790 786 1803
rect 570 1738 590 1790
rect 642 1738 662 1790
rect 714 1738 734 1790
rect 518 1725 786 1738
rect 570 1673 590 1725
rect 642 1673 662 1725
rect 714 1673 734 1725
rect 518 1660 786 1673
rect 570 1608 590 1660
rect 642 1608 662 1660
rect 714 1608 734 1660
rect 518 1595 786 1608
rect 570 1543 590 1595
rect 642 1543 662 1595
rect 714 1543 734 1595
rect 1061 4119 1251 4125
rect 1061 4067 1066 4119
rect 1118 4067 1130 4119
rect 1182 4067 1194 4119
rect 1246 4067 1251 4119
rect 1061 4054 1251 4067
rect 1061 4002 1066 4054
rect 1118 4002 1130 4054
rect 1182 4002 1194 4054
rect 1246 4002 1251 4054
rect 1061 3989 1251 4002
rect 1061 3937 1066 3989
rect 1118 3937 1130 3989
rect 1182 3937 1194 3989
rect 1246 3937 1251 3989
rect 1061 3924 1251 3937
rect 1061 1568 1066 3924
rect 1246 1568 1251 3924
rect 1061 1562 1251 1568
rect 1557 4124 1747 4130
rect 1557 4072 1562 4124
rect 1614 4072 1626 4124
rect 1678 4072 1690 4124
rect 1742 4072 1747 4124
rect 1557 4059 1747 4072
rect 1557 4007 1562 4059
rect 1614 4007 1626 4059
rect 1678 4007 1690 4059
rect 1742 4007 1747 4059
rect 1557 3994 1747 4007
rect 1557 3942 1562 3994
rect 1614 3942 1626 3994
rect 1678 3942 1690 3994
rect 1742 3942 1747 3994
rect 1557 3929 1747 3942
rect 1557 3877 1562 3929
rect 1614 3877 1626 3929
rect 1678 3877 1690 3929
rect 1742 3877 1747 3929
rect 1557 3864 1747 3877
rect 1557 3812 1562 3864
rect 1614 3812 1626 3864
rect 1678 3812 1690 3864
rect 1742 3812 1747 3864
rect 1557 3799 1747 3812
rect 1557 3747 1562 3799
rect 1614 3747 1626 3799
rect 1678 3747 1690 3799
rect 1742 3747 1747 3799
rect 1557 3734 1747 3747
rect 1557 3682 1562 3734
rect 1614 3682 1626 3734
rect 1678 3682 1690 3734
rect 1742 3682 1747 3734
rect 1557 3669 1747 3682
rect 1557 3617 1562 3669
rect 1614 3617 1626 3669
rect 1678 3617 1690 3669
rect 1742 3617 1747 3669
rect 1557 3604 1747 3617
rect 1557 1568 1562 3604
rect 1742 1568 1747 3604
rect 1557 1562 1747 1568
rect 2053 4119 2243 4125
rect 2053 4067 2058 4119
rect 2110 4067 2122 4119
rect 2174 4067 2186 4119
rect 2238 4067 2243 4119
rect 2053 4054 2243 4067
rect 2053 4002 2058 4054
rect 2110 4002 2122 4054
rect 2174 4002 2186 4054
rect 2238 4002 2243 4054
rect 2053 3989 2243 4002
rect 2053 3937 2058 3989
rect 2110 3937 2122 3989
rect 2174 3937 2186 3989
rect 2238 3937 2243 3989
rect 2053 3924 2243 3937
rect 2053 1568 2058 3924
rect 2238 1568 2243 3924
rect 2053 1562 2243 1568
rect 2549 4124 2739 4130
rect 2549 4072 2554 4124
rect 2606 4072 2618 4124
rect 2670 4072 2682 4124
rect 2734 4072 2739 4124
rect 2549 4059 2739 4072
rect 2549 4007 2554 4059
rect 2606 4007 2618 4059
rect 2670 4007 2682 4059
rect 2734 4007 2739 4059
rect 2549 3994 2739 4007
rect 2549 3942 2554 3994
rect 2606 3942 2618 3994
rect 2670 3942 2682 3994
rect 2734 3942 2739 3994
rect 2549 3929 2739 3942
rect 2549 3877 2554 3929
rect 2606 3877 2618 3929
rect 2670 3877 2682 3929
rect 2734 3877 2739 3929
rect 2549 3864 2739 3877
rect 2549 3812 2554 3864
rect 2606 3812 2618 3864
rect 2670 3812 2682 3864
rect 2734 3812 2739 3864
rect 2549 3799 2739 3812
rect 2549 3747 2554 3799
rect 2606 3747 2618 3799
rect 2670 3747 2682 3799
rect 2734 3747 2739 3799
rect 2549 3734 2739 3747
rect 2549 3682 2554 3734
rect 2606 3682 2618 3734
rect 2670 3682 2682 3734
rect 2734 3682 2739 3734
rect 2549 3669 2739 3682
rect 2549 3617 2554 3669
rect 2606 3617 2618 3669
rect 2670 3617 2682 3669
rect 2734 3617 2739 3669
rect 2549 3604 2739 3617
rect 2549 1568 2554 3604
rect 2734 1568 2739 3604
rect 2549 1562 2739 1568
rect 3045 4119 3235 4125
rect 3045 4067 3050 4119
rect 3102 4067 3114 4119
rect 3166 4067 3178 4119
rect 3230 4067 3235 4119
rect 3045 4054 3235 4067
rect 3045 4002 3050 4054
rect 3102 4002 3114 4054
rect 3166 4002 3178 4054
rect 3230 4002 3235 4054
rect 3045 3989 3235 4002
rect 3045 3937 3050 3989
rect 3102 3937 3114 3989
rect 3166 3937 3178 3989
rect 3230 3937 3235 3989
rect 3045 3924 3235 3937
rect 3045 1568 3050 3924
rect 3230 1568 3235 3924
rect 3045 1562 3235 1568
rect 3541 4124 3731 4130
rect 3541 4072 3546 4124
rect 3598 4072 3610 4124
rect 3662 4072 3674 4124
rect 3726 4072 3731 4124
rect 3541 4059 3731 4072
rect 3541 4007 3546 4059
rect 3598 4007 3610 4059
rect 3662 4007 3674 4059
rect 3726 4007 3731 4059
rect 3541 3994 3731 4007
rect 3541 3942 3546 3994
rect 3598 3942 3610 3994
rect 3662 3942 3674 3994
rect 3726 3942 3731 3994
rect 3541 3929 3731 3942
rect 3541 3877 3546 3929
rect 3598 3877 3610 3929
rect 3662 3877 3674 3929
rect 3726 3877 3731 3929
rect 3541 3864 3731 3877
rect 3541 3812 3546 3864
rect 3598 3812 3610 3864
rect 3662 3812 3674 3864
rect 3726 3812 3731 3864
rect 3541 3799 3731 3812
rect 3541 3747 3546 3799
rect 3598 3747 3610 3799
rect 3662 3747 3674 3799
rect 3726 3747 3731 3799
rect 3541 3734 3731 3747
rect 3541 3682 3546 3734
rect 3598 3682 3610 3734
rect 3662 3682 3674 3734
rect 3726 3682 3731 3734
rect 3541 3669 3731 3682
rect 3541 3617 3546 3669
rect 3598 3617 3610 3669
rect 3662 3617 3674 3669
rect 3726 3617 3731 3669
rect 3541 3604 3731 3617
rect 3541 1568 3546 3604
rect 3726 1568 3731 3604
rect 3541 1562 3731 1568
rect 4037 4119 4227 4125
rect 4037 4067 4042 4119
rect 4094 4067 4106 4119
rect 4158 4067 4170 4119
rect 4222 4067 4227 4119
rect 4037 4054 4227 4067
rect 4037 4002 4042 4054
rect 4094 4002 4106 4054
rect 4158 4002 4170 4054
rect 4222 4002 4227 4054
rect 4037 3989 4227 4002
rect 4037 3937 4042 3989
rect 4094 3937 4106 3989
rect 4158 3937 4170 3989
rect 4222 3937 4227 3989
rect 4037 3924 4227 3937
rect 4037 1568 4042 3924
rect 4222 1568 4227 3924
rect 4037 1562 4227 1568
rect 4533 4124 4723 4130
rect 4533 4072 4538 4124
rect 4590 4072 4602 4124
rect 4654 4072 4666 4124
rect 4718 4072 4723 4124
rect 4533 4059 4723 4072
rect 4533 4007 4538 4059
rect 4590 4007 4602 4059
rect 4654 4007 4666 4059
rect 4718 4007 4723 4059
rect 4533 3994 4723 4007
rect 4533 3942 4538 3994
rect 4590 3942 4602 3994
rect 4654 3942 4666 3994
rect 4718 3942 4723 3994
rect 4533 3929 4723 3942
rect 4533 3877 4538 3929
rect 4590 3877 4602 3929
rect 4654 3877 4666 3929
rect 4718 3877 4723 3929
rect 4533 3864 4723 3877
rect 4533 3812 4538 3864
rect 4590 3812 4602 3864
rect 4654 3812 4666 3864
rect 4718 3812 4723 3864
rect 4533 3799 4723 3812
rect 4533 3747 4538 3799
rect 4590 3747 4602 3799
rect 4654 3747 4666 3799
rect 4718 3747 4723 3799
rect 4533 3734 4723 3747
rect 4533 3682 4538 3734
rect 4590 3682 4602 3734
rect 4654 3682 4666 3734
rect 4718 3682 4723 3734
rect 4533 3669 4723 3682
rect 4533 3617 4538 3669
rect 4590 3617 4602 3669
rect 4654 3617 4666 3669
rect 4718 3617 4723 3669
rect 4533 3604 4723 3617
rect 4533 1568 4538 3604
rect 4718 1568 4723 3604
rect 4533 1562 4723 1568
rect 5029 4119 5219 4125
rect 5029 4067 5034 4119
rect 5086 4067 5098 4119
rect 5150 4067 5162 4119
rect 5214 4067 5219 4119
rect 5029 4054 5219 4067
rect 5029 4002 5034 4054
rect 5086 4002 5098 4054
rect 5150 4002 5162 4054
rect 5214 4002 5219 4054
rect 5029 3989 5219 4002
rect 5029 3937 5034 3989
rect 5086 3937 5098 3989
rect 5150 3937 5162 3989
rect 5214 3937 5219 3989
rect 5029 3924 5219 3937
rect 5029 1568 5034 3924
rect 5214 1568 5219 3924
rect 5029 1562 5219 1568
rect 5525 4124 5715 4130
rect 5525 4072 5530 4124
rect 5582 4072 5594 4124
rect 5646 4072 5658 4124
rect 5710 4072 5715 4124
rect 5525 4059 5715 4072
rect 5525 4007 5530 4059
rect 5582 4007 5594 4059
rect 5646 4007 5658 4059
rect 5710 4007 5715 4059
rect 5525 3994 5715 4007
rect 5525 3942 5530 3994
rect 5582 3942 5594 3994
rect 5646 3942 5658 3994
rect 5710 3942 5715 3994
rect 5525 3929 5715 3942
rect 5525 3877 5530 3929
rect 5582 3877 5594 3929
rect 5646 3877 5658 3929
rect 5710 3877 5715 3929
rect 5525 3864 5715 3877
rect 5525 3812 5530 3864
rect 5582 3812 5594 3864
rect 5646 3812 5658 3864
rect 5710 3812 5715 3864
rect 5525 3799 5715 3812
rect 5525 3747 5530 3799
rect 5582 3747 5594 3799
rect 5646 3747 5658 3799
rect 5710 3747 5715 3799
rect 5525 3734 5715 3747
rect 5525 3682 5530 3734
rect 5582 3682 5594 3734
rect 5646 3682 5658 3734
rect 5710 3682 5715 3734
rect 5525 3669 5715 3682
rect 5525 3617 5530 3669
rect 5582 3617 5594 3669
rect 5646 3617 5658 3669
rect 5710 3617 5715 3669
rect 5525 3604 5715 3617
rect 5525 1568 5530 3604
rect 5710 1568 5715 3604
rect 5525 1562 5715 1568
rect 6021 4119 6211 4125
rect 6021 4067 6026 4119
rect 6078 4067 6090 4119
rect 6142 4067 6154 4119
rect 6206 4067 6211 4119
rect 6021 4054 6211 4067
rect 6021 4002 6026 4054
rect 6078 4002 6090 4054
rect 6142 4002 6154 4054
rect 6206 4002 6211 4054
rect 6021 3989 6211 4002
rect 6021 3937 6026 3989
rect 6078 3937 6090 3989
rect 6142 3937 6154 3989
rect 6206 3937 6211 3989
rect 6021 3924 6211 3937
rect 6021 1568 6026 3924
rect 6206 1568 6211 3924
rect 6021 1562 6211 1568
rect 6517 4124 6707 4130
rect 6517 4072 6522 4124
rect 6574 4072 6586 4124
rect 6638 4072 6650 4124
rect 6702 4072 6707 4124
rect 6517 4059 6707 4072
rect 6517 4007 6522 4059
rect 6574 4007 6586 4059
rect 6638 4007 6650 4059
rect 6702 4007 6707 4059
rect 6517 3994 6707 4007
rect 6517 3942 6522 3994
rect 6574 3942 6586 3994
rect 6638 3942 6650 3994
rect 6702 3942 6707 3994
rect 6517 3929 6707 3942
rect 6517 3877 6522 3929
rect 6574 3877 6586 3929
rect 6638 3877 6650 3929
rect 6702 3877 6707 3929
rect 6517 3864 6707 3877
rect 6517 3812 6522 3864
rect 6574 3812 6586 3864
rect 6638 3812 6650 3864
rect 6702 3812 6707 3864
rect 6517 3799 6707 3812
rect 6517 3747 6522 3799
rect 6574 3747 6586 3799
rect 6638 3747 6650 3799
rect 6702 3747 6707 3799
rect 6517 3734 6707 3747
rect 6517 3682 6522 3734
rect 6574 3682 6586 3734
rect 6638 3682 6650 3734
rect 6702 3682 6707 3734
rect 6517 3669 6707 3682
rect 6517 3617 6522 3669
rect 6574 3617 6586 3669
rect 6638 3617 6650 3669
rect 6702 3617 6707 3669
rect 6517 3604 6707 3617
rect 6517 1568 6522 3604
rect 6702 1568 6707 3604
rect 6517 1562 6707 1568
rect 7013 4119 7203 4125
rect 7013 4067 7018 4119
rect 7070 4067 7082 4119
rect 7134 4067 7146 4119
rect 7198 4067 7203 4119
rect 7013 4054 7203 4067
rect 7013 4002 7018 4054
rect 7070 4002 7082 4054
rect 7134 4002 7146 4054
rect 7198 4002 7203 4054
rect 7013 3989 7203 4002
rect 7013 3937 7018 3989
rect 7070 3937 7082 3989
rect 7134 3937 7146 3989
rect 7198 3937 7203 3989
rect 7013 3924 7203 3937
rect 7013 1568 7018 3924
rect 7198 1568 7203 3924
rect 7013 1562 7203 1568
rect 7509 4124 7699 4130
rect 7509 4072 7514 4124
rect 7566 4072 7578 4124
rect 7630 4072 7642 4124
rect 7694 4072 7699 4124
rect 7509 4059 7699 4072
rect 7509 4007 7514 4059
rect 7566 4007 7578 4059
rect 7630 4007 7642 4059
rect 7694 4007 7699 4059
rect 7509 3994 7699 4007
rect 7509 3942 7514 3994
rect 7566 3942 7578 3994
rect 7630 3942 7642 3994
rect 7694 3942 7699 3994
rect 7509 3929 7699 3942
rect 7509 3877 7514 3929
rect 7566 3877 7578 3929
rect 7630 3877 7642 3929
rect 7694 3877 7699 3929
rect 7509 3864 7699 3877
rect 7509 3812 7514 3864
rect 7566 3812 7578 3864
rect 7630 3812 7642 3864
rect 7694 3812 7699 3864
rect 7509 3799 7699 3812
rect 7509 3747 7514 3799
rect 7566 3747 7578 3799
rect 7630 3747 7642 3799
rect 7694 3747 7699 3799
rect 7509 3734 7699 3747
rect 7509 3682 7514 3734
rect 7566 3682 7578 3734
rect 7630 3682 7642 3734
rect 7694 3682 7699 3734
rect 7509 3669 7699 3682
rect 7509 3617 7514 3669
rect 7566 3617 7578 3669
rect 7630 3617 7642 3669
rect 7694 3617 7699 3669
rect 7509 3604 7699 3617
rect 7509 1568 7514 3604
rect 7694 1568 7699 3604
rect 7509 1562 7699 1568
rect 8005 4119 8195 4125
rect 8005 4067 8010 4119
rect 8062 4067 8074 4119
rect 8126 4067 8138 4119
rect 8190 4067 8195 4119
rect 8005 4054 8195 4067
rect 8005 4002 8010 4054
rect 8062 4002 8074 4054
rect 8126 4002 8138 4054
rect 8190 4002 8195 4054
rect 8005 3989 8195 4002
rect 8005 3937 8010 3989
rect 8062 3937 8074 3989
rect 8126 3937 8138 3989
rect 8190 3937 8195 3989
rect 8005 3924 8195 3937
rect 8005 1568 8010 3924
rect 8190 1568 8195 3924
rect 8005 1562 8195 1568
rect 8501 4124 8691 4130
rect 8501 4072 8506 4124
rect 8558 4072 8570 4124
rect 8622 4072 8634 4124
rect 8686 4072 8691 4124
rect 8501 4059 8691 4072
rect 8501 4007 8506 4059
rect 8558 4007 8570 4059
rect 8622 4007 8634 4059
rect 8686 4007 8691 4059
rect 8501 3994 8691 4007
rect 8501 3942 8506 3994
rect 8558 3942 8570 3994
rect 8622 3942 8634 3994
rect 8686 3942 8691 3994
rect 8501 3929 8691 3942
rect 8501 3877 8506 3929
rect 8558 3877 8570 3929
rect 8622 3877 8634 3929
rect 8686 3877 8691 3929
rect 8501 3864 8691 3877
rect 8501 3812 8506 3864
rect 8558 3812 8570 3864
rect 8622 3812 8634 3864
rect 8686 3812 8691 3864
rect 8501 3799 8691 3812
rect 8501 3747 8506 3799
rect 8558 3747 8570 3799
rect 8622 3747 8634 3799
rect 8686 3747 8691 3799
rect 8501 3734 8691 3747
rect 8501 3682 8506 3734
rect 8558 3682 8570 3734
rect 8622 3682 8634 3734
rect 8686 3682 8691 3734
rect 8501 3669 8691 3682
rect 8501 3617 8506 3669
rect 8558 3617 8570 3669
rect 8622 3617 8634 3669
rect 8686 3617 8691 3669
rect 8501 3604 8691 3617
rect 8501 1568 8506 3604
rect 8686 1568 8691 3604
rect 8501 1562 8691 1568
rect 8997 4119 9187 4125
rect 8997 4067 9002 4119
rect 9054 4067 9066 4119
rect 9118 4067 9130 4119
rect 9182 4067 9187 4119
rect 8997 4054 9187 4067
rect 8997 4002 9002 4054
rect 9054 4002 9066 4054
rect 9118 4002 9130 4054
rect 9182 4002 9187 4054
rect 8997 3989 9187 4002
rect 8997 3937 9002 3989
rect 9054 3937 9066 3989
rect 9118 3937 9130 3989
rect 9182 3937 9187 3989
rect 8997 3924 9187 3937
rect 8997 1568 9002 3924
rect 9182 1568 9187 3924
rect 8997 1562 9187 1568
rect 9493 4124 9683 4130
rect 9493 4072 9498 4124
rect 9550 4072 9562 4124
rect 9614 4072 9626 4124
rect 9678 4072 9683 4124
rect 9493 4059 9683 4072
rect 9493 4007 9498 4059
rect 9550 4007 9562 4059
rect 9614 4007 9626 4059
rect 9678 4007 9683 4059
rect 9493 3994 9683 4007
rect 9493 3942 9498 3994
rect 9550 3942 9562 3994
rect 9614 3942 9626 3994
rect 9678 3942 9683 3994
rect 9493 3929 9683 3942
rect 9493 3877 9498 3929
rect 9550 3877 9562 3929
rect 9614 3877 9626 3929
rect 9678 3877 9683 3929
rect 9493 3864 9683 3877
rect 9493 3812 9498 3864
rect 9550 3812 9562 3864
rect 9614 3812 9626 3864
rect 9678 3812 9683 3864
rect 9493 3799 9683 3812
rect 9493 3747 9498 3799
rect 9550 3747 9562 3799
rect 9614 3747 9626 3799
rect 9678 3747 9683 3799
rect 9493 3734 9683 3747
rect 9493 3682 9498 3734
rect 9550 3682 9562 3734
rect 9614 3682 9626 3734
rect 9678 3682 9683 3734
rect 9493 3669 9683 3682
rect 9493 3617 9498 3669
rect 9550 3617 9562 3669
rect 9614 3617 9626 3669
rect 9678 3617 9683 3669
rect 9493 3604 9683 3617
rect 9493 1568 9498 3604
rect 9678 1568 9683 3604
rect 9493 1562 9683 1568
rect 9989 4119 10179 4125
rect 9989 4067 9994 4119
rect 10046 4067 10058 4119
rect 10110 4067 10122 4119
rect 10174 4067 10179 4119
rect 9989 4054 10179 4067
rect 9989 4002 9994 4054
rect 10046 4002 10058 4054
rect 10110 4002 10122 4054
rect 10174 4002 10179 4054
rect 9989 3989 10179 4002
rect 9989 3937 9994 3989
rect 10046 3937 10058 3989
rect 10110 3937 10122 3989
rect 10174 3937 10179 3989
rect 9989 3924 10179 3937
rect 9989 1568 9994 3924
rect 10174 1568 10179 3924
rect 9989 1562 10179 1568
rect 10485 4124 10675 4130
rect 10485 4072 10490 4124
rect 10542 4072 10554 4124
rect 10606 4072 10618 4124
rect 10670 4072 10675 4124
rect 10485 4059 10675 4072
rect 10485 4007 10490 4059
rect 10542 4007 10554 4059
rect 10606 4007 10618 4059
rect 10670 4007 10675 4059
rect 10485 3994 10675 4007
rect 10485 3942 10490 3994
rect 10542 3942 10554 3994
rect 10606 3942 10618 3994
rect 10670 3942 10675 3994
rect 10485 3929 10675 3942
rect 10485 3877 10490 3929
rect 10542 3877 10554 3929
rect 10606 3877 10618 3929
rect 10670 3877 10675 3929
rect 10485 3864 10675 3877
rect 10485 3812 10490 3864
rect 10542 3812 10554 3864
rect 10606 3812 10618 3864
rect 10670 3812 10675 3864
rect 10485 3799 10675 3812
rect 10485 3747 10490 3799
rect 10542 3747 10554 3799
rect 10606 3747 10618 3799
rect 10670 3747 10675 3799
rect 10485 3734 10675 3747
rect 10485 3682 10490 3734
rect 10542 3682 10554 3734
rect 10606 3682 10618 3734
rect 10670 3682 10675 3734
rect 10485 3669 10675 3682
rect 10485 3617 10490 3669
rect 10542 3617 10554 3669
rect 10606 3617 10618 3669
rect 10670 3617 10675 3669
rect 10485 3604 10675 3617
rect 10485 1568 10490 3604
rect 10670 1568 10675 3604
rect 10485 1562 10675 1568
rect 10981 4119 11171 4125
rect 10981 4067 10986 4119
rect 11038 4067 11050 4119
rect 11102 4067 11114 4119
rect 11166 4067 11171 4119
rect 10981 4054 11171 4067
rect 10981 4002 10986 4054
rect 11038 4002 11050 4054
rect 11102 4002 11114 4054
rect 11166 4002 11171 4054
rect 10981 3989 11171 4002
rect 10981 3937 10986 3989
rect 11038 3937 11050 3989
rect 11102 3937 11114 3989
rect 11166 3937 11171 3989
rect 10981 3924 11171 3937
rect 10981 1568 10986 3924
rect 11166 1568 11171 3924
rect 10981 1562 11171 1568
rect 11477 4124 11667 4130
rect 11477 4072 11482 4124
rect 11534 4072 11546 4124
rect 11598 4072 11610 4124
rect 11662 4072 11667 4124
rect 11477 4059 11667 4072
rect 11477 4007 11482 4059
rect 11534 4007 11546 4059
rect 11598 4007 11610 4059
rect 11662 4007 11667 4059
rect 11477 3994 11667 4007
rect 11477 3942 11482 3994
rect 11534 3942 11546 3994
rect 11598 3942 11610 3994
rect 11662 3942 11667 3994
rect 11477 3929 11667 3942
rect 11477 3877 11482 3929
rect 11534 3877 11546 3929
rect 11598 3877 11610 3929
rect 11662 3877 11667 3929
rect 11477 3864 11667 3877
rect 11477 3812 11482 3864
rect 11534 3812 11546 3864
rect 11598 3812 11610 3864
rect 11662 3812 11667 3864
rect 11477 3799 11667 3812
rect 11477 3747 11482 3799
rect 11534 3747 11546 3799
rect 11598 3747 11610 3799
rect 11662 3747 11667 3799
rect 11477 3734 11667 3747
rect 11477 3682 11482 3734
rect 11534 3682 11546 3734
rect 11598 3682 11610 3734
rect 11662 3682 11667 3734
rect 11477 3669 11667 3682
rect 11477 3617 11482 3669
rect 11534 3617 11546 3669
rect 11598 3617 11610 3669
rect 11662 3617 11667 3669
rect 11477 3604 11667 3617
rect 11477 1568 11482 3604
rect 11662 1568 11667 3604
rect 11477 1562 11667 1568
rect 11973 4119 12163 4125
rect 11973 4067 11978 4119
rect 12030 4067 12042 4119
rect 12094 4067 12106 4119
rect 12158 4067 12163 4119
rect 11973 4054 12163 4067
rect 11973 4002 11978 4054
rect 12030 4002 12042 4054
rect 12094 4002 12106 4054
rect 12158 4002 12163 4054
rect 11973 3989 12163 4002
rect 11973 3937 11978 3989
rect 12030 3937 12042 3989
rect 12094 3937 12106 3989
rect 12158 3937 12163 3989
rect 11973 3924 12163 3937
rect 11973 1568 11978 3924
rect 12158 1568 12163 3924
rect 11973 1562 12163 1568
rect 12469 4124 12659 4130
rect 12469 4072 12474 4124
rect 12526 4072 12538 4124
rect 12590 4072 12602 4124
rect 12654 4072 12659 4124
rect 12469 4059 12659 4072
rect 12469 4007 12474 4059
rect 12526 4007 12538 4059
rect 12590 4007 12602 4059
rect 12654 4007 12659 4059
rect 12469 3994 12659 4007
rect 12469 3942 12474 3994
rect 12526 3942 12538 3994
rect 12590 3942 12602 3994
rect 12654 3942 12659 3994
rect 12469 3929 12659 3942
rect 12469 3877 12474 3929
rect 12526 3877 12538 3929
rect 12590 3877 12602 3929
rect 12654 3877 12659 3929
rect 12469 3864 12659 3877
rect 12469 3812 12474 3864
rect 12526 3812 12538 3864
rect 12590 3812 12602 3864
rect 12654 3812 12659 3864
rect 12469 3799 12659 3812
rect 12469 3747 12474 3799
rect 12526 3747 12538 3799
rect 12590 3747 12602 3799
rect 12654 3747 12659 3799
rect 12469 3734 12659 3747
rect 12469 3682 12474 3734
rect 12526 3682 12538 3734
rect 12590 3682 12602 3734
rect 12654 3682 12659 3734
rect 12469 3669 12659 3682
rect 12469 3617 12474 3669
rect 12526 3617 12538 3669
rect 12590 3617 12602 3669
rect 12654 3617 12659 3669
rect 12469 3604 12659 3617
rect 12469 1568 12474 3604
rect 12654 1568 12659 3604
rect 12469 1562 12659 1568
rect 12965 4119 13155 4125
rect 12965 4067 12970 4119
rect 13022 4067 13034 4119
rect 13086 4067 13098 4119
rect 13150 4067 13155 4119
rect 12965 4054 13155 4067
rect 12965 4002 12970 4054
rect 13022 4002 13034 4054
rect 13086 4002 13098 4054
rect 13150 4002 13155 4054
rect 12965 3989 13155 4002
rect 12965 3937 12970 3989
rect 13022 3937 13034 3989
rect 13086 3937 13098 3989
rect 13150 3937 13155 3989
rect 12965 3924 13155 3937
rect 12965 1568 12970 3924
rect 13150 1568 13155 3924
rect 12965 1562 13155 1568
rect 13461 4124 13651 4130
rect 13461 4072 13466 4124
rect 13518 4072 13530 4124
rect 13582 4072 13594 4124
rect 13646 4072 13651 4124
rect 13461 4059 13651 4072
rect 13461 4007 13466 4059
rect 13518 4007 13530 4059
rect 13582 4007 13594 4059
rect 13646 4007 13651 4059
rect 13461 3994 13651 4007
rect 13461 3942 13466 3994
rect 13518 3942 13530 3994
rect 13582 3942 13594 3994
rect 13646 3942 13651 3994
rect 13461 3929 13651 3942
rect 13461 3877 13466 3929
rect 13518 3877 13530 3929
rect 13582 3877 13594 3929
rect 13646 3877 13651 3929
rect 13461 3864 13651 3877
rect 13461 3812 13466 3864
rect 13518 3812 13530 3864
rect 13582 3812 13594 3864
rect 13646 3812 13651 3864
rect 13461 3799 13651 3812
rect 13461 3747 13466 3799
rect 13518 3747 13530 3799
rect 13582 3747 13594 3799
rect 13646 3747 13651 3799
rect 13461 3734 13651 3747
rect 13461 3682 13466 3734
rect 13518 3682 13530 3734
rect 13582 3682 13594 3734
rect 13646 3682 13651 3734
rect 13461 3669 13651 3682
rect 13461 3617 13466 3669
rect 13518 3617 13530 3669
rect 13582 3617 13594 3669
rect 13646 3617 13651 3669
rect 13461 3604 13651 3617
rect 13461 1568 13466 3604
rect 13646 1568 13651 3604
rect 13461 1562 13651 1568
rect 13991 4124 14135 4130
rect 14043 4072 14083 4124
rect 13991 4060 14135 4072
rect 14043 4008 14083 4060
rect 13991 3996 14135 4008
rect 14043 3944 14083 3996
rect 13991 3932 14135 3944
rect 14043 3880 14083 3932
rect 13991 3868 14135 3880
rect 14043 3816 14083 3868
rect 13991 3804 14135 3816
rect 14043 3752 14083 3804
rect 13991 3740 14135 3752
rect 14043 3688 14083 3740
rect 13991 3676 14135 3688
rect 14043 3624 14083 3676
rect 13991 3612 14135 3624
rect 14043 3560 14083 3612
rect 13991 3548 14135 3560
rect 14043 3496 14083 3548
rect 13991 3484 14135 3496
rect 14043 3432 14083 3484
rect 13991 3420 14135 3432
rect 14043 3368 14083 3420
rect 13991 3356 14135 3368
rect 14043 3304 14083 3356
rect 13991 3292 14135 3304
rect 14043 3240 14083 3292
rect 13991 3228 14135 3240
rect 14043 3176 14083 3228
rect 13991 3164 14135 3176
rect 14043 3112 14083 3164
rect 13991 3100 14135 3112
rect 14043 3048 14083 3100
rect 13991 3036 14135 3048
rect 14043 2984 14083 3036
rect 13991 2972 14135 2984
rect 14043 2920 14083 2972
rect 13991 2908 14135 2920
rect 14043 2856 14083 2908
rect 13991 2844 14135 2856
rect 14043 2792 14083 2844
rect 13991 2780 14135 2792
rect 14043 2728 14083 2780
rect 13991 2716 14135 2728
rect 14043 2664 14083 2716
rect 13991 2652 14135 2664
rect 14043 2600 14083 2652
rect 13991 2588 14135 2600
rect 14043 2536 14083 2588
rect 13991 2524 14135 2536
rect 14043 2472 14083 2524
rect 13991 2460 14135 2472
rect 14043 2408 14083 2460
rect 13991 2396 14135 2408
rect 14043 2344 14083 2396
rect 13991 2332 14135 2344
rect 14043 2280 14083 2332
rect 13991 2268 14135 2280
rect 14043 2216 14083 2268
rect 13991 2204 14135 2216
rect 14043 2152 14083 2204
rect 13991 2140 14135 2152
rect 14043 2088 14083 2140
rect 13991 2075 14135 2088
rect 14043 2023 14083 2075
rect 13991 2010 14135 2023
rect 14043 1958 14083 2010
rect 13991 1945 14135 1958
rect 14043 1893 14083 1945
rect 13991 1880 14135 1893
rect 14043 1828 14083 1880
rect 13991 1815 14135 1828
rect 14043 1763 14083 1815
rect 13991 1750 14135 1763
rect 14043 1698 14083 1750
rect 13991 1685 14135 1698
rect 14043 1633 14083 1685
rect 13991 1620 14135 1633
rect 14043 1568 14083 1620
rect 13991 1562 14135 1568
rect 14350 4124 14618 4130
rect 14402 4072 14422 4124
rect 14474 4072 14494 4124
rect 14546 4072 14566 4124
rect 14350 4059 14618 4072
rect 14402 4007 14422 4059
rect 14474 4007 14494 4059
rect 14546 4007 14566 4059
rect 14350 3994 14618 4007
rect 14402 3942 14422 3994
rect 14474 3942 14494 3994
rect 14546 3942 14566 3994
rect 14350 3929 14618 3942
rect 14402 3877 14422 3929
rect 14474 3877 14494 3929
rect 14546 3877 14566 3929
rect 14350 3864 14618 3877
rect 14402 3812 14422 3864
rect 14474 3812 14494 3864
rect 14546 3812 14566 3864
rect 14350 3799 14618 3812
rect 14402 3747 14422 3799
rect 14474 3747 14494 3799
rect 14546 3747 14566 3799
rect 14350 3734 14618 3747
rect 14402 3682 14422 3734
rect 14474 3682 14494 3734
rect 14546 3682 14566 3734
rect 14350 3669 14618 3682
rect 14402 3617 14422 3669
rect 14474 3617 14494 3669
rect 14546 3617 14566 3669
rect 14350 3604 14618 3617
rect 14402 3552 14422 3604
rect 14474 3552 14494 3604
rect 14546 3552 14566 3604
rect 14350 3540 14618 3552
rect 14402 3488 14422 3540
rect 14474 3488 14494 3540
rect 14546 3488 14566 3540
rect 14350 3476 14618 3488
rect 14402 3424 14422 3476
rect 14474 3424 14494 3476
rect 14546 3424 14566 3476
rect 14350 3412 14618 3424
rect 14402 3360 14422 3412
rect 14474 3360 14494 3412
rect 14546 3360 14566 3412
rect 14350 3348 14618 3360
rect 14402 3296 14422 3348
rect 14474 3296 14494 3348
rect 14546 3296 14566 3348
rect 14350 3284 14618 3296
rect 14402 3232 14422 3284
rect 14474 3232 14494 3284
rect 14546 3232 14566 3284
rect 14350 3220 14618 3232
rect 14402 3168 14422 3220
rect 14474 3168 14494 3220
rect 14546 3168 14566 3220
rect 14350 3156 14618 3168
rect 14402 3104 14422 3156
rect 14474 3104 14494 3156
rect 14546 3104 14566 3156
rect 14350 3092 14618 3104
rect 14402 3040 14422 3092
rect 14474 3040 14494 3092
rect 14546 3040 14566 3092
rect 14350 3028 14618 3040
rect 14402 2976 14422 3028
rect 14474 2976 14494 3028
rect 14546 2976 14566 3028
rect 14350 2964 14618 2976
rect 14402 2912 14422 2964
rect 14474 2912 14494 2964
rect 14546 2912 14566 2964
rect 14350 2900 14618 2912
rect 14402 2848 14422 2900
rect 14474 2848 14494 2900
rect 14546 2848 14566 2900
rect 14350 2836 14618 2848
rect 14402 2784 14422 2836
rect 14474 2784 14494 2836
rect 14546 2784 14566 2836
rect 14350 2772 14618 2784
rect 14402 2720 14422 2772
rect 14474 2720 14494 2772
rect 14546 2720 14566 2772
rect 14350 2708 14618 2720
rect 14402 2656 14422 2708
rect 14474 2656 14494 2708
rect 14546 2656 14566 2708
rect 14350 2644 14618 2656
rect 14402 2592 14422 2644
rect 14474 2592 14494 2644
rect 14546 2592 14566 2644
rect 14350 2580 14618 2592
rect 14402 2528 14422 2580
rect 14474 2528 14494 2580
rect 14546 2528 14566 2580
rect 14350 2516 14618 2528
rect 14402 2464 14422 2516
rect 14474 2464 14494 2516
rect 14546 2464 14566 2516
rect 14350 2452 14618 2464
rect 14402 2400 14422 2452
rect 14474 2400 14494 2452
rect 14546 2400 14566 2452
rect 14350 2388 14618 2400
rect 14402 2336 14422 2388
rect 14474 2336 14494 2388
rect 14546 2336 14566 2388
rect 14350 2324 14618 2336
rect 14402 2272 14422 2324
rect 14474 2272 14494 2324
rect 14546 2272 14566 2324
rect 14350 2260 14618 2272
rect 14402 2208 14422 2260
rect 14474 2208 14494 2260
rect 14546 2208 14566 2260
rect 14350 2196 14618 2208
rect 14402 2144 14422 2196
rect 14474 2144 14494 2196
rect 14546 2144 14566 2196
rect 14350 2132 14618 2144
rect 14402 2080 14422 2132
rect 14474 2080 14494 2132
rect 14546 2080 14566 2132
rect 14350 2068 14618 2080
rect 14402 2016 14422 2068
rect 14474 2016 14494 2068
rect 14546 2016 14566 2068
rect 14350 2004 14618 2016
rect 14402 1952 14422 2004
rect 14474 1952 14494 2004
rect 14546 1952 14566 2004
rect 14350 1940 14618 1952
rect 14402 1888 14422 1940
rect 14474 1888 14494 1940
rect 14546 1888 14566 1940
rect 14350 1876 14618 1888
rect 14402 1824 14422 1876
rect 14474 1824 14494 1876
rect 14546 1824 14566 1876
rect 14350 1812 14618 1824
rect 14402 1760 14422 1812
rect 14474 1760 14494 1812
rect 14546 1760 14566 1812
rect 14350 1748 14618 1760
rect 14402 1696 14422 1748
rect 14474 1696 14494 1748
rect 14546 1696 14566 1748
rect 14350 1684 14618 1696
rect 14402 1632 14422 1684
rect 14474 1632 14494 1684
rect 14546 1632 14566 1684
rect 14350 1620 14618 1632
rect 14402 1568 14422 1620
rect 14474 1568 14494 1620
rect 14546 1568 14566 1620
rect 14350 1562 14618 1568
rect 518 1530 786 1543
rect 570 1478 590 1530
rect 642 1478 662 1530
rect 714 1478 734 1530
rect 518 1465 786 1478
rect 570 1413 590 1465
rect 642 1413 662 1465
rect 714 1413 734 1465
rect 518 1400 786 1413
rect 570 1348 590 1400
rect 642 1348 662 1400
rect 714 1348 734 1400
rect 518 1335 786 1348
rect 570 1283 590 1335
rect 642 1283 662 1335
rect 714 1283 734 1335
rect 518 1270 786 1283
rect 570 1218 590 1270
rect 642 1218 662 1270
rect 714 1218 734 1270
rect 518 1205 786 1218
rect 570 1153 590 1205
rect 642 1153 662 1205
rect 714 1153 734 1205
rect 518 1140 786 1153
rect 570 1088 590 1140
rect 642 1088 662 1140
rect 714 1088 734 1140
rect 518 1075 786 1088
rect 570 1023 590 1075
rect 642 1023 662 1075
rect 714 1023 734 1075
rect 518 1010 786 1023
rect 570 958 590 1010
rect 642 958 662 1010
rect 714 958 734 1010
rect 518 945 786 958
rect 570 893 590 945
rect 642 893 662 945
rect 714 893 734 945
rect 518 880 786 893
rect 570 828 590 880
rect 642 828 662 880
rect 714 828 734 880
rect 518 822 786 828
use sky130_fd_pr__via_l1m1_centered__example_559591418086  sky130_fd_pr__via_l1m1_centered__example_559591418086_0
timestamp 1624884095
transform 1 0 941 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_0
timestamp 1624884095
transform 1 0 1371 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_1
timestamp 1624884095
transform 1 0 7885 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_2
timestamp 1624884095
transform 1 0 6893 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_3
timestamp 1624884095
transform 1 0 5901 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_4
timestamp 1624884095
transform 1 0 4909 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_5
timestamp 1624884095
transform 1 0 3917 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_6
timestamp 1624884095
transform 1 0 2925 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_7
timestamp 1624884095
transform 1 0 1933 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_8
timestamp 1624884095
transform 1 0 10861 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_9
timestamp 1624884095
transform 1 0 9869 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_10
timestamp 1624884095
transform 1 0 8877 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_11
timestamp 1624884095
transform 1 0 11291 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_12
timestamp 1624884095
transform 1 0 10299 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_13
timestamp 1624884095
transform 1 0 9307 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_14
timestamp 1624884095
transform 1 0 2363 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_15
timestamp 1624884095
transform 1 0 3355 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_16
timestamp 1624884095
transform 1 0 4347 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_17
timestamp 1624884095
transform 1 0 5339 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_18
timestamp 1624884095
transform 1 0 6331 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_19
timestamp 1624884095
transform 1 0 7323 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_20
timestamp 1624884095
transform 1 0 8315 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_21
timestamp 1624884095
transform 1 0 11853 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_22
timestamp 1624884095
transform 1 0 12283 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_23
timestamp 1624884095
transform 1 0 13275 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_24
timestamp 1624884095
transform 1 0 12845 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_25
timestamp 1624884095
transform 1 0 13837 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_26
timestamp 1624884095
transform 1 0 14195 0 1 1197
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_5595914180812  sky130_fd_pr__via_l1m1_centered__example_5595914180812_0
timestamp 1624884095
transform -1 0 142 0 1 348
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_5595914180811  sky130_fd_pr__via_l1m1_centered__example_5595914180811_0
timestamp 1624884095
transform -1 0 14924 0 1 437
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_0
timestamp 1624884095
transform -1 0 8164 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_1
timestamp 1624884095
transform 1 0 8036 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_2
timestamp 1624884095
transform -1 0 7172 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_3
timestamp 1624884095
transform -1 0 6180 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_4
timestamp 1624884095
transform -1 0 5188 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_5
timestamp 1624884095
transform -1 0 4196 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_6
timestamp 1624884095
transform -1 0 3204 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_7
timestamp 1624884095
transform -1 0 2212 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_8
timestamp 1624884095
transform 1 0 7044 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_9
timestamp 1624884095
transform -1 0 1220 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_10
timestamp 1624884095
transform 1 0 6052 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_11
timestamp 1624884095
transform 1 0 5060 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_12
timestamp 1624884095
transform 1 0 1092 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_13
timestamp 1624884095
transform 1 0 2084 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_14
timestamp 1624884095
transform 1 0 3076 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_15
timestamp 1624884095
transform 1 0 4068 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_16
timestamp 1624884095
transform 1 0 9028 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_17
timestamp 1624884095
transform 1 0 10020 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_18
timestamp 1624884095
transform 1 0 11012 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_19
timestamp 1624884095
transform 1 0 12004 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_20
timestamp 1624884095
transform -1 0 9156 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_21
timestamp 1624884095
transform -1 0 10148 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_22
timestamp 1624884095
transform -1 0 11140 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_23
timestamp 1624884095
transform -1 0 12132 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_24
timestamp 1624884095
transform 1 0 12996 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_25
timestamp 1624884095
transform -1 0 13124 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_26
timestamp 1624884095
transform -1 0 13124 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_27
timestamp 1624884095
transform 1 0 12996 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_28
timestamp 1624884095
transform -1 0 12132 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_29
timestamp 1624884095
transform -1 0 11140 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_30
timestamp 1624884095
transform -1 0 10148 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_31
timestamp 1624884095
transform -1 0 9156 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_32
timestamp 1624884095
transform 1 0 12004 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_33
timestamp 1624884095
transform 1 0 11012 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_34
timestamp 1624884095
transform 1 0 10020 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_35
timestamp 1624884095
transform 1 0 9028 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_36
timestamp 1624884095
transform 1 0 4068 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_37
timestamp 1624884095
transform 1 0 3076 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_38
timestamp 1624884095
transform 1 0 2084 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_39
timestamp 1624884095
transform 1 0 1092 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_40
timestamp 1624884095
transform 1 0 5060 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_41
timestamp 1624884095
transform 1 0 6052 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_42
timestamp 1624884095
transform -1 0 1220 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_43
timestamp 1624884095
transform 1 0 7044 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_44
timestamp 1624884095
transform -1 0 2212 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_45
timestamp 1624884095
transform -1 0 3204 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_46
timestamp 1624884095
transform -1 0 4196 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_47
timestamp 1624884095
transform -1 0 5188 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_48
timestamp 1624884095
transform -1 0 6180 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_49
timestamp 1624884095
transform -1 0 7172 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_50
timestamp 1624884095
transform 1 0 8036 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_51
timestamp 1624884095
transform -1 0 8164 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_52
timestamp 1624884095
transform 1 0 734 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_53
timestamp 1624884095
transform -1 0 14401 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_54
timestamp 1624884095
transform 1 0 13988 0 1 1552
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_55
timestamp 1624884095
transform 1 0 13988 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_56
timestamp 1624884095
transform -1 0 14401 0 1 3152
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_57
timestamp 1624884095
transform 1 0 734 0 1 3152
box 0 0 1 1
use sky130_fd_pr__pfet_01v8__example_55959141808658  sky130_fd_pr__pfet_01v8__example_55959141808658_0
timestamp 1624884095
transform 1 0 881 0 -1 2552
box -25 0 13041 500
use sky130_fd_pr__pfet_01v8__example_55959141808658  sky130_fd_pr__pfet_01v8__example_55959141808658_1
timestamp 1624884095
transform 1 0 881 0 1 3152
box -25 0 13041 500
use sky130_fd_pr__pfet_01v8__example_55959141808657  sky130_fd_pr__pfet_01v8__example_55959141808657_0
timestamp 1624884095
transform 1 0 14135 0 1 1552
box -25 500 145 501
use sky130_fd_pr__pfet_01v8__example_55959141808657  sky130_fd_pr__pfet_01v8__example_55959141808657_1
timestamp 1624884095
transform 1 0 14135 0 1 3152
box -25 500 145 501
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 976038
string GDS_START 186236
<< end >>
