magic
tech sky130A
magscale 1 2
timestamp 1624883981
<< checkpaint >>
rect -1246 -1260 2128 1968
<< pwell >>
rect 15 163 867 545
<< nmos >>
rect 171 189 201 519
rect 257 189 307 519
rect 363 189 413 519
rect 469 189 519 519
rect 575 189 625 519
rect 681 189 711 519
<< ndiff >>
rect 111 507 171 519
rect 111 473 126 507
rect 160 473 171 507
rect 111 439 171 473
rect 111 405 126 439
rect 160 405 171 439
rect 111 371 171 405
rect 111 337 126 371
rect 160 337 171 371
rect 111 303 171 337
rect 111 269 126 303
rect 160 269 171 303
rect 111 235 171 269
rect 111 201 126 235
rect 160 201 171 235
rect 111 189 171 201
rect 201 507 257 519
rect 201 473 212 507
rect 246 473 257 507
rect 201 439 257 473
rect 201 405 212 439
rect 246 405 257 439
rect 201 371 257 405
rect 201 337 212 371
rect 246 337 257 371
rect 201 303 257 337
rect 201 269 212 303
rect 246 269 257 303
rect 201 235 257 269
rect 201 201 212 235
rect 246 201 257 235
rect 201 189 257 201
rect 307 507 363 519
rect 307 473 318 507
rect 352 473 363 507
rect 307 439 363 473
rect 307 405 318 439
rect 352 405 363 439
rect 307 371 363 405
rect 307 337 318 371
rect 352 337 363 371
rect 307 303 363 337
rect 307 269 318 303
rect 352 269 363 303
rect 307 235 363 269
rect 307 201 318 235
rect 352 201 363 235
rect 307 189 363 201
rect 413 507 469 519
rect 413 473 424 507
rect 458 473 469 507
rect 413 439 469 473
rect 413 405 424 439
rect 458 405 469 439
rect 413 371 469 405
rect 413 337 424 371
rect 458 337 469 371
rect 413 303 469 337
rect 413 269 424 303
rect 458 269 469 303
rect 413 235 469 269
rect 413 201 424 235
rect 458 201 469 235
rect 413 189 469 201
rect 519 507 575 519
rect 519 473 530 507
rect 564 473 575 507
rect 519 439 575 473
rect 519 405 530 439
rect 564 405 575 439
rect 519 371 575 405
rect 519 337 530 371
rect 564 337 575 371
rect 519 303 575 337
rect 519 269 530 303
rect 564 269 575 303
rect 519 235 575 269
rect 519 201 530 235
rect 564 201 575 235
rect 519 189 575 201
rect 625 507 681 519
rect 625 473 636 507
rect 670 473 681 507
rect 625 439 681 473
rect 625 405 636 439
rect 670 405 681 439
rect 625 371 681 405
rect 625 337 636 371
rect 670 337 681 371
rect 625 303 681 337
rect 625 269 636 303
rect 670 269 681 303
rect 625 235 681 269
rect 625 201 636 235
rect 670 201 681 235
rect 625 189 681 201
rect 711 507 771 519
rect 711 473 722 507
rect 756 473 771 507
rect 711 439 771 473
rect 711 405 722 439
rect 756 405 771 439
rect 711 371 771 405
rect 711 337 722 371
rect 756 337 771 371
rect 711 303 771 337
rect 711 269 722 303
rect 756 269 771 303
rect 711 235 771 269
rect 711 201 722 235
rect 756 201 771 235
rect 711 189 771 201
<< ndiffc >>
rect 126 473 160 507
rect 126 405 160 439
rect 126 337 160 371
rect 126 269 160 303
rect 126 201 160 235
rect 212 473 246 507
rect 212 405 246 439
rect 212 337 246 371
rect 212 269 246 303
rect 212 201 246 235
rect 318 473 352 507
rect 318 405 352 439
rect 318 337 352 371
rect 318 269 352 303
rect 318 201 352 235
rect 424 473 458 507
rect 424 405 458 439
rect 424 337 458 371
rect 424 269 458 303
rect 424 201 458 235
rect 530 473 564 507
rect 530 405 564 439
rect 530 337 564 371
rect 530 269 564 303
rect 530 201 564 235
rect 636 473 670 507
rect 636 405 670 439
rect 636 337 670 371
rect 636 269 670 303
rect 636 201 670 235
rect 722 473 756 507
rect 722 405 756 439
rect 722 337 756 371
rect 722 269 756 303
rect 722 201 756 235
<< psubdiff >>
rect 41 507 111 519
rect 41 473 58 507
rect 92 473 111 507
rect 41 439 111 473
rect 41 405 58 439
rect 92 405 111 439
rect 41 371 111 405
rect 41 337 58 371
rect 92 337 111 371
rect 41 303 111 337
rect 41 269 58 303
rect 92 269 111 303
rect 41 235 111 269
rect 41 201 58 235
rect 92 201 111 235
rect 41 189 111 201
rect 771 507 841 519
rect 771 473 790 507
rect 824 473 841 507
rect 771 439 841 473
rect 771 405 790 439
rect 824 405 841 439
rect 771 371 841 405
rect 771 337 790 371
rect 824 337 841 371
rect 771 303 841 337
rect 771 269 790 303
rect 824 269 841 303
rect 771 235 841 269
rect 771 201 790 235
rect 824 201 841 235
rect 771 189 841 201
<< psubdiffcont >>
rect 58 473 92 507
rect 58 405 92 439
rect 58 337 92 371
rect 58 269 92 303
rect 58 201 92 235
rect 790 473 824 507
rect 790 405 824 439
rect 790 337 824 371
rect 790 269 824 303
rect 790 201 824 235
<< poly >>
rect 243 687 639 708
rect 120 595 201 611
rect 120 561 136 595
rect 170 561 201 595
rect 243 585 288 687
rect 594 585 639 687
rect 243 569 639 585
rect 681 595 762 611
rect 120 545 201 561
rect 171 519 201 545
rect 257 519 307 569
rect 363 519 413 569
rect 469 519 519 569
rect 575 519 625 569
rect 681 561 712 595
rect 746 561 762 595
rect 681 545 762 561
rect 681 519 711 545
rect 171 163 201 189
rect 120 147 201 163
rect 120 113 136 147
rect 170 113 201 147
rect 257 139 307 189
rect 363 139 413 189
rect 469 139 519 189
rect 575 139 625 189
rect 681 163 711 189
rect 681 147 762 163
rect 120 97 201 113
rect 243 123 639 139
rect 243 21 288 123
rect 594 21 639 123
rect 681 113 712 147
rect 746 113 762 147
rect 681 97 762 113
rect 243 0 639 21
<< polycont >>
rect 136 561 170 595
rect 288 585 594 687
rect 712 561 746 595
rect 136 113 170 147
rect 288 21 594 123
rect 712 113 746 147
<< locali >>
rect 266 689 616 708
rect 120 595 186 611
rect 120 561 136 595
rect 170 561 186 595
rect 266 583 280 689
rect 602 583 616 689
rect 266 569 616 583
rect 696 595 762 611
rect 120 545 186 561
rect 696 561 712 595
rect 746 561 762 595
rect 696 545 762 561
rect 120 523 160 545
rect 722 523 762 545
rect 41 507 160 523
rect 41 473 58 507
rect 92 479 126 507
rect 94 473 126 479
rect 41 445 60 473
rect 94 445 160 473
rect 41 439 160 445
rect 41 405 58 439
rect 92 407 126 439
rect 94 405 126 407
rect 41 373 60 405
rect 94 373 160 405
rect 41 371 160 373
rect 41 337 58 371
rect 92 337 126 371
rect 41 335 160 337
rect 41 303 60 335
rect 94 303 160 335
rect 41 269 58 303
rect 94 301 126 303
rect 92 269 126 301
rect 41 263 160 269
rect 41 235 60 263
rect 94 235 160 263
rect 41 201 58 235
rect 94 229 126 235
rect 92 201 126 229
rect 41 185 160 201
rect 212 507 246 523
rect 212 439 246 445
rect 212 371 246 373
rect 212 335 246 337
rect 212 263 246 269
rect 212 185 246 201
rect 318 507 352 523
rect 318 439 352 445
rect 318 371 352 373
rect 318 335 352 337
rect 318 263 352 269
rect 318 185 352 201
rect 424 507 458 523
rect 424 439 458 445
rect 424 371 458 373
rect 424 335 458 337
rect 424 263 458 269
rect 424 185 458 201
rect 530 507 564 523
rect 530 439 564 445
rect 530 371 564 373
rect 530 335 564 337
rect 530 263 564 269
rect 530 185 564 201
rect 636 507 670 523
rect 636 439 670 445
rect 636 371 670 373
rect 636 335 670 337
rect 636 263 670 269
rect 636 185 670 201
rect 722 507 841 523
rect 756 479 790 507
rect 756 473 788 479
rect 824 473 841 507
rect 722 445 788 473
rect 822 445 841 473
rect 722 439 841 445
rect 756 407 790 439
rect 756 405 788 407
rect 824 405 841 439
rect 722 373 788 405
rect 822 373 841 405
rect 722 371 841 373
rect 756 337 790 371
rect 824 337 841 371
rect 722 335 841 337
rect 722 303 788 335
rect 822 303 841 335
rect 756 301 788 303
rect 756 269 790 301
rect 824 269 841 303
rect 722 263 841 269
rect 722 235 788 263
rect 822 235 841 263
rect 756 229 788 235
rect 756 201 790 229
rect 824 201 841 235
rect 722 185 841 201
rect 120 163 160 185
rect 722 163 762 185
rect 120 147 186 163
rect 120 113 136 147
rect 170 113 186 147
rect 696 147 762 163
rect 120 97 186 113
rect 266 125 616 139
rect 266 19 280 125
rect 602 19 616 125
rect 696 113 712 147
rect 746 113 762 147
rect 696 97 762 113
rect 266 0 616 19
<< viali >>
rect 280 687 602 689
rect 280 585 288 687
rect 288 585 594 687
rect 594 585 602 687
rect 280 583 602 585
rect 60 473 92 479
rect 92 473 94 479
rect 60 445 94 473
rect 60 405 92 407
rect 92 405 94 407
rect 60 373 94 405
rect 60 303 94 335
rect 60 301 92 303
rect 92 301 94 303
rect 60 235 94 263
rect 60 229 92 235
rect 92 229 94 235
rect 212 473 246 479
rect 212 445 246 473
rect 212 405 246 407
rect 212 373 246 405
rect 212 303 246 335
rect 212 301 246 303
rect 212 235 246 263
rect 212 229 246 235
rect 318 473 352 479
rect 318 445 352 473
rect 318 405 352 407
rect 318 373 352 405
rect 318 303 352 335
rect 318 301 352 303
rect 318 235 352 263
rect 318 229 352 235
rect 424 473 458 479
rect 424 445 458 473
rect 424 405 458 407
rect 424 373 458 405
rect 424 303 458 335
rect 424 301 458 303
rect 424 235 458 263
rect 424 229 458 235
rect 530 473 564 479
rect 530 445 564 473
rect 530 405 564 407
rect 530 373 564 405
rect 530 303 564 335
rect 530 301 564 303
rect 530 235 564 263
rect 530 229 564 235
rect 636 473 670 479
rect 636 445 670 473
rect 636 405 670 407
rect 636 373 670 405
rect 636 303 670 335
rect 636 301 670 303
rect 636 235 670 263
rect 636 229 670 235
rect 788 473 790 479
rect 790 473 822 479
rect 788 445 822 473
rect 788 405 790 407
rect 790 405 822 407
rect 788 373 822 405
rect 788 303 822 335
rect 788 301 790 303
rect 790 301 822 303
rect 788 235 822 263
rect 788 229 790 235
rect 790 229 822 235
rect 280 123 602 125
rect 280 21 288 123
rect 288 21 594 123
rect 594 21 602 123
rect 280 19 602 21
<< metal1 >>
rect 264 689 618 708
rect 264 583 280 689
rect 602 583 618 689
rect 264 571 618 583
rect 41 479 100 507
rect 41 445 60 479
rect 94 445 100 479
rect 41 407 100 445
rect 41 373 60 407
rect 94 373 100 407
rect 41 335 100 373
rect 41 301 60 335
rect 94 301 100 335
rect 41 263 100 301
rect 41 229 60 263
rect 94 229 100 263
rect 41 201 100 229
rect 203 479 255 507
rect 203 445 212 479
rect 246 445 255 479
rect 203 407 255 445
rect 203 373 212 407
rect 246 373 255 407
rect 203 335 255 373
rect 203 323 212 335
rect 246 323 255 335
rect 203 263 255 271
rect 203 259 212 263
rect 246 259 255 263
rect 203 201 255 207
rect 309 501 361 507
rect 309 445 318 449
rect 352 445 361 449
rect 309 437 361 445
rect 309 373 318 385
rect 352 373 361 385
rect 309 335 361 373
rect 309 301 318 335
rect 352 301 361 335
rect 309 263 361 301
rect 309 229 318 263
rect 352 229 361 263
rect 309 201 361 229
rect 415 479 467 507
rect 415 445 424 479
rect 458 445 467 479
rect 415 407 467 445
rect 415 373 424 407
rect 458 373 467 407
rect 415 335 467 373
rect 415 323 424 335
rect 458 323 467 335
rect 415 263 467 271
rect 415 259 424 263
rect 458 259 467 263
rect 415 201 467 207
rect 521 501 573 507
rect 521 445 530 449
rect 564 445 573 449
rect 521 437 573 445
rect 521 373 530 385
rect 564 373 573 385
rect 521 335 573 373
rect 521 301 530 335
rect 564 301 573 335
rect 521 263 573 301
rect 521 229 530 263
rect 564 229 573 263
rect 521 201 573 229
rect 627 479 679 507
rect 627 445 636 479
rect 670 445 679 479
rect 627 407 679 445
rect 627 373 636 407
rect 670 373 679 407
rect 627 335 679 373
rect 627 323 636 335
rect 670 323 679 335
rect 627 263 679 271
rect 627 259 636 263
rect 670 259 679 263
rect 627 201 679 207
rect 782 479 841 507
rect 782 445 788 479
rect 822 445 841 479
rect 782 407 841 445
rect 782 373 788 407
rect 822 373 841 407
rect 782 335 841 373
rect 782 301 788 335
rect 822 301 841 335
rect 782 263 841 301
rect 782 229 788 263
rect 822 229 841 263
rect 782 201 841 229
rect 264 125 618 137
rect 264 19 280 125
rect 602 19 618 125
rect 264 0 618 19
<< via1 >>
rect 203 301 212 323
rect 212 301 246 323
rect 246 301 255 323
rect 203 271 255 301
rect 203 229 212 259
rect 212 229 246 259
rect 246 229 255 259
rect 203 207 255 229
rect 309 479 361 501
rect 309 449 318 479
rect 318 449 352 479
rect 352 449 361 479
rect 309 407 361 437
rect 309 385 318 407
rect 318 385 352 407
rect 352 385 361 407
rect 415 301 424 323
rect 424 301 458 323
rect 458 301 467 323
rect 415 271 467 301
rect 415 229 424 259
rect 424 229 458 259
rect 458 229 467 259
rect 415 207 467 229
rect 521 479 573 501
rect 521 449 530 479
rect 530 449 564 479
rect 564 449 573 479
rect 521 407 573 437
rect 521 385 530 407
rect 530 385 564 407
rect 564 385 573 407
rect 627 301 636 323
rect 636 301 670 323
rect 670 301 679 323
rect 627 271 679 301
rect 627 229 636 259
rect 636 229 670 259
rect 670 229 679 259
rect 627 207 679 229
<< metal2 >>
rect 14 501 868 507
rect 14 449 309 501
rect 361 449 521 501
rect 573 449 868 501
rect 14 437 868 449
rect 14 385 309 437
rect 361 385 521 437
rect 573 385 868 437
rect 14 379 868 385
rect 14 323 868 329
rect 14 271 203 323
rect 255 271 415 323
rect 467 271 627 323
rect 679 271 868 323
rect 14 259 868 271
rect 14 207 203 259
rect 255 207 415 259
rect 467 207 627 259
rect 679 207 868 259
rect 14 201 868 207
<< labels >>
flabel comment s 183 365 183 365 0 FreeSans 180 90 0 0 dummy_poly
flabel comment s 693 352 693 352 0 FreeSans 180 90 0 0 dummy_poly
flabel metal1 s 321 606 571 656 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel metal1 s 321 42 571 92 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel metal1 s 41 339 87 369 0 FreeSans 200 90 0 0 SUBSTRATE
port 4 nsew
flabel metal1 s 795 339 841 369 0 FreeSans 200 90 0 0 SUBSTRATE
port 4 nsew
flabel metal2 s 14 201 35 329 7 FreeSans 300 180 0 0 SOURCE
port 3 nsew
flabel metal2 s 14 379 35 507 7 FreeSans 300 180 0 0 DRAIN
port 1 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 5533936
string GDS_START 5518500
<< end >>
