* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__nfet_01v8__toxe_slope_spectre = 0.0
.param sky130_fd_pr__nfet_01v8__vth0_slope_spectre = 0.0
.param sky130_fd_pr__nfet_01v8__voff_slope_spectre = 0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__nfet_01v8__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_01v8__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_01v8__voff_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt  sky130_fd_pr__nfet_01v8 d g s b
+ 
.param  l = 1 w = 1 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1 
msky130_fd_pr__nfet_01v8 d g s b sky130_fd_pr__nfet_01v8__model l = {l} w = {w} nf = {nf} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd} 
.model sky130_fd_pr__nfet_01v8__model.0 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {0.521494355+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.54086565
+ k2 = -0.026725491
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.1052686+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 2.5784
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0319905
+ ua = -7.5751847e-10
+ ub = 1.734885e-18
+ uc = 4.9242e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.314494
+ ags = 0.423558
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 2.1073424e-24
+ keta = -0.0087946
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.026316
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0030734587
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 754674160.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.31303
+ kt2 = -0.045313337
+ at = 140000.0
+ ute = -1.8134
+ ua1 = 3.7602e-10
+ ub1 = -6.3962e-19
+ uc1 = 1.5829713e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.1 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {0.521494355+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.54086565
+ k2 = -0.026725491
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.1052686+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 2.5784
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0319905
+ ua = -7.5751847e-10
+ ub = 1.734885e-18
+ uc = 4.9242e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.314494
+ ags = 0.423558
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 2.1073424e-24
+ keta = -0.0087946
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.026316
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0030734587
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 754674160.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.31303
+ kt2 = -0.045313337
+ at = 140000.0
+ ute = -1.8134
+ ua1 = 3.7602e-10
+ ub1 = -6.3962e-19
+ uc1 = 1.5829713e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.2 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.218129600e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -2.533509204e-09 wvth0 = -3.186707545e-08 pvth0 = 2.534031918e-13
+ k1 = 5.415479012e-01 lk1 = -5.425180173e-09 wk1 = -6.823919393e-08 pk1 = 5.426299497e-13
+ k2 = -2.720722062e-02 lk2 = 3.830656641e-09 wk2 = 4.818290141e-08 pk2 = -3.831446982e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.049986455e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.146645748e-09 wvoff = -2.700101578e-08 pvoff = 2.147088644e-13
+ nfactor = 2.583165078e+00 lnfactor = -3.789133339e-08 wnfactor = -4.766061153e-07 pnfactor = 3.789915113e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.198065511e-02 lu0 = 7.828542819e-11 wu0 = 9.846925531e-10 pu0 = -7.830158004e-15
+ ua = -7.571315321e-10 lua = -3.076884210e-18 wua = -3.870177424e-17 pua = 3.077519033e-22
+ ub = 1.735654766e-18 lub = -6.121090184e-27 wub = -7.699251394e-26 pub = 6.122353088e-31
+ uc = 4.876862466e-11 luc = 3.764224339e-18 wuc = 4.734730026e-17 puc = -3.765000973e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.308117268e+00 la0 = 5.070701382e-08 wa0 = 6.378047621e-07 pa0 = -5.071747569e-12
+ ags = 4.237412493e-01 lags = -1.457176493e-09 wags = -1.832870911e-08 pags = 1.457477137e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 1.950171466e-24 lb1 = 1.249804562e-30 wb1 = 1.572033612e-29 pb1 = -1.250062421e-34
+ keta = -8.286491579e-03 lketa = -4.040417702e-09 wketa = -5.082132543e-08 pketa = 4.041251321e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.813472448e-02 lpclm = -3.325375207e-07 wpclm = -4.182735252e-06 ppclm = 3.326061298e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 3.074736097e-03 lpdiblc2 = -1.015771223e-11 wpdiblc2 = -1.277660967e-10 ppdiblc2 = 1.015980797e-15
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 7.580546759e+08 lpscbe1 = -2.688146055e+01 wpscbe1 = -3.381213417e+02 ppscbe1 = 2.688700673e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.131873691e-01 lkt1 = 1.251380708e-09 wkt1 = 1.574016127e-08 pkt1 = -1.251638893e-13
+ kt2 = -4.539697534e-02 lkt2 = 6.650821582e-10 wkt2 = 8.365560022e-09 pkt2 = -6.652193779e-14
+ at = 140000.0
+ ute = -1.816368385e+00 lute = 2.360424274e-08 wute = 2.968997243e-07 pute = -2.360911277e-12
+ ua1 = 3.613302243e-10 lua1 = 1.168113480e-16 wua1 = 1.469280646e-15 pua1 = -1.168354485e-20
+ ub1 = -6.203888939e-19 lub1 = -1.529234671e-25 wub1 = -1.923507385e-24 pub1 = 1.529550183e-29
+ uc1 = 1.691322611e-11 luc1 = -8.615967309e-18 wuc1 = -1.083736660e-16 puc1 = 8.617744955e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.3 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.172193813e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.561976709e-08 wvth0 = 1.059289624e-08 pvth0 = 8.560643642e-14
+ k1 = 5.305642003e-01 lk1 = 3.798109855e-08 wk1 = 1.374219832e-07 pk1 = -2.701185486e-13
+ k2 = -1.951904366e-02 lk2 = -2.655210381e-08 wk2 = -9.030202569e-08 pk2 = 1.641312539e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 5.378976803e-01 ldsub = 8.734573725e-08 wdsub = 2.210687984e-06 pdsub = -8.736375842e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.093607521e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.509188017e-08 wvoff = 5.598118683e-08 pvoff = -1.132269255e-13
+ nfactor = 2.513649424e+00 lnfactor = 2.368262590e-07 wnfactor = 2.398232180e-07 pnfactor = 9.586716424e-13
+ eta0 = 7.414288528e-02 leta0 = 2.314662037e-08 weta0 = 5.858323158e-07 peta0 = -2.315139598e-12
+ etab = -6.487968019e-02 letab = -2.023489459e-08 wetab = -5.121376239e-07 petab = 2.023906945e-12
+ u0 = 3.200913334e-02 lu0 = -3.425715201e-11 wu0 = 1.102135439e-08 pu0 = -4.749385120e-14
+ ua = -7.760011693e-10 lua = 7.149367668e-17 wua = 1.342223993e-15 pua = -5.149502397e-21
+ ub = 1.731569260e-18 lub = 1.002434650e-26 wub = -6.758335518e-25 pub = 2.978783828e-30
+ uc = 5.869782097e-11 luc = -3.547477787e-17 wuc = -3.262199531e-16 puc = 1.099793233e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.407957701e+00 la0 = -3.438504978e-07 wa0 = -1.002383227e-06 pa0 = 1.410080182e-12
+ ags = 4.347153216e-01 lags = -4.482540441e-08 wags = -1.355800413e-06 pags = 5.431276727e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 4.478325063e-24 lb1 = -8.741157602e-30 wb1 = -3.144067224e-29 pb1 = 6.136845078e-35
+ keta = -1.632297162e-02 lketa = 2.771879508e-08 wketa = 8.797632511e-08 pketa = -1.443866660e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -6.065884966e-01 lpclm = 2.333888357e-06 wpclm = 8.570843418e-06 ppclm = -1.714001225e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 3.181049172e-03 lpdiblc2 = -4.302943326e-10 wpdiblc2 = -1.243313447e-08 ppdiblc2 = 4.964533227e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 7.036778051e+08 lpscbe1 = 1.880094620e+02 wpscbe1 = 6.762426835e+02 ppscbe1 = -1.319945245e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.113073089e-01 lkt1 = -6.178393478e-09 wkt1 = 3.366128340e-08 pkt1 = -1.959860314e-13
+ kt2 = -4.405263989e-02 lkt2 = -4.647571595e-09 wkt2 = -1.662922207e-08 pkt2 = 3.225446664e-14
+ at = 1.381537196e+05 lat = 7.296280585e-03 wat = 1.846661363e-01 pat = -7.297785953e-7
+ ute = -1.758431629e+00 lute = -2.053549213e-07 wute = -1.612926609e-06 pute = 5.186495125e-12
+ ua1 = 6.201857871e-10 lua1 = -9.061550323e-16 wua1 = -5.195526344e-15 pua1 = 1.465497926e-20
+ ub1 = -9.432506693e-19 lub1 = 1.122987849e-24 wub1 = 5.199513679e-24 pub1 = -1.285382978e-29
+ uc1 = -6.765134883e-14 luc1 = 5.849043968e-17 wuc1 = 1.719542394e-16 puc1 = -2.460480276e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.4 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.269226307e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.319821014e-09 wvth0 = -1.156669319e-07 pvth0 = 3.320505960e-13
+ k1 = 5.524481767e-01 lk1 = -4.733819062e-09 wk1 = -2.435429029e-07 pk1 = 4.734795743e-13
+ k2 = -3.403716059e-02 lk2 = 1.785532771e-09 wk2 = 8.528315095e-08 pk2 = -1.785901162e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 5.826472000e-01 wdsub = -2.265187257e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.029738619e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.625430530e-09 wvoff = 1.325075199e-07 pvoff = -2.625972209e-13
+ nfactor = 2.626480551e+00 lnfactor = 1.659332642e-08 wnfactor = 1.581271102e-06 pnfactor = -1.659674996e-12
+ eta0 = 8.614746983e-02 leta0 = -2.849001211e-10 weta0 = -6.148738175e-07 peta0 = 2.849589016e-14
+ etab = -7.523302611e-02 letab = -2.639540117e-11 wetab = 5.234105783e-07 petab = 2.640084707e-15
+ u0 = 3.168571117e-02 lu0 = 5.970244211e-10 wu0 = 1.728244751e-08 pu0 = -5.971475991e-14
+ ua = -7.764945590e-10 lua = 7.245671468e-17 wua = 2.416912458e-15 pua = -7.247166394e-21
+ ub = 1.767613406e-18 lub = -6.032953795e-26 wub = -2.241202899e-24 pub = 6.034198514e-30
+ uc = 3.955731360e-11 luc = 1.885214783e-18 wuc = 3.338375030e-16 puc = -1.885603740e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.145872006e+04 lvsat = -2.847247979e-03 wvsat = -1.459021028e-01 pvsat = 2.847835423e-7
+ a0 = 1.225512924e+00 la0 = 1.225999733e-08 wa0 = 3.482794738e-07 pa0 = -1.226252682e-12
+ ags = 4.303748814e-01 lags = -3.635338168e-08 wags = -4.360780954e-07 pags = 3.636088211e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -6.788693384e-03 lketa = 9.109018544e-09 wketa = 4.807785122e-07 pketa = -9.110897917e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.770898436e-01 lpclm = 2.348909453e-08 wpclm = 9.932205155e-07 ppclm = -2.349394080e-12
+ pdiblc1 = 4.127907046e-01 lpdiblc1 = -4.448474321e-08 wpdiblc1 = -2.279540674e-06 ppdiblc1 = 4.449392130e-12
+ pdiblc2 = 2.903034209e-03 lpdiblc2 = 1.123577912e-10 wpdiblc2 = 1.875904864e-08 ppdiblc2 = -1.123809728e-14
+ pdiblcb = -2.321731417e-02 lpdiblcb = -3.479590594e-09 wpdiblcb = -1.783053630e-07 ppdiblcb = 3.480308503e-13
+ drout = 5.384425606e-01 ldrout = 4.207755634e-08 wdrout = 2.156188711e-06 pdrout = -4.208623778e-12
+ pscbe1 = 7.612738250e+08 lpscbe1 = 7.558888522e+01 wpscbe1 = 3.873416500e+03 ppscbe1 = -7.560448072e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.175497226e-07 lalpha0 = -3.660747402e-13 walpha0 = -1.875884179e-11 palpha0 = 3.661502687e-17
+ alpha1 = 8.524431765e-01 lalpha1 = -4.768789719e-09 walpha1 = -2.443680540e-07 palpha1 = 4.769773615e-13
+ beta0 = 1.405919074e+01 lbeta0 = -3.887966206e-07 wbeta0 = -1.992318369e-05 pbeta0 = 3.888768371e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.107870590e-01 lkt1 = -7.193859549e-09 wkt1 = -4.353839145e-07 pkt1 = 7.195343786e-13
+ kt2 = -4.499211016e-02 lkt2 = -2.813837418e-09 wkt2 = -1.442944487e-07 pkt2 = 2.814417968e-13
+ at = 1.381857848e+05 lat = 7.233692969e-03 wat = 1.814589465e-01 pat = -7.235185425e-7
+ ute = -1.804136022e+00 lute = -1.161453856e-07 wute = -4.907410108e-06 pute = 1.161693487e-11
+ ua1 = 2.794532101e-10 lua1 = -2.410855892e-16 wua1 = -1.004139232e-14 pua1 = 2.411353299e-20
+ ub1 = -4.327624759e-19 lub1 = 1.265756432e-25 wub1 = 5.100299665e-24 pub1 = -1.266017583e-29
+ uc1 = 3.129483059e-11 luc1 = -2.725392919e-18 wuc1 = -9.376049924e-17 puc1 = 2.725955222e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.5 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.171125310e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.018226499e-09 wvth0 = 2.136630052e-07 pvth0 = 1.856768615e-14
+ k1 = 5.409208001e-01 lk1 = 6.238871633e-09 wk1 = 9.210076425e-07 pk1 = -6.350339634e-13
+ k2 = -2.872661670e-02 lk2 = -3.269473057e-09 wk2 = -3.714966036e-07 pk2 = 2.562098533e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.834881500e-01 ldsub = -2.863647844e-07 wdsub = -5.237035285e-06 pdsub = 2.828845673e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.008853338e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 6.374003522e-10 wvoff = -5.211012878e-08 pvoff = -8.686318891e-14
+ nfactor = 2.558418908e+00 lnfactor = 8.137991121e-08 wnfactor = -3.622854331e-07 pnfactor = 1.903595430e-13
+ eta0 = 1.963790274e-01 leta0 = -1.052122254e-07 weta0 = -4.453913582e-06 peta0 = 3.682804900e-12
+ etab = -1.428132220e-01 letab = 6.430190908e-08 wetab = 1.000445129e-06 petab = -4.514400406e-13
+ u0 = 3.383241305e-02 lu0 = -1.446380308e-09 wu0 = -3.807495614e-08 pu0 = -7.021099164e-15
+ ua = -5.446606297e-10 lua = -1.482215978e-16 wua = -5.255743085e-15 pua = 5.628863722e-23
+ ub = 1.593961595e-18 lub = 1.049663211e-25 wub = 4.948197280e-24 pub = -8.092549166e-31
+ uc = 1.249145366e-11 luc = 2.764869261e-17 wuc = 2.008662409e-16 puc = -6.198755604e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.887838036e+04 lvsat = -3.910716404e-04 wvsat = 1.121851053e-01 pvsat = 3.911523263e-8
+ a0 = 1.301414784e+00 la0 = -5.998954116e-08 wa0 = -3.891812428e-06 pa0 = 2.809810238e-12
+ ags = 2.341559776e-01 lags = 1.504236647e-07 wags = 2.108615474e-06 pags = 1.213842752e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 3.585808579e-03 lketa = -7.662727592e-10 wketa = -7.245302051e-07 pketa = 2.362206755e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.387428945e-01 lpclm = -3.519727316e-08 wpclm = -2.654052225e-06 ppclm = 1.122375543e-12
+ pdiblc1 = 3.860362044e-01 lpdiblc1 = -1.901764281e-08 wpdiblc1 = 3.964613441e-07 ppdiblc1 = 1.902156653e-12
+ pdiblc2 = 1.307411195e-03 lpdiblc2 = 1.631201021e-09 wpdiblc2 = 2.270271598e-08 ppdiblc2 = -1.499199929e-14
+ pdiblcb = -2.856537165e-02 lpdiblcb = 1.611123708e-09 wpdiblcb = 3.566107261e-07 ppdiblcb = -1.611456115e-13
+ drout = 5.989362241e-01 ldrout = -1.550521253e-08 wdrout = -3.894425740e-06 pdrout = 1.550841156e-12
+ pscbe1 = 8.611341629e+08 lpscbe1 = -1.946627312e+01 wpscbe1 = -6.114677612e+03 ppscbe1 = 1.947028940e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 6.220736218e-08 lalpha0 = -2.182072988e-13 walpha0 = -3.221400721e-12 palpha0 = 2.182523193e-17
+ alpha1 = 8.451136471e-01 lalpha1 = 2.208050047e-09 walpha1 = 4.887361079e-07 palpha1 = -2.208505612e-13
+ beta0 = 1.379865296e+01 lbeta0 = -1.407956618e-07 wbeta0 = 6.135969324e-06 pbeta0 = 1.408247108e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.100292044e-01 lkt1 = -7.915246926e-09 wkt1 = 2.879054336e-07 pkt1 = 3.104899066e-14
+ kt2 = -4.859593454e-02 lkt2 = 6.165745338e-10 wkt2 = 2.174123230e-07 pkt2 = -6.286000670e-14
+ at = 1.694651349e+05 lat = -2.254052607e-02 wat = -6.818265665e-01 pat = 9.822653489e-8
+ ute = -2.097439592e+00 lute = 1.630447101e-07 wute = 1.192739109e-05 pute = -4.407792531e-12
+ ua1 = -3.453099276e-10 lua1 = 3.536145712e-16 wua1 = 2.476167800e-14 pua1 = -9.014848391e-21
+ ub1 = -1.030730348e-19 lub1 = -1.872494717e-25 wub1 = -1.128437649e-23 pub1 = 2.936086094e-30
+ uc1 = 1.777556596e-11 luc1 = 1.014333821e-17 wuc1 = 7.089691523e-16 puc1 = -4.915075813e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.6 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.273663950e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.384700175e-09 wvth0 = 5.612462690e-07 pvth0 = -1.384985867e-13
+ k1 = 5.715529117e-01 lk1 = -7.603197571e-09 wk1 = -2.167218217e-06 pk1 = 7.604766262e-13
+ k2 = -4.015512610e-02 lk2 = 1.894853201e-09 wk2 = 6.149008506e-07 pk2 = -1.895244147e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.596726871e-01 ldsub = -4.474429138e-09 wdsub = 3.273804614e-08 pdsub = 4.475352302e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-9.996576440e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.218644100e-10 wvoff = -1.952278310e-07 pvoff = -2.219101850e-14
+ nfactor = 2.723311816e+00 lnfactor = 6.867938774e-09 wnfactor = 1.579144102e-06 pnfactor = -6.869355767e-13
+ eta0 = -3.645268133e-02 weta0 = 3.696030541e-6
+ etab = -5.500922860e-04 letab = 1.590374692e-11 wetab = 4.941140841e-09 petab = -1.590702818e-15
+ u0 = 3.035087852e-02 lu0 = 1.268589979e-10 wu0 = -2.553311884e-08 pu0 = -1.268851715e-14
+ ua = -9.050069043e-10 lua = 1.461203710e-17 wua = -1.896907855e-15 pua = -1.461505186e-21
+ ub = 1.848530684e-18 lub = -1.006861344e-26 wub = 9.287231345e-25 pub = 1.007069080e-30
+ uc = 7.378934263e-11 luc = -5.065875470e-20 wuc = 5.247656150e-17 puc = 5.066920662e-24
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.889396347e+04 lvsat = -3.981133522e-04 wvsat = 1.106264726e-01 pvsat = 3.981954910e-8
+ a0 = 1.168659609e+00 wa0 = 2.326218952e-6
+ ags = 4.920292993e-01 lags = 3.389561025e-08 wags = 1.229736674e-05 pags = -3.390260359e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.176432020e-03 lketa = 3.224787296e-10 wketa = -1.304021010e-07 pketa = -3.225452634e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.532560235e-01 lpclm = 3.432619589e-09 wpclm = 5.895192546e-07 ppclm = -3.433327807e-13
+ pdiblc1 = 2.901930816e-01 lpdiblc1 = 2.429204335e-08 wpdiblc1 = 9.982751056e-06 ppdiblc1 = -2.429705528e-12
+ pdiblc2 = 4.863234098e-03 lpdiblc2 = 2.439221243e-11 wpdiblc2 = -5.075116665e-09 ppdiblc2 = -2.439724503e-15
+ pdiblcb = -3.719210502e-02 lpdiblcb = 5.509380609e-09 wpdiblcb = 1.219462050e-06 ppdiblcb = -5.510517305e-13
+ drout = 5.951799404e-01 ldrout = -1.380781932e-08 wdrout = -3.518719875e-06 pdrout = 1.381066814e-12
+ pscbe1 = 8.326363742e+08 lpscbe1 = -6.588663863e+00 wpscbe1 = -3.264310775e+03 ppscbe1 = 6.590023236e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.255066444e-07 lalpha0 = 9.255759424e-14 walpha0 = 6.556418885e-11 palpha0 = -9.257669072e-18
+ alpha1 = 0.85
+ beta0 = 1.350701020e+01 lbeta0 = -9.007837296e-09 wbeta0 = 3.530626305e-05 pbeta0 = 9.009695793e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.284544700e-01 lkt1 = 4.107805201e-10 wkt1 = 4.475393148e-07 pkt1 = -4.108652723e-14
+ kt2 = -4.746758796e-02 lkt2 = 1.066961524e-10 wkt2 = 1.019213196e-07 pkt2 = -1.067181660e-14
+ at = 1.179069490e+05 lat = 7.576385343e-04 wat = -2.967561167e-01 pat = -7.577948503e-8
+ ute = -1.702597379e+00 lute = -1.537698402e-08 wute = -1.230515948e-06 pute = 1.538015660e-12
+ ua1 = 4.578239744e-10 lua1 = -9.306379613e-18 wua1 = 2.752170275e-15 pua1 = 9.308299705e-22
+ ub1 = -4.911172607e-19 lub1 = -1.189965884e-26 wub1 = -7.420804672e-24 pub1 = 1.190211398e-30
+ uc1 = 4.654934639e-11 luc1 = -2.858986461e-18 wuc1 = -1.011539597e-15 puc1 = 2.859576327e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.7 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.229406475e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.278174521e-09 wvth0 = 1.003912338e-06 pvth0 = -2.278644554e-13
+ k1 = 5.516656744e-01 lk1 = -3.588342226e-09 wk1 = -1.780841779e-07 pk1 = 3.589082573e-13
+ k2 = -3.408768906e-02 lk2 = 6.699529435e-10 wk2 = 8.031963081e-09 pk2 = -6.700911682e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.148966321e-01 ldsub = 4.565005612e-09 wdsub = 4.511267361e-06 pdsub = -4.565947464e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.006486646e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 3.597289941e-10 wvoff = -1.269237170e-07 pvoff = -3.598032134e-14
+ nfactor = 2.844957734e+00 lnfactor = -1.769006076e-08 wnfactor = -1.058795748e-05 pnfactor = 1.769371058e-12
+ eta0 = -1.017366340e-01 leta0 = 1.317958964e-08 weta0 = 1.022577274e-05 peta0 = -1.318230885e-12
+ etab = -4.377919339e-03 letab = 7.886693003e-10 wetab = 3.878028219e-07 petab = -7.888320185e-14
+ u0 = 3.223541334e-02 lu0 = -2.535927756e-10 wu0 = -2.140254823e-07 pu0 = 2.536450969e-14
+ ua = -6.344417395e-10 lua = -4.000992895e-17 wua = -2.895900664e-14 pua = 4.001818380e-21
+ ub = 1.644104504e-18 lub = 3.120114826e-26 wub = 2.137555888e-23 pub = -3.120758568e-30
+ uc = 7.379597926e-11 luc = -5.199856395e-20 wuc = 5.181276169e-17 puc = 5.200929230e-24
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.832386026e+04 lvsat = -2.830203450e-04 wvsat = 1.676485565e-01 pvsat = 2.830787378e-8
+ a0 = 1.168659609e+00 wa0 = 2.326218952e-6
+ ags = 8.349323227e-01 lags = -3.532999502e-08 wags = -2.200001038e-05 pags = 3.533728431e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.676169291e-03 lketa = 1.971026958e-11 wketa = -2.804067707e-07 pketa = -1.971433620e-15
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.524013734e-01 lpclm = 3.605157200e-09 wpclm = 6.750018952e-07 ppclm = -3.605901016e-13
+ pdiblc1 = 4.470333421e-01 lpdiblc1 = -7.371025280e-09 wpdiblc1 = -5.704510921e-06 ppdiblc1 = 7.372546070e-13
+ pdiblc2 = 5.878611694e-03 lpdiblc2 = -1.805932321e-10 wpdiblc2 = -1.066338256e-07 ppdiblc2 = 1.806304921e-14
+ pdiblcb = 9.816828002e-03 lpdiblcb = -3.980829798e-09 wpdiblcb = -3.482401141e-06 ppdiblcb = 3.981651123e-13
+ drout = 4.865202783e-01 ldrout = 8.128501942e-09 wdrout = 7.349488207e-06 pdrout = -8.130179015e-13
+ pscbe1 = 7.994163763e+08 lpscbe1 = 1.178225440e-01 wpscbe1 = 5.837441519e+01 ppscbe1 = -1.178468531e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.411118510e-07 lalpha0 = 7.551988896e-14 walpha0 = 5.712296828e-11 palpha0 = -7.553547023e-18
+ alpha1 = 8.985131162e-01 lalpha1 = -9.793876402e-09 walpha1 = -4.852312538e-06 palpha1 = 9.795897075e-13
+ beta0 = 1.287542604e+01 lbeta0 = 1.184970036e-07 wbeta0 = 9.847770942e-05 pbeta0 = -1.185214519e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.217926112e-01 lkt1 = -9.341221868e-10 wkt1 = -2.187840080e-07 pkt1 = 9.343149149e-14
+ kt2 = -4.640002116e-02 lkt2 = -1.088252994e-10 wkt2 = -4.857385744e-09 pkt2 = 1.088477522e-14
+ at = 1.230880761e+05 lat = -2.883325827e-04 wat = -8.149757222e-01 pat = 2.883920714e-8
+ ute = -1.914671295e+00 lute = 2.743671035e-08 wute = 1.998125123e-05 pute = -2.744237109e-12
+ ua1 = 1.250765445e-10 lua1 = 5.786900428e-17 wua1 = 3.603377851e-14 pua1 = -5.788094381e-21
+ ub1 = -3.105051378e-19 lub1 = -4.836181482e-26 wub1 = -2.548574335e-23 pub1 = 4.837179283e-30
+ uc1 = 3.829960631e-11 luc1 = -1.193520684e-18 wuc1 = -1.863953801e-16 puc1 = 1.193766931e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.8 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.273923193e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.691083593e-09 wvth0 = 5.586533116e-07 pvth0 = -1.691432497e-13
+ k1 = 5.285591841e-01 lk1 = -5.410351761e-10 wk1 = 2.133041587e-06 pk1 = 5.411468025e-14
+ k2 = -2.795698838e-02 lk2 = -1.385699937e-10 wk2 = -6.051645941e-07 pk2 = 1.385985834e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.309471627e-01 ldsub = 2.448245588e-09 wdsub = 2.905883148e-06 pdsub = -2.448750710e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 4.015608772e-03 lcdscd = 1.825749525e-10 wcdscd = 1.384677258e-07 pcdscd = -1.826126214e-14
+ cit = 0.0
+ voff = {-1.140722216e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.130041113e-09 wvoff = 1.215708936e-06 pvoff = -2.130480583e-13
+ nfactor = 2.404810399e+00 lnfactor = 4.035700990e-08 wnfactor = 3.343585712e-05 pnfactor = -4.036533636e-12
+ eta0 = -9.543751350e-03 leta0 = 1.021100089e-09 weta0 = 1.004582358e-06 peta0 = -1.021310763e-13
+ etab = -2.046012849e-03 letab = 4.811351404e-10 wetab = 1.545640610e-07 petab = -4.812344083e-14
+ u0 = 2.729167991e-02 lu0 = 3.983917324e-10 wu0 = 2.804498594e-07 pu0 = -3.984739286e-14
+ ua = -1.361176209e-09 lua = 5.583253961e-17 wua = 4.372943428e-14 pua = -5.584405897e-21
+ ub = 2.230433597e-18 lub = -4.612451884e-26 wub = -3.726944755e-23 pub = 4.613403526e-30
+ uc = 6.487204827e-11 luc = 1.124898379e-18 wuc = 9.443899792e-16 puc = -1.125130468e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.974571693e+04 lvsat = -4.705362249e-04 wvsat = 2.543355348e-02 pvsat = 4.706333060e-8
+ a0 = 1.168659609e+00 wa0 = 2.326218952e-6
+ ags = 5.670393357e-01 wags = 4.794815495e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.865639891e-02 lketa = -2.087778393e-09 wketa = -1.878759436e-06 pketa = 2.088209143e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.497580448e-01 lpclm = 3.953762028e-09 wpclm = 9.393892987e-07 ppclm = -3.954577768e-13
+ pdiblc1 = 3.941760871e-01 lpdiblc1 = -4.001576379e-10 wpdiblc1 = -4.176948735e-07 ppdiblc1 = 4.002401985e-14
+ pdiblc2 = 4.694446634e-03 lpdiblc2 = -2.442435986e-11 wpdiblc2 = 1.180711210e-08 ppdiblc2 = 2.442939909e-15
+ pdiblcb = 1.768372043e-03 lpdiblcb = -2.919391378e-09 wpdiblcb = -2.677389489e-06 ppdiblcb = 2.919993707e-13
+ drout = 5.019275418e-01 ldrout = 6.096576626e-09 wdrout = 5.808443976e-06 pdrout = -6.097834471e-13
+ pscbe1 = 7.989354065e+08 lpscbe1 = 1.812533128e-01 wpscbe1 = 1.064813114e+02 ppscbe1 = -1.812907089e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.670289792e-08 lalpha0 = -6.828979429e-16 walpha0 = -6.704280861e-13 palpha0 = 6.830388384e-20
+ alpha1 = 7.368027290e-01 lalpha1 = 1.153265117e-08 walpha1 = 1.132206259e-05 palpha1 = -1.153503059e-12
+ beta0 = 1.348168018e+01 lbeta0 = 3.854360109e-08 wbeta0 = 3.783978701e-05 pbeta0 = -3.855155341e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.176701731e-01 lkt1 = -1.477793447e-09 wkt1 = -6.311128733e-07 pkt1 = 1.478098346e-13
+ kt2 = -4.550045638e-02 lkt2 = -2.274608018e-10 wkt2 = -9.483242330e-08 pkt2 = 2.275077315e-14
+ at = 1.200717910e+05 lat = 1.094581132e-04 wat = -5.132849798e-01 pat = -1.094806966e-8
+ ute = -1.238897372e+00 lute = -6.168503042e-08 wute = -4.761008367e-05 pute = 6.169775728e-12
+ ua1 = 1.215299084e-09 lua1 = -8.591063445e-17 wua1 = -7.301096891e-14 pua1 = 8.592835954e-21
+ ub1 = -1.050533218e-18 lub1 = 4.923382844e-26 wub1 = 4.853233294e-23 pub1 = -4.924398636e-30
+ uc1 = 3.621735192e-11 luc1 = -9.189108935e-19 wuc1 = 2.187301941e-17 puc1 = 9.191004832e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.9 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.181802239e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.312536362e-07 wvth0 = 2.326729478e-08 pvth0 = -2.325609879e-12
+ k1 = 5.418283439e-01 lk1 = -9.622306586e-08 wk1 = -6.758719581e-09 pk1 = 6.755467353e-13
+ k2 = -2.562399133e-02 lk2 = -1.100969642e-07 wk2 = -7.733223846e-09 pk2 = 7.729502696e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.045248049e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.434371986e-08 wvoff = -5.221911719e-09 pvoff = 5.219398987e-13
+ nfactor = 2.825822499e+00 lnfactor = -2.473034417e-05 wnfactor = -1.737062314e-06 pnfactor = 1.736226457e-10
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.133419179e-02 lu0 = 6.559924037e-08 wu0 = 4.607698440e-09 pu0 = -4.605481261e-13
+ ua = -7.330860930e-10 lua = -2.442062039e-15 wua = -1.715307278e-16 pua = 1.714481890e-20
+ ub = 1.660844193e-18 lub = 7.400517948e-24 wub = 5.198132601e-25 pub = -5.195631312e-29
+ uc = 4.770249614e-11 luc = 1.538763065e-16 wuc = 1.080829005e-17 puc = -1.080308921e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.338536054e+00 la0 = -2.403048544e-06 wa0 = -1.687904153e-07 pa0 = 1.687091951e-11
+ ags = 4.157296323e-01 lags = 7.824600798e-07 wags = 5.496008899e-08 pags = -5.493364275e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 7.880004902e-25 lb1 = 1.318707056e-28 wb1 = 9.262614031e-30 pb1 = -9.258156954e-34
+ keta = -7.162031474e-03 lketa = -1.631782950e-07 wketa = -1.146166284e-08 pketa = 1.145614760e-12
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.797380891e-02 lpclm = -3.164257549e-06 wpclm = -2.222578263e-07 ppclm = 2.221508781e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 3.148731110e-03 lpdiblc2 = -7.523618993e-09 wpdiblc2 = -5.284598922e-10 ppdiblc2 = 5.282056026e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 7.170199491e+08 lpscbe1 = 3.763609205e+03 wpscbe1 = 2.643563578e+02 ppscbe1 = -2.642291522e-2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.201484054e-01 lkt1 = 7.114980092e-07 wkt1 = 4.997570472e-08 pkt1 = -4.995165691e-12
+ kt2 = -4.543615047e-02 lkt2 = 1.227543698e-08 wkt2 = 8.622281524e-10 pkt2 = -8.618132568e-14
+ at = 140000.0
+ ute = -1.857412656e+00 lute = 4.399147761e-06 wute = 3.089966616e-07 pute = -3.088479755e-11
+ ua1 = 3.028200036e-10 lua1 = 7.316477330e-15 wua1 = 5.139102371e-16 pua1 = -5.136629487e-20
+ ub1 = -5.508621871e-19 lub1 = -8.871510358e-24 wub1 = -6.231359418e-25 pub1 = 6.228360950e-29
+ uc1 = 1.657925166e-11 luc1 = -7.491779926e-17 wuc1 = -5.262235124e-18 puc1 = 5.259702989e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.10 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.347828508e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = -9.329363894e-8
+ k1 = 5.370055873e-01 wk1 = 2.710007976e-8
+ k2 = -3.114211587e-02 wk2 = 3.100749787e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.082509558e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = 2.093802271e-8
+ nfactor = 1.586323117e+00 wnfactor = 6.965006713e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.462206426e-02 wu0 = -1.847524427e-8
+ ua = -8.554836774e-10 wua = 6.877776701e-16
+ ub = 2.031762501e-18 wub = -2.084267684e-24
+ uc = 5.541486704e-11 wuc = -4.333742790e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.218093849e+00 wa0 = 6.767899843e-7
+ ags = 4.549469913e-01 wags = -2.203705565e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 7.397437744e-24 wb1 = -3.713981266e-29
+ keta = -1.534062351e-02 wketa = 4.595722212e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.006206389e-01 wpclm = 8.911754287e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.771642905e-03 wpdiblc2 = 2.118937627e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 9.056542541e+08 wpscbe1 = -1.059975680e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.844877071e-01 wkt1 = -2.003849350e-7
+ kt2 = -4.482089835e-02 wkt2 = -3.457230533e-9
+ at = 140000.0
+ ute = -1.636924785e+00 wute = -1.238967540e-6
+ ua1 = 6.695261467e-10 wua1 = -2.060598646e-15
+ ub1 = -9.955074993e-19 wub1 = 2.498555166e-24
+ uc1 = 1.282432754e-11 wuc1 = 2.109970533e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.11 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.439583902e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.296279764e-08 wvth0 = -1.873419915e-07 pvth0 = 7.478613079e-13
+ k1 = 5.246951187e-01 lk1 = 9.789138099e-08 wk1 = 5.007798974e-08 pk1 = -1.827176058e-13
+ k2 = -2.829774244e-02 lk2 = -2.261811904e-08 wk2 = 5.583905375e-08 pk2 = -1.974575774e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.176997976e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 7.513606508e-08 wvoff = 6.216909851e-08 pvoff = -3.278646083e-13
+ nfactor = 4.853469164e-01 lnfactor = 8.754831730e-06 wnfactor = 1.425140320e-05 pnfactor = -5.794055779e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.698210199e-02 lu0 = -1.876673918e-08 wu0 = -3.412862550e-08 pu0 = 1.244738248e-13
+ ua = -8.958090789e-10 lua = 3.206627938e-16 wua = 9.349022485e-16 pua = -1.965105240e-21
+ ub = 2.237502053e-18 lub = -1.636016432e-24 wub = -3.600277633e-24 pub = 1.205513070e-29
+ uc = 1.762669439e-10 luc = -9.610013340e-16 wuc = -8.477714799e-16 puc = 6.396763854e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.533573376e+00 la0 = -2.508655659e-06 wa0 = -9.450396069e-07 pa0 = 1.289659591e-11
+ ags = 6.131245190e-01 lags = -1.257808877e-06 wags = -1.347918953e-06 pags = 8.966130668e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 1.470588616e-23 lb1 = -5.811591211e-29 wb1 = -7.383284265e-29 pb1 = 2.917786081e-34
+ keta = -2.858576715e-02 lketa = 1.053238060e-07 wketa = 9.169241821e-08 pketa = -3.636808368e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.019940503e+00 lpclm = 7.310322164e-06 wpclm = 3.456240511e-06 ppclm = -2.039709229e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 2.811239553e-03 lpdiblc2 = -3.148678279e-10 wpdiblc2 = 1.722146178e-09 ppdiblc2 = 3.155238385e-15
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 1.007386963e+09 lpscbe1 = -8.089663926e+02 wpscbe1 = -2.088591572e+03 ppscbe1 = 8.179431173e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.591643886e-01 lkt1 = -2.013680148e-07 wkt1 = -3.635353044e-07 pkt1 = 1.297352323e-12
+ kt2 = -3.207210312e-02 lkt2 = -1.013769025e-07 wkt2 = -8.518346428e-08 pkt2 = 6.498772853e-13
+ at = 140000.0
+ ute = -1.114228663e+00 lute = -4.156417360e-06 wute = -4.632564872e-06 pute = 2.698548215e-11
+ ua1 = 1.929252841e-09 lua1 = -1.001719677e-14 wua1 = -9.538527051e-15 pua1 = 5.946359680e-20
+ ub1 = -2.202620758e-18 lub1 = 9.598820989e-24 wub1 = 9.184760274e-24 pub1 = -5.316790736e-29
+ uc1 = -2.787028429e-11 luc1 = 3.235987106e-16 wuc1 = 2.060348802e-16 puc1 = -1.470582503e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.12 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.096268598e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.271132523e-08 wvth0 = 6.389719598e-08 pvth0 = -2.450060636e-13
+ k1 = 5.755396052e-01 lk1 = -1.030399791e-07 wk1 = -1.783337836e-07 pk1 = 7.199385416e-13
+ k2 = -4.478792741e-02 lk2 = 4.254912964e-08 wk2 = 8.710150814e-08 pk2 = -3.210030769e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.527821500e-01 ldsub = -1.157040216e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-8.868120019e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -3.954197852e-08 wvoff = -8.920233687e-08 pvoff = 2.703372911e-13
+ nfactor = 2.856287491e+00 lnfactor = -6.148432801e-07 wnfactor = -2.165712561e-06 pnfactor = 6.937930062e-12
+ eta0 = 1.575872698e-01 leta0 = -3.066156572e-7
+ etab = -1.378254975e-01 letab = 2.680382949e-07 wetab = -1.188449825e-11 petab = 4.696612282e-17
+ u0 = 3.427618503e-02 lu0 = -8.073277361e-09 wu0 = -4.894781303e-09 pu0 = 8.945151329e-15
+ ua = -4.134632304e-10 lua = -1.585510600e-15 wua = -1.203021463e-15 pua = 6.483714854e-21
+ ub = 1.399537536e-18 lub = 1.675519622e-24 wub = 1.655238993e-24 pub = -8.714045596e-30
+ uc = -2.108046154e-10 luc = 5.686594070e-16 wuc = 1.565857476e-15 puc = -3.141610557e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 6.165625135e-01 la0 = 1.115262147e-06 wa0 = 4.553711154e-06 pa0 = -8.833812744e-12
+ ags = -9.340263153e-02 lags = 1.534302345e-06 wags = 2.351921389e-06 pags = -5.655198080e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 9.885208938e-06 lketa = -7.682809191e-09 wketa = -2.669065219e-08 pketa = 1.041549698e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 8.375421807e-01 lpclm = -3.022836338e-08 wpclm = -1.567866627e-06 ppclm = -5.424187508e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 1.346347235e-03 lpdiblc2 = 5.474212287e-09 wpdiblc2 = 4.476326575e-10 ppdiblc2 = 8.191964150e-15
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 8.053011024e+08 lpscbe1 = -1.034712106e+01 wpscbe1 = -3.721708918e+01 ppscbe1 = 7.264332925e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.047259471e-01 lkt1 = -2.131415747e-08 wkt1 = -1.254403595e-08 pkt1 = -8.972340239e-14
+ kt2 = -5.829284529e-02 lkt2 = 2.244350219e-09 wkt2 = 8.334601966e-08 pkt2 = -1.613118019e-14
+ at = 1.674704694e+05 lat = -1.085600259e-01 wat = -2.115597552e-02 pat = 8.360589768e-8
+ ute = -2.536150174e+00 lute = 1.462847241e-06 wute = 3.847149092e-06 pute = -6.525338356e-12
+ ua1 = -1.728309101e-09 lua1 = 4.437052779e-15 wua1 = 1.129239202e-14 pua1 = -2.285771648e-20
+ ub1 = 1.245897194e-18 lub1 = -4.029311585e-24 wub1 = -1.016968786e-23 pub1 = 2.331856850e-29
+ uc1 = 6.765861793e-11 luc1 = -5.392014302e-17 wuc1 = -3.035269739e-16 puc1 = 5.431453065e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.13 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.338473676e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.543577620e-08 wvth0 = -1.642829613e-07 pvth0 = 2.003744500e-13
+ k1 = 4.352435178e-01 lk1 = 1.708012883e-07 wk1 = 5.793078755e-07 pk1 = -7.588878177e-13
+ k2 = 1.069414574e-02 lk2 = -6.574527479e-08 wk2 = -2.287588897e-07 pk2 = 2.955188323e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.122467418e+00 ldsub = -1.683433766e-06 wdsub = -6.055066352e-06 pdsub = 1.181876897e-11
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.044535435e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -8.756241257e-09 wvoff = 1.428958202e-07 pvoff = -1.826906918e-13
+ nfactor = 2.276853150e+00 lnfactor = 5.161436005e-07 wnfactor = 4.035876418e-06 pnfactor = -5.166833635e-12
+ eta0 = -6.301712752e-03 leta0 = 1.327613389e-08 weta0 = 3.417787209e-08 peta0 = -6.671113916e-14
+ etab = -9.552859247e-04 letab = 8.839294674e-10 wetab = 1.933898733e-09 petab = -3.750971196e-15
+ u0 = 3.416963449e-02 lu0 = -7.865303385e-09 wu0 = -1.562640200e-10 pu0 = -3.038705237e-16
+ ua = -9.685279801e-10 lua = -5.020902616e-16 wua = 3.765108439e-15 pua = -3.213483507e-21
+ ub = 2.160490419e-18 lub = 1.902301466e-25 wub = -4.999447830e-24 pub = 4.275111175e-30
+ uc = 7.459494227e-11 luc = 1.159343294e-17 wuc = 8.785120596e-17 puc = -2.567182011e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.141218848e+04 lvsat = 1.143564361e-01 wvsat = 2.756624983e-01 pvsat = -5.380603929e-7
+ a0 = 1.957627994e+00 la0 = -1.502338083e-06 wa0 = -4.791631013e-06 pa0 = 9.407183070e-12
+ ags = 1.410381489e+00 lags = -1.400905307e-06 wags = -7.316343842e-06 pags = 1.321610513e-11
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 4.991952291e-02 lketa = -1.051004827e-07 wketa = 8.265099420e-08 pketa = -1.092669123e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.094706358e+00 lpclm = -5.321822355e-07 wpclm = -2.640774551e-06 ppclm = 1.551769841e-12
+ pdiblc1 = -1.774724204e-01 lpdiblc1 = 1.107638636e-06 wpdiblc1 = 1.864479510e-06 ppdiblc1 = -3.639242130e-12
+ pdiblc2 = 6.764259455e-03 lpdiblc2 = -5.100907633e-09 wpdiblc2 = -8.349192880e-09 ppdiblc2 = 2.536232078e-14
+ pdiblcb = -4.838830672e-02 lpdiblcb = 4.565119150e-08 wpdiblcb = -1.589087323e-09 ppdiblcb = 3.101709352e-15
+ drout = 8.455643000e-01 ldrout = -5.573875314e-7
+ pscbe1 = 2.301647263e+09 lpscbe1 = -2.931036761e+03 wpscbe1 = -6.940978551e+03 ppscbe1 = 1.354796416e-2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 4.130171153e-07 lalpha0 = -7.476038300e-13 walpha0 = -2.013114642e-11 palpha0 = 3.929360221e-17
+ alpha1 = 8.176360460e-01 lalpha1 = 6.317058690e-8
+ beta0 = 1.188328349e+01 lbeta0 = 3.858315396e-06 wbeta0 = -4.646939632e-06 pbeta0 = 9.070273176e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.586691458e-01 lkt1 = 8.397654703e-08 wkt1 = -9.922140364e-08 pkt1 = 7.946050472e-14
+ kt2 = -8.651182867e-02 lkt2 = 5.732444773e-08 wkt2 = 1.472002157e-07 pkt2 = -1.407669723e-13
+ at = 1.549976129e+05 lat = -8.421449430e-02 wat = 6.342928877e-02 pat = -8.149447255e-8
+ ute = -2.543197859e+00 lute = 1.476603484e-06 wute = 2.812710781e-07 pute = 4.348311882e-13
+ ua1 = -8.170805901e-10 lua1 = 2.658443162e-15 wua1 = -2.343032036e-15 pua1 = 3.757008658e-21
+ ub1 = -3.665462189e-19 lub1 = -8.820139240e-25 wub1 = 4.635419692e-24 pub1 = -5.579239637e-30
+ uc1 = 1.240513015e-11 luc1 = 5.392808997e-17 wuc1 = 3.885713613e-17 puc1 = -1.251477327e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.14 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.464437866e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.445484319e-09 wvth0 = 7.739053809e-09 pvth0 = 3.662996222e-14
+ k1 = 7.126925567e-01 lk1 = -9.329718025e-08 wk1 = -2.849386482e-07 pk1 = 6.377202754e-14
+ k2 = -1.011625105e-01 lk2 = 4.072895104e-08 wk2 = 1.370491506e-07 pk2 = -5.268689088e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -1.675701909e+00 ldsub = 9.800904509e-07 wdsub = 1.273009634e-05 pdsub = -6.062470478e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.073774119e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -5.973066530e-09 wvoff = -6.531637841e-09 pvoff = -4.045353359e-14
+ nfactor = 2.791748920e+00 lnfactor = 2.602410070e-08 wnfactor = -2.000409581e-06 pnfactor = 5.789923176e-13
+ eta0 = -4.282880735e-01 leta0 = 4.149569329e-07 weta0 = -6.835574418e-08 peta0 = 3.088866204e-14
+ etab = 2.316475173e-04 letab = -2.458899243e-10 wetab = -3.820259473e-09 petab = 1.726302671e-15
+ u0 = 2.947163865e-02 lu0 = -3.393370401e-09 wu0 = -7.459563813e-09 pu0 = 6.648001786e-15
+ ua = -1.275739257e-09 lua = -2.096616843e-16 wua = -1.231090814e-16 pua = 4.876368743e-22
+ ub = 2.327649863e-18 lub = 3.111424813e-26 wub = -2.027580489e-25 pub = -2.907666901e-31
+ uc = 8.765824459e-11 luc = -8.412763313e-19 wuc = -3.268521369e-16 puc = 1.380300316e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.886355565e+05 lvsat = -4.482031060e-02 wvsat = -6.583796375e-01 pvsat = 3.510365694e-7
+ a0 = -6.334613824e-01 la0 = 9.640706629e-07 wa0 = 9.692241100e-06 pa0 = -4.379739601e-12
+ ags = -1.246482431e+00 lags = 1.128112978e-06 wags = 1.250363287e-05 pags = -5.650154124e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -7.980152066e-02 lketa = 1.837851394e-08 wketa = -1.390984530e-07 pketa = 1.018121733e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.789834749e-01 lpclm = 2.442888785e-07 wpclm = -1.283137318e-07 ppclm = -8.397938765e-13
+ pdiblc1 = 6.979695736e-01 lpdiblc1 = 2.743220347e-07 wpdiblc1 = -1.793508050e-06 ppdiblc1 = -1.572732738e-13
+ pdiblc2 = -1.380705581e-03 lpdiblc2 = 2.652129830e-09 wpdiblc2 = 4.157499463e-08 ppdiblc2 = -2.215956476e-14
+ pdiblcb = 2.177661343e-02 lpdiblcb = -2.113746285e-08 wpdiblcb = 3.178174645e-09 ppdiblcb = -1.436156737e-15
+ drout = 9.937327017e-01 ldrout = -6.984262178e-07 wdrout = -6.666146524e-06 pdrout = 6.345378220e-12
+ pscbe1 = -1.444498826e+09 lpscbe1 = 6.348485235e+02 wpscbe1 = 1.007232313e+04 ppscbe1 = -2.646674459e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.967580078e-05 lalpha0 = 1.837456023e-11 walpha0 = 1.353518908e-10 palpha0 = -1.087077468e-16
+ alpha1 = 9.147279080e-01 lalpha1 = -2.924931179e-8
+ beta0 = 2.141331387e+00 lbeta0 = 1.313149451e-05 wbeta0 = 8.797773422e-05 pbeta0 = -7.909739400e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.687445832e-01 lkt1 = -1.620935531e-09 wkt1 = -1.938699117e-09 pkt1 = -1.314105334e-14
+ kt2 = -1.802566897e-02 lkt2 = -7.866226457e-09 wkt2 = 2.789738289e-09 pkt2 = -3.305382607e-15
+ at = 7.930253889e+04 lat = -1.216179160e-02 wat = -4.882815952e-02 pat = 2.536125958e-8
+ ute = -6.999961772e-01 lute = -2.779051763e-07 wute = 2.116455136e-06 pute = -1.312045648e-12
+ ua1 = 2.543325005e-09 lua1 = -5.402630759e-16 wua1 = 4.481635161e-15 pua1 = -2.739262378e-21
+ ub1 = -1.236256342e-18 lub1 = -5.415338227e-26 wub1 = -3.328713499e-24 pub1 = 2.001667429e-30
+ uc1 = 1.460582847e-10 luc1 = -7.329380841e-17 wuc1 = -1.916566077e-16 puc1 = 9.427392030e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.15 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.837470629e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.341115750e-08 wvth0 = 1.654183478e-07 pvth0 = -3.462231481e-14
+ k1 = 3.068429378e-01 lk1 = 9.009855138e-08 wk1 = -3.087869038e-07 pk1 = 7.454860112e-14
+ k2 = 3.883422862e-02 lk2 = -2.253291544e-08 wk2 = 6.034565914e-08 pk2 = -1.802604046e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.002933194e-01 ldsub = 4.198765118e-08 wdsub = -9.545076652e-07 pdsub = 1.213420623e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.047052420e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.180569310e-09 wvoff = -1.619537028e-07 pvoff = 2.977874455e-14
+ nfactor = 3.598500438e+00 lnfactor = -3.385315822e-07 wnfactor = -4.565233141e-06 pnfactor = 1.737987353e-12
+ eta0 = 0.49
+ etab = -2.683563039e-04 letab = -1.994769753e-11 wetab = 2.963176190e-09 petab = -1.339003020e-15
+ u0 = 2.389414900e-02 lu0 = -8.730088019e-10 wu0 = 1.979720304e-08 pu0 = -5.668813275e-15
+ ua = -1.387352258e-09 lua = -1.592258898e-16 wua = 1.489461369e-15 pua = -2.410530733e-22
+ ub = 2.080114045e-18 lub = 1.429709812e-25 wub = -6.971384153e-25 pub = -6.736559575e-32
+ uc = 1.190810864e-11 luc = 3.338877085e-17 wuc = 4.869219331e-16 puc = -2.296990089e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.952416086e+04 lvsat = 1.352267595e-02 wvsat = 2.466147287e-01 pvsat = -5.791318977e-8
+ a0 = 1.5
+ ags = 2.243633756e+00 lags = -4.490042151e-07 wags = -3.557951722e-12 pags = 1.607770782e-18
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.698741901e-02 lketa = -5.487175127e-09 wketa = 6.732593279e-08 pketa = 8.532915438e-15
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.175856166e+00 lpclm = -1.609908502e-07 wpclm = -3.781527232e-06 ppclm = 8.110238931e-13
+ pdiblc1 = 3.036609324e+00 lpdiblc1 = -7.824648342e-07 wpdiblc1 = -9.298826698e-06 ppdiblc1 = 3.234237622e-12
+ pdiblc2 = 6.046156329e-03 lpdiblc2 = -7.039279567e-10 wpdiblc2 = -1.337997833e-08 ppdiblc2 = 2.673543383e-15
+ pdiblcb = 5.419328835e-01 lpdiblcb = -2.561861983e-07 wpdiblcb = -2.846361377e-06 ppdiblcb = 1.286216625e-12
+ drout = -1.805033163e+00 ldrout = 5.662829001e-07 wdrout = 1.333229305e-05 pdrout = -2.691536653e-12
+ pscbe1 = -7.175914011e+08 lpscbe1 = 3.063728696e+02 wpscbe1 = 7.619267951e+03 ppscbe1 = -1.538185433e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.957237663e-05 lalpha0 = -8.398565421e-12 walpha0 = -2.166503568e-10 palpha0 = 5.035538088e-17
+ alpha1 = 0.85
+ beta0 = 4.151249225e+01 lbeta0 = -4.659585035e-06 wbeta0 = -1.613099204e-04 pbeta0 = 3.355096067e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.200317414e-01 lkt1 = -2.363334316e-08 wkt1 = -3.136567626e-07 pkt1 = 1.277184169e-13
+ kt2 = -4.388916277e-03 lkt2 = -1.402841590e-08 wkt2 = -2.005181813e-07 pkt2 = 8.856560340e-14
+ at = 7.631558333e+04 lat = -1.081204314e-02 wat = -4.758443768e-03 pat = 5.446992356e-9
+ ute = -1.215157672e+00 lute = -4.511348475e-08 wute = -4.652650750e-06 pute = 1.746784689e-12
+ ua1 = 1.714603108e-09 lua1 = -1.657793964e-16 wua1 = -6.071213526e-15 pua1 = 2.029369440e-21
+ ub1 = -2.029427825e-18 lub1 = 3.042657406e-25 wub1 = 3.379107700e-24 pub1 = -1.029469523e-30
+ uc1 = -1.233366081e-10 luc1 = 4.844062513e-17 wuc1 = 1.811671720e-16 puc1 = -7.419806207e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.16 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.933526007e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.535033307e-08 wvth0 = 5.095759264e-07 pvth0 = -1.041011909e-13
+ k1 = 5.036432250e-01 lk1 = 5.036831260e-08 wk1 = 1.590637675e-07 pk1 = -1.990156026e-14
+ k2 = -9.014653428e-03 lk2 = -1.287313529e-08 wk2 = -1.679965932e-07 pk2 = 2.807192179e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 9.851946489e-01 ldsub = -7.609281412e-08 wdsub = -8.967115455e-07 pdsub = 1.096741239e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-7.249742839e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.368271493e-08 wvoff = -3.245631871e-07 pvoff = 6.260650986e-14
+ nfactor = 6.197083821e-01 lnfactor = 2.628299369e-07 wnfactor = 5.034699331e-06 pnfactor = -2.000566145e-13
+ eta0 = 1.386034242e+00 leta0 = -1.808922888e-07 weta0 = -2.193190777e-07 peta0 = 4.427635473e-14
+ etab = 6.731936023e-02 letab = -1.366462350e-08 wetab = -1.155573934e-07 petab = 2.258804808e-14
+ u0 = -1.873414963e-03 lu0 = 4.328972778e-09 wu0 = 2.544004910e-08 pu0 = -6.807996681e-15
+ ua = -4.766767181e-09 lua = 5.230137743e-16 wua = 5.252958532e-17 pua = 4.903615210e-23
+ ub = 4.373588145e-18 lub = -3.200378636e-25 wub = 2.212858690e-24 pub = -6.548387214e-31
+ uc = 3.246411690e-10 luc = -2.974609210e-17 wuc = -1.709279004e-15 puc = 2.136722325e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.104885540e+04 lvsat = 1.321486910e-02 wvsat = 2.889300084e-01 pvsat = -6.645584076e-8
+ a0 = 1.5
+ ags = -2.298691984e+00 lags = 4.680050476e-07 wags = 1.270697043e-11 pags = -1.675807967e-18
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.048909338e-01 lketa = 1.024006434e-08 wketa = 4.747822755e-07 pketa = -7.372477848e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.057117069e+00 lpclm = -1.370196824e-07 wpclm = -2.868421266e-06 ppclm = 6.266851476e-13
+ pdiblc1 = -3.124198466e+00 lpdiblc1 = 4.612852032e-07 wpdiblc1 = 1.936779339e-05 ppdiblc1 = -2.553008308e-12
+ pdiblc2 = -7.063513872e-03 lpdiblc2 = 1.942665373e-09 wpdiblc2 = -1.577192467e-08 ppdiblc2 = 3.156431900e-15
+ pdiblcb = -2.027975080e+00 lpdiblcb = 2.626293912e-07 wpdiblcb = 1.082418594e-05 ppdiblcb = -1.473607137e-12
+ drout = 1.940375001e+00 ldrout = -1.898438455e-07 wdrout = -2.857490781e-06 pdrout = 5.768730964e-13
+ pscbe1 = 8.157026898e+08 lpscbe1 = -3.170074713e+00 wpscbe1 = -5.596579857e+01 ppscbe1 = 1.129843138e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.240360062e-06 lalpha0 = -8.619405840e-13 walpha0 = 3.759527756e-11 palpha0 = -9.719820277e-19
+ alpha1 = -2.250685343e+00 lalpha1 = 6.259694576e-07 walpha1 = 1.725705094e-05 palpha1 = -3.483870700e-12
+ beta0 = 4.093927223e+01 lbeta0 = -4.543862804e-06 wbeta0 = -9.854822717e-05 pbeta0 = 2.088056728e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.487777652e-01 lkt1 = 4.273423286e-08 wkt1 = 1.374795228e-06 pkt1 = -2.131479593e-13
+ kt2 = -1.438741777e-01 lkt2 = 1.413100817e-08 wkt2 = 6.794727969e-07 pkt2 = -8.908785527e-14
+ at = 3.640858180e+04 lat = -2.755577762e-03 wat = -2.064308906e-01 pat = 4.616082760e-8
+ ute = -7.557782616e-01 lute = -1.378534596e-07 wute = 1.184508971e-05 pute = -1.583795653e-12
+ ua1 = 3.687410867e-09 lua1 = -5.640517997e-16 wua1 = 1.102394017e-14 pua1 = -1.421817283e-21
+ ub1 = -3.872944109e-18 lub1 = 6.764366515e-25 wub1 = -4.751703146e-25 pub1 = -2.513640227e-31
+ uc1 = -6.615015636e-11 luc1 = 3.689576707e-17 wuc1 = 5.469079661e-16 puc1 = -1.480341793e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.17 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.840807109e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -9.394469691e-10 wvth0 = 8.627281753e-07 pvth0 = -1.506752627e-13
+ k1 = 8.182619762e-01 lk1 = 8.876077074e-09 wk1 = 9.914489443e-08 pk1 = -1.199939936e-14
+ k2 = -5.194733661e-02 lk2 = -7.211130095e-09 wk2 = -4.367371876e-07 pk2 = 6.351370011e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.248986900e+00 ldsub = -1.108820000e-07 wdsub = -4.241399208e-06 pdsub = 5.507748774e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 5.320138903e-02 lcdscd = -6.304094285e-09 wcdscd = -2.068475025e-07 pcdscd = 2.727925548e-14
+ cit = 0.0
+ voff = {4.187749292e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.847220473e-08 wvoff = -2.525214822e-06 pvoff = 3.528306481e-13
+ nfactor = 1.899302995e+01 lnfactor = -2.160262085e-06 wnfactor = -8.302392790e-05 pnfactor = 1.141320320e-11
+ eta0 = 6.007280197e-02 leta0 = -6.023168140e-09 weta0 = 5.158301557e-07 peta0 = -5.267586132e-14
+ etab = 2.138091657e-02 letab = -7.606215610e-09 wetab = -9.907789327e-09 petab = 8.654872652e-15
+ u0 = 5.074416411e-02 lu0 = -2.610286167e-09 wu0 = 1.157985984e-07 pu0 = -1.872457252e-14
+ ua = 4.832378658e-09 lua = -7.429311781e-16 wua = 2.467647860e-16 pua = 2.342021960e-23
+ ub = -4.579732589e-18 lub = 8.607350280e-25 wub = 1.054222310e-23 pub = -1.753323629e-30
+ uc = 1.575002746e-10 luc = -7.703383806e-18 wuc = 2.940812895e-16 puc = -5.053292638e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.753359793e+05 lvsat = -1.857431086e-03 wvsat = -6.456705011e-01 pvsat = 5.680020903e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.912013126e-01 lketa = 1.139394634e-07 wketa = 4.509016728e-06 pketa = -6.057636523e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.174476039e-01 lpclm = 9.701168114e-08 wpclm = 9.835973826e-06 ppclm = -1.048783182e-12
+ pdiblc1 = -3.636638727e-02 lpdiblc1 = 5.405882083e-08 wpdiblc1 = 2.604985400e-06 ppdiblc1 = -3.423124271e-13
+ pdiblc2 = -4.237141443e-03 lpdiblc2 = 1.569920551e-09 wpdiblc2 = 7.451250516e-08 ppdiblc2 = -8.750368990e-15
+ pdiblcb = -4.660076154e-01 lpdiblcb = 5.663556003e-08 wpdiblcb = 6.066935773e-07 ppdiblcb = -1.261140269e-13
+ drout = -1.226762679e-01 ldrout = 8.223341884e-08 wdrout = 1.019355747e-05 pdrout = -1.144312198e-12
+ pscbe1 = 8.099648223e+08 lpscbe1 = -2.413359009e+00 wpscbe1 = 2.904784237e+01 ppscbe1 = 8.674740096e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.898453629e-05 lalpha0 = 1.937219971e-12 walpha0 = 1.328706924e-10 palpha0 = -1.353699901e-17
+ alpha1 = 8.084932466e+00 lalpha1 = -7.371021546e-07 walpha1 = -4.026645218e-05 palpha1 = 4.102386415e-12
+ beta0 = -1.856071010e+01 lbeta0 = 3.303054366e-06 wbeta0 = 2.627976176e-04 pbeta0 = -2.677408408e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.697073507e-01 lkt1 = 3.230634752e-08 wkt1 = 4.362842009e-07 pkt1 = -8.937618662e-14
+ kt2 = -5.934352408e-02 lkt2 = 2.983021033e-09 wkt2 = 2.354660740e-09 pkt2 = 2.111616443e-16
+ at = 1.793791159e+05 lat = -2.161067476e-02 wat = -9.296598824e-01 pat = 1.415409903e-7
+ ute = -7.917541749e+00 lute = 8.066470710e-07 wute = -7.217792350e-07 pute = 7.353559025e-14
+ ua1 = -1.080475665e-08 lua1 = 1.347189745e-15 wua1 = 1.137741903e-14 pua1 = -1.468434429e-21
+ ub1 = 6.739153551e-18 lub1 = -7.230974000e-25 wub1 = -6.156191259e-24 pub1 = 4.978547005e-31
+ uc1 = 2.405016708e-10 luc1 = -3.545782549e-18 wuc1 = -1.412332007e-15 puc1 = 1.103523475e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.18 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.242783392e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.782644595e-07 wvth0 = -7.349098088e-09 pvth0 = 7.345561776e-13
+ k1 = 5.438963270e-01 lk1 = -3.029218688e-07 wk1 = -1.714130182e-08 pk1 = 1.713305360e-12
+ k2 = -2.827807665e-02 lk2 = 1.551838561e-07 wk2 = 5.591961849e-09 pk2 = -5.589271053e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.061930727e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 9.240278277e-08 wvoff = 3.153846883e-09 pvoff = -3.152329284e-13
+ nfactor = 2.489367473e+00 lnfactor = 8.898968531e-06 wnfactor = -4.784544444e-08 pnfactor = 4.782242169e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.202281576e-02 lu0 = -3.230020667e-09 wu0 = 1.150370903e-09 pu0 = -1.149817356e-13
+ ua = -7.600960480e-10 lua = 2.576337686e-16 wua = -3.592368347e-17 pua = 3.590639735e-21
+ ub = 1.751104992e-18 lub = -1.621218738e-24 wub = 6.664700209e-26 pub = -6.661493222e-30
+ uc = 5.896655521e-11 luc = -9.719875851e-16 wuc = -4.574440536e-17 puc = 4.572239361e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.328513376e+00 la0 = -1.401263024e-06 wa0 = -1.184702374e-07 pa0 = 1.184132307e-11
+ ags = 4.331596951e-01 lags = -9.597074838e-07 wags = -3.254984210e-08 pags = 3.253417944e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 7.937578791e-25 lb0 = -7.933759308e-29 wb0 = -3.985166208e-30 pb0 = 3.983248586e-34
+ b1 = 2.632910460e-24 lb1 = -5.253151618e-29
+ keta = -9.245665968e-03 lketa = 4.508489201e-08 wketa = -1.000500816e-09 pketa = 1.000019385e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.620939740e-02 lpclm = 1.010173941e-06 wpclm = -1.257408538e-08 ppclm = 1.256803485e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 2.768070182e-03 lpdiblc2 = 3.052415685e-08 wpdiblc2 = 1.382698548e-09 ppdiblc2 = -1.382033207e-13
+ pdiblcb = -9.616352767e-01 lpdiblcb = 9.361845772e-05 wpdiblcb = 4.702501042e-06 ppdiblcb = -4.700238246e-10
+ drout = 0.56
+ pscbe1 = 8.069588658e+08 lpscbe1 = -5.225954690e+03 wpscbe1 = -1.871938452e+02 ppscbe1 = 1.871037694e-2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.071583742e-01 lkt1 = -5.868800464e-07 wkt1 = -1.524246175e-08 pkt1 = 1.523512723e-12
+ kt2 = -4.358904271e-02 lkt2 = -1.723464573e-07 wkt2 = -8.411420136e-09 pkt2 = 8.407372645e-13
+ at = 140000.0
+ ute = -1.760686254e+00 lute = -5.268838076e-06 wute = -1.766310083e-07 pute = 1.765460152e-11
+ ua1 = 4.322170872e-10 lua1 = -5.617004568e-15 wua1 = -1.357449013e-16 pua1 = 1.356795822e-20
+ ub1 = -6.475970438e-19 lub1 = 7.973205360e-25 wub1 = -1.374658244e-25 pub1 = 1.373996772e-29
+ uc1 = 1.483067491e-11 luc1 = 9.985573607e-17 wuc1 = 3.516725267e-18 puc1 = -3.515033054e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.19 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.103315610e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = 2.946728918e-8
+ k1 = 5.287137050e-01 wk1 = 6.873056959e-8
+ k2 = -2.050017059e-02 wk2 = -2.242179311e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.015617909e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = -1.264581273e-8
+ nfactor = 2.935389005e+00 wnfactor = 1.918433432e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.186092522e-02 wu0 = -4.612581253e-9
+ ua = -7.471832921e-10 wua = 1.440412900e-16
+ ub = 1.669848556e-18 wub = -2.672309527e-25
+ uc = 1.024996628e-11 wuc = 1.834189182e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.258281250e+00 wa0 = 4.750238330e-7
+ ags = 3.850585920e-01 wags = 1.305133771e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -3.182688907e-24 wb0 = 1.597910977e-29
+ b1 = 0.0
+ keta = -6.985984688e-03 wketa = 4.011655107e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.683990892e-02 wpclm = 5.041764384e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 4.297958860e-03 wpdiblc2 = -5.544133097e-9
+ pdiblcb = 3.730576837e+00 wpdiblcb = -1.885536925e-5
+ drout = 0.56
+ pscbe1 = 5.450309458e+08 wpscbe1 = 7.505812417e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.365731470e-01 wkt1 = 6.111689117e-8
+ kt2 = -5.222714843e-02 wkt2 = 3.372682560e-8
+ at = 140000.0
+ ute = -2.024763514e+00 wute = 7.082279944e-7
+ ua1 = 1.506895175e-10 wua1 = 5.442891375e-16
+ ub1 = -6.076348700e-19 wub1 = 5.511894316e-25
+ uc1 = 1.983550308e-11 wuc1 = -1.410082695e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.20 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.900072432e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.616165564e-07 wvth0 = 8.352686370e-08 pvth0 = -4.298753035e-13
+ k1 = 5.140076064e-01 lk1 = 1.169411458e-07 wk1 = 1.037360563e-07 pk1 = -2.783594647e-13
+ k2 = -6.745359820e-03 lk2 = -1.093766184e-07 wk2 = -5.236752809e-08 pk2 = 2.381249211e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.016172852e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 4.412838967e-10 wvoff = -1.857527776e-08 pvoff = 4.715040035e-14
+ nfactor = 4.219757848e+00 lnfactor = -1.021314820e-05 wnfactor = -4.497699826e-06 pnfactor = 3.729068922e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.916724017e-02 lu0 = 2.141986303e-08 wu0 = 5.106919861e-09 pu0 = -7.728831624e-14
+ ua = -6.537445677e-10 lua = -7.430136177e-16 wua = -2.804145827e-16 pua = 3.375222589e-21
+ ub = 1.289097530e-18 lub = 3.027686853e-24 wub = 1.161312464e-24 pub = -1.135960725e-29
+ uc = -1.039980703e-10 luc = 9.084867911e-16 wuc = 5.593360188e-16 puc = -2.989248050e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.028273433e+00 la0 = 1.828994790e-06 wa0 = 1.591885458e-06 pa0 = -8.881150736e-12
+ ags = 2.276293407e-01 lags = 1.251858672e-06 wags = 5.875104751e-07 pags = -3.633986541e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -6.327090862e-24 lb0 = 2.500391016e-29 wb0 = 3.176599485e-29 pb0 = -1.255354315e-34
+ b1 = 0.0
+ keta = -9.949582930e-03 lketa = 2.356618055e-08 wketa = -1.873004631e-09 pketa = 4.679411396e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.536152732e-01 lpclm = 3.343409574e-06 wpclm = 1.108667378e-07 ppclm = -4.806840016e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 5.733887536e-03 lpdiblc2 = -1.141833396e-08 wpdiblc2 = -1.295139381e-08 ppdiblc2 = 5.890165575e-14
+ pdiblcb = 7.440975023e+00 lpdiblcb = -2.950464484e-05 wpdiblcb = -3.748391311e-05 ppdiblcb = 1.481319640e-10
+ drout = 0.56
+ pscbe1 = 2.957796568e+08 lpscbe1 = 1.982016589e+03 wpscbe1 = 1.484126839e+03 ppscbe1 = -5.833067298e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.578913672e-01 lkt1 = 1.695199501e-07 wkt1 = 1.321365232e-07 pkt1 = -5.647396623e-13
+ kt2 = -6.272827337e-02 lkt2 = 8.350369592e-08 wkt2 = 6.872988506e-08 pkt2 = -2.783401635e-13
+ at = 140000.0
+ ute = -2.368694122e+00 lute = 2.734895264e-06 wute = 1.665644552e-06 pute = -7.613262537e-12
+ ua1 = -4.919840822e-10 lua1 = 5.110463987e-15 wua1 = 2.617612526e-15 pua1 = -1.648682086e-20
+ ub1 = -1.837194745e-19 lub1 = -3.370924780e-24 wub1 = -9.514001169e-25 pub1 = 1.194841328e-29
+ uc1 = 2.802841252e-11 luc1 = -6.514904086e-17 wuc1 = -7.461190576e-17 puc1 = 4.811768978e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.21 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.370774918e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.439946480e-08 wvth0 = -7.392232566e-08 pvth0 = 1.923451564e-13
+ k1 = 5.393751731e-01 lk1 = 1.669154093e-08 wk1 = 3.234521560e-09 pk1 = 1.188106409e-13
+ k2 = -3.353326717e-02 lk2 = -3.513996358e-09 wk2 = 3.059600080e-08 pk2 = -8.973707248e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.294975716e+00 ldsub = -2.904536566e-06 wdsub = -2.220091166e-06 pdsub = 8.773536097e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.064943691e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.971493928e-08 wvoff = 2.310291441e-10 pvoff = -2.716988659e-14
+ nfactor = 5.601714499e-01 lnfactor = 4.249101755e-06 wnfactor = 9.362241111e-06 pnfactor = -1.748214803e-11
+ eta0 = 2.747685646e-01 leta0 = -7.697021900e-07 weta0 = -5.883241590e-07 peta0 = 2.324987066e-12
+ etab = -2.402693739e-01 letab = 6.728843034e-07 wetab = 5.143211193e-07 petab = -2.032535859e-12
+ u0 = 3.851999148e-02 lu0 = -1.554109720e-08 wu0 = -2.620137176e-08 pu0 = 4.643832656e-14
+ ua = -8.605867453e-10 lua = 7.440205406e-17 wua = 1.041821164e-15 pua = -1.850095736e-21
+ ub = 2.416343257e-18 lub = -1.427054118e-24 wub = -3.449768350e-24 pub = 6.862835406e-30
+ uc = 1.672537765e-10 luc = -1.634682285e-16 wuc = -3.322345846e-16 puc = 5.341328776e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 2.269020746e+00 la0 = -3.074290942e-06 wa0 = -3.742673527e-06 pa0 = 1.220039156e-11
+ ags = 6.299887533e-01 lags = -3.382178455e-07 wags = -1.279960546e-06 pags = 3.746036707e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.106115003e-24 lb0 = -1.227499686e-29 wb0 = -1.559466038e-29 pb0 = 6.162824206e-35
+ b1 = 0.0
+ keta = -1.069866621e-02 lketa = 2.652646854e-08 wketa = 2.707304374e-08 pketa = -6.759722463e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.026634605e-01 lpclm = -4.356901846e-07 wpclm = -3.886270084e-07 ppclm = 1.493255844e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 3.319665137e-04 lpdiblc2 = 9.929415094e-09 wpdiblc2 = 5.540464969e-09 ppdiblc2 = -1.417596963e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 7.824079358e+08 lpscbe1 = 5.891953937e+01 wpscbe1 = 7.772107556e+01 ppscbe1 = -2.751190827e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.953515374e-01 lkt1 = -7.763001502e-08 wkt1 = -5.960949764e-08 pkt1 = 1.930177941e-13
+ kt2 = -4.017600980e-02 lkt2 = -5.620165998e-09 wkt2 = -7.611944328e-09 pkt2 = 2.335366159e-14
+ at = 1.616795051e+05 lat = -8.567482415e-02 wat = 7.918325159e-03 pat = -3.129227875e-8
+ ute = -1.518792910e+00 lute = -6.238131861e-07 wute = -1.260627340e-06 pute = 3.951015756e-12
+ ua1 = 1.258548293e-09 lua1 = -1.807431647e-15 wua1 = -3.703519794e-15 pua1 = 8.493541853e-21
+ ub1 = -1.511586973e-18 lub1 = 1.876649558e-24 wub1 = 3.674625385e-24 pub1 = -6.333089004e-30
+ uc1 = 3.187787385e-12 luc1 = 3.301815362e-17 wuc1 = 2.015734097e-17 puc1 = 1.066601123e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.22 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.058189185e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.661355049e-08 wvth0 = -2.356243299e-08 pvth0 = 9.404863871e-14
+ k1 = 4.326648764e-01 lk1 = 2.249773415e-07 wk1 = 5.922542850e-07 pk1 = -1.030885844e-12
+ k2 = 5.188525143e-03 lk2 = -7.909432706e-08 wk2 = -2.011171947e-07 pk2 = 3.625395113e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -1.486854549e+00 ldsub = 2.525265073e-06 wdsub = 7.045379013e-06 pdsub = -9.311559101e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-8.555778923e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.115077323e-08 wvoff = 4.802719159e-08 pvoff = -1.204623079e-13
+ nfactor = 2.570217394e+00 lnfactor = 3.257312671e-07 wnfactor = 2.563002507e-06 pnfactor = -4.210843381e-12
+ eta0 = -2.309278936e-01 leta0 = 2.173571186e-07 weta0 = 1.161943264e-06 peta0 = -1.091326662e-12
+ etab = 8.362490895e-02 letab = 4.068120681e-08 wetab = -4.227121342e-07 petab = -2.035584553e-13
+ u0 = 3.449825574e-02 lu0 = -7.691147623e-09 wu0 = -1.806150391e-09 pu0 = -1.178242518e-15
+ ua = -3.398391863e-10 lua = -9.420352121e-16 wua = 6.086933631e-16 pua = -1.004681810e-21
+ ub = 1.234660257e-18 lub = 8.794504773e-25 wub = -3.511952922e-25 pub = 8.147895277e-31
+ uc = 1.498308902e-10 luc = -1.294608276e-16 wuc = -2.898808016e-16 puc = 4.514633333e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.441014302e+04 lvsat = 3.042954562e-02 wvsat = 5.978559181e-02 pvsat = -1.166943607e-7
+ a0 = -6.008028347e-01 la0 = 2.527263178e-06 wa0 = 8.053308673e-06 pa0 = -1.082396197e-11
+ ags = -5.928539822e-01 lags = 2.048625656e-06 wags = 2.741164266e-06 pags = -4.102720413e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -6.212230006e-24 lb0 = 5.913303710e-30 wb0 = 3.118932076e-29 pb0 = -2.968852183e-35
+ b1 = 0.0
+ keta = 9.171951258e-02 lketa = -1.733816287e-07 wketa = -1.272113715e-07 pketa = 2.335475941e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.220103576e+00 lpclm = -1.640859814e-06 wpclm = -3.270347834e-06 ppclm = 7.118031971e-12
+ pdiblc1 = 2.291815534e-01 lpdiblc1 = 3.138984703e-07 wpdiblc1 = -1.771804442e-07 ppdiblc1 = 3.458351426e-13
+ pdiblc2 = 3.226925169e-03 lpdiblc2 = 4.278800299e-09 wpdiblc2 = 9.410460830e-09 ppdiblc2 = -2.172974102e-14
+ pdiblcb = -4.884111431e-02 lpdiblcb = 4.653501805e-08 wpdiblcb = 6.842929999e-10 ppdiblcb = -1.335658505e-15
+ drout = 8.455643000e-01 ldrout = -5.573875314e-07 pdrout = -8.881784197e-28
+ pscbe1 = 5.769753976e+08 lpscbe1 = 4.598994075e+02 wpscbe1 = 1.717964206e+03 ppscbe1 = -3.476678484e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -9.032675154e-06 lalpha0 = 1.768926344e-11 walpha0 = 2.729219845e-11 palpha0 = -5.327112360e-17
+ alpha1 = 1.086474933e+00 lalpha1 = -4.615709278e-07 walpha1 = -1.349741117e-06 palpha1 = 2.634534040e-12
+ beta0 = 7.536129003e+00 lbeta0 = 1.234344365e-05 wbeta0 = 1.717852330e-05 pbeta0 = -3.353043324e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.669142542e-01 lkt1 = 6.205189237e-08 wkt1 = -5.782574820e-08 pkt1 = 1.895361275e-13
+ kt2 = -7.240722758e-02 lkt2 = 5.729133559e-08 wkt2 = 7.638620412e-08 pkt2 = -1.406007284e-13
+ at = 1.758501549e+05 lat = -1.133342462e-01 wat = -4.126365090e-02 pat = 6.470508586e-8
+ ute = -3.256385789e+00 lute = 2.767761340e-06 wute = 3.861925222e-06 pute = -6.047597262e-12
+ ua1 = -2.485904305e-09 lua1 = 5.501294235e-15 wua1 = 6.035517711e-15 pua1 = -1.051590041e-20
+ ub1 = 5.163814222e-19 lub1 = -2.081703421e-24 wub1 = 2.025649231e-25 pub1 = 4.439598422e-31
+ uc1 = -1.035408583e-10 luc1 = 2.413397694e-16 wuc1 = 6.209792762e-16 puc1 = -1.066072807e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.23 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.120355648e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.069604305e-08 wvth0 = 1.804900732e-07 pvth0 = -1.001850650e-13
+ k1 = 9.779785293e-01 lk1 = -2.940963637e-07 wk1 = -1.616841891e-06 pk1 = 1.071910834e-12
+ k2 = -1.867046085e-01 lk2 = 1.035651009e-07 wk2 = 5.665245449e-07 pk2 = -3.681640754e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.861196590e+00 ldsub = -6.616811938e-07 wdsub = -5.027369449e-06 pdsub = 2.180260778e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-7.849352461e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.787511250e-08 wvoff = -1.515470065e-07 pvoff = 6.950857927e-14
+ nfactor = 3.162673733e+00 lnfactor = -2.382166651e-07 wnfactor = -3.862686568e-06 pnfactor = 1.905647962e-12
+ eta0 = -4.477608914e-01 leta0 = 4.237563294e-07 weta0 = 2.941010842e-08 peta0 = -1.328986920e-14
+ etab = 2.404202112e-01 letab = -1.085692623e-07 wetab = -1.209718648e-06 petab = 5.455780924e-13
+ u0 = 2.765063597e-02 lu0 = -1.173028469e-09 wu0 = 1.683020473e-09 pu0 = -4.499517970e-15
+ ua = -1.188075671e-09 lua = -1.346150188e-16 wua = -5.632356850e-16 pua = 1.108551838e-22
+ ub = 2.125890712e-18 lub = 3.110514034e-26 wub = 8.102003979e-25 pub = -2.907209632e-31
+ uc = -5.518879117e-11 luc = 6.569351167e-17 wuc = 3.903302619e-16 puc = -1.960166541e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.350679447e+04 lvsat = 1.225180595e-02 wvsat = -1.305668109e-01 pvsat = 6.449847474e-8
+ a0 = 2.555097751e+00 la0 = -4.767786267e-07 wa0 = -6.316340918e-06 pa0 = 2.854234450e-12
+ ags = 1.749354146e+00 lags = -1.808777591e-07 wags = -2.537360118e-06 pags = 9.218066563e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.708802463e-01 lketa = 7.658209239e-08 wketa = 3.181743114e-07 pketa = -1.904065752e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.374592147e+00 lpclm = 8.289817453e-07 wpclm = 8.173680951e-06 ppclm = -3.775321594e-12
+ pdiblc1 = -2.464605840e-01 lpdiblc1 = 7.666531837e-07 wpdiblc1 = 2.948128221e-06 ppdiblc1 = -2.629086795e-12
+ pdiblc2 = 9.383319755e-03 lpdiblc2 = -1.581354736e-09 wpdiblc2 = -1.246721542e-08 ppdiblc2 = -9.047966717e-16
+ pdiblcb = 2.268222863e-02 lpdiblcb = -2.154669316e-08 wpdiblcb = -1.368586000e-09 ppdiblcb = 6.184380102e-16
+ drout = -2.210973268e-01 ldrout = 4.579474045e-07 wdrout = -5.669320086e-07 pdrout = 5.396518073e-13
+ pscbe1 = 1.295213052e+09 lpscbe1 = -2.237773691e+02 wpscbe1 = -3.682761996e+03 ppscbe1 = 1.664170174e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.253689184e-05 lalpha0 = -1.236120756e-11 walpha0 = -7.658250451e-11 palpha0 = 4.560523253e-17
+ alpha1 = 3.770501350e-01 lalpha1 = 2.137170580e-07 walpha1 = 2.699482233e-06 palpha1 = -1.219844731e-12
+ beta0 = 3.218327149e+01 lbeta0 = -1.111770299e-05 wbeta0 = -6.285179161e-05 pbeta0 = 4.264890295e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.236262667e-01 lkt1 = 2.084687954e-08 wkt1 = 2.736020376e-07 pkt1 = -1.259436847e-13
+ kt2 = 8.771857069e-03 lkt2 = -1.998149268e-08 wkt2 = -1.317507784e-07 pkt2 = 5.752091070e-14
+ at = 4.955415599e+04 lat = 6.884515460e-03 wat = 1.005275236e-01 pat = -7.026323915e-8
+ ute = 9.647843608e-01 lute = -1.250290323e-06 wute = -6.241795306e-06 pute = 3.569942338e-12
+ ua1 = 5.348312815e-09 lua1 = -1.955948191e-15 wua1 = -9.601176399e-15 pua1 = 4.368371615e-21
+ ub1 = -1.391645313e-18 lub1 = -2.654890240e-25 wub1 = -2.548562657e-24 pub1 = 3.062705915e-30
+ uc1 = 3.855317782e-10 luc1 = -2.241991810e-16 wuc1 = -1.393964893e-15 puc1 = 8.519142630e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.24 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {6.272563756e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.137005217e-08 wvth0 = -5.302589977e-08 pvth0 = 5.336366430e-15
+ k1 = -9.842068180e-03 lk1 = 1.522809957e-07 wk1 = 1.281171971e-06 pk1 = -2.376465687e-13
+ k2 = 1.359112136e-01 lk2 = -4.221885943e-08 wk2 = -4.270421580e-07 pk2 = 8.080983986e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 3.265054909e-01 ldsub = 3.181655489e-08 wdsub = -5.840461320e-07 pdsub = 1.724073938e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.400973809e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -3.750030739e-11 wvoff = 1.573720230e-08 pvoff = -6.083976262e-15
+ nfactor = 2.793853105e+00 lnfactor = -7.155363080e-08 wnfactor = -5.253949915e-07 pnfactor = 3.975893069e-13
+ eta0 = 0.49
+ etab = 1.751876472e-03 letab = -7.195765343e-10 wetab = -7.179669130e-09 petab = 2.173575906e-15
+ u0 = 3.021057267e-02 lu0 = -2.329815222e-09 wu0 = -1.191523576e-08 pu0 = 1.645275657e-15
+ ua = -9.455415431e-10 lua = -2.442115831e-16 wua = -7.287076436e-16 pua = 1.856288179e-22
+ ub = 1.827956372e-18 lub = 1.657360080e-25 wub = 5.688524647e-25 pub = -1.816604178e-31
+ uc = 1.571656521e-10 luc = -3.026542653e-17 wuc = -2.423627380e-16 puc = 8.988529140e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.183300764e+05 lvsat = -3.484173490e-03 wvsat = -4.862813243e-02 pvsat = 2.747194277e-8
+ a0 = 1.5
+ ags = 2.422716309e+00 lags = -4.851573266e-07 wags = -8.991111543e-07 pags = 1.815130762e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.432787832e-02 lketa = -7.109940171e-09 wketa = -1.401029711e-07 pketa = 1.668022154e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.609333087e-01 lpclm = 4.473076669e-08 wpclm = 3.099005450e-07 ppclm = -2.218286399e-13
+ pdiblc1 = 1.798001305e+00 lpdiblc1 = -1.572002990e-07 wpdiblc1 = -3.080231643e-06 ppdiblc1 = 9.501448864e-14
+ pdiblc2 = 8.650677437e-03 lpdiblc2 = -1.250287593e-09 wpdiblc2 = -2.645632035e-08 ppdiblc2 = 5.416614054e-15
+ pdiblcb = -2.689232835e-01 lpdiblcb = 1.102242973e-07 wpdiblcb = 1.224649043e-06 ppdiblcb = -5.533956341e-13
+ drout = 6.246268936e-01 ldrout = 7.578069809e-08 wdrout = 1.133864017e-06 pdrout = -2.289056016e-13
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.380625504e-05 lalpha0 = 4.061569999e-12 walpha0 = 5.134410949e-11 palpha0 = -1.220237373e-17
+ alpha1 = 0.85
+ beta0 = -2.305805796e+00 lbeta0 = 4.467255741e-06 wbeta0 = 5.868562893e-05 pbeta0 = -1.227154819e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.474428469e-01 lkt1 = -1.357896042e-08 wkt1 = -1.760356897e-07 pkt1 = 7.723906117e-14
+ kt2 = -3.134935994e-02 lkt2 = -1.851477022e-09 wkt2 = -6.515971511e-08 pkt2 = 2.742967441e-14
+ at = 8.967589036e+04 lat = -1.124573399e-02 wat = -7.183562875e-02 pat = 7.624394514e-9
+ ute = -2.298161102e+00 lute = 2.241727353e-07 wute = 7.847109267e-07 pute = 3.947976750e-13
+ ua1 = 1.337735152e-09 lua1 = -1.436443466e-16 wua1 = -4.179098209e-15 pua1 = 1.918237500e-21
+ ub1 = -3.585450663e-18 lub1 = 7.258499312e-25 wub1 = 1.119132576e-23 pub1 = -3.146088601e-30
+ uc1 = -2.991611115e-10 luc1 = 8.520052668e-17 wuc1 = 1.063917300e-15 puc1 = -2.587560001e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.25 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {7.901161519e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -5.424834666e-08 wvth0 = -4.783014553e-07 pvth0 = 9.119142085e-14
+ k1 = 5.321541783e-01 lk1 = 4.286225147e-08 wk1 = 1.592076295e-08 pk1 = 1.778361048e-14
+ k2 = -5.235602683e-02 lk2 = -4.211280667e-09 wk2 = 4.960449301e-08 pk2 = -1.541606270e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.318673889e-01 ldsub = -7.020641044e-08 wdsub = -1.269117974e-07 pdsub = 8.012065719e-14
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = -4.126589768e-03 lcdscd = 1.923237469e-09 wcdscd = 4.782950144e-08 pcdscd = -9.655867580e-15
+ cit = 0.0
+ voff = {-2.304547281e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.820393130e-08 wvoff = 4.684822864e-07 pvoff = -9.748460659e-14
+ nfactor = -1.976982395e+00 lnfactor = 8.915874106e-07 wnfactor = 1.807172814e-05 pnfactor = -3.356816508e-12
+ eta0 = 1.237370810e+00 leta0 = -1.508799665e-07 weta0 = 5.270653056e-07 peta0 = -1.064044710e-13
+ etab = -3.163989299e-02 letab = 6.021587276e-09 wetab = 3.812806000e-07 petab = -7.624917170e-14
+ u0 = 9.129506221e-03 lu0 = 1.926051553e-09 wu0 = -2.980156909e-08 pu0 = 5.256186514e-15
+ ua = -6.164745406e-09 lua = 8.094465120e-16 wua = 7.071263799e-15 pua = -1.389037217e-21
+ ub = 7.379459720e-18 lub = -9.550070394e-25 wub = -1.287851633e-23 pub = 2.533107842e-30
+ uc = -1.938246050e-10 luc = 4.059283756e-17 wuc = 8.937468513e-16 puc = -1.394736486e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.878873057e+04 lvsat = 4.608529371e-04 wvsat = 9.945198344e-02 pvsat = -2.422619106e-9
+ a0 = 1.5
+ ags = -2.298688364e+00 lags = 4.680045702e-07 wags = -5.467183228e-12 pags = 7.210175909e-19
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 3.585833577e-03 lketa = -4.941325437e-09 wketa = -6.983965412e-08 pketa = 2.495392854e-15
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.463772615e-01 lpclm = 7.293156065e-09 wpclm = -3.041846461e-07 ppclm = -9.785650747e-14
+ pdiblc1 = 2.180020560e+00 lpdiblc1 = -2.343227284e-07 wpdiblc1 = -7.262738388e-06 ppdiblc1 = 9.393831330e-13
+ pdiblc2 = -1.294253471e-02 lpdiblc2 = 3.108971668e-09 wpdiblc2 = 1.374447547e-08 ppdiblc2 = -2.699162808e-15
+ pdiblcb = 1.007359921e+00 lpdiblcb = -1.474330323e-07 wpdiblcb = -4.415114100e-06 ppdiblcb = 5.851653889e-13
+ drout = 5.186304277e-01 ldrout = 9.717937062e-08 wdrout = 4.280565518e-06 pdrout = -8.641648474e-13
+ pscbe1 = 7.870214523e+08 lpscbe1 = 2.620122198e+00 wpscbe1 = 8.803214030e+01 ppscbe1 = -1.777201651e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.013296356e-05 lalpha0 = -7.713033915e-13 walpha0 = -2.030580133e-12 palpha0 = -1.427038016e-18
+ alpha1 = 1.694825441e+00 lalpha1 = -1.705542049e-07 walpha1 = -2.551906763e-06 palpha1 = 5.151814892e-13
+ beta0 = 1.073128899e+01 lbeta0 = 1.835314008e-06 wbeta0 = 5.311494013e-05 pbeta0 = -1.114693196e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.313850971e-01 lkt1 = 3.367385010e-09 wkt1 = 2.833466417e-07 pkt1 = -1.550150328e-14
+ kt2 = -2.907444431e-02 lkt2 = -2.310739263e-09 wkt2 = 1.031055818e-07 pkt2 = -6.539892002e-15
+ at = 1.047980119e+05 lat = -1.429860301e-02 wat = -5.497890520e-01 pat = 1.041141095e-7
+ ute = 1.494009605e+00 lute = -5.413944792e-07 wute = 5.497327555e-07 pute = 4.422353031e-13
+ ua1 = 4.297664718e-09 lua1 = -7.411978872e-16 wua1 = 7.960080158e-15 pua1 = -5.324319677e-22
+ ub1 = -1.655415541e-18 lub1 = 3.362125108e-25 wub1 = -1.160856520e-23 pub1 = 1.456776185e-30
+ uc1 = 3.050852914e-10 luc1 = -3.678534137e-17 wuc1 = -1.316928602e-15 puc1 = 2.218915515e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.26 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.490431167e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.245539371e-08 wvth0 = 5.365758418e-07 pvth0 = -4.265161196e-14
+ k1 = 7.337009731e-01 lk1 = 1.628205862e-08 wk1 = 5.236945724e-07 pk1 = -4.918210728e-14
+ k2 = -1.191116681e-01 lk2 = 4.592520064e-09 wk2 = -9.952979551e-08 pk2 = 4.251916409e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 3.219506298e-01 ldsub = -2.958078336e-09 wdsub = 4.129087547e-07 pdsub = 8.928582966e-15
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.702936505e-02 lcdscd = -2.185641009e-09 wcdscd = -7.544742815e-08 pcdscd = 6.602017172e-15
+ cit = 0.0
+ voff = {6.358791888e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.057470703e-08 wvoff = -7.419515519e-07 pvoff = 6.214861844e-14
+ nfactor = 8.233019118e+00 lnfactor = -4.549177988e-07 wnfactor = -2.900187318e-05 pnfactor = 2.851297107e-12
+ eta0 = 4.076684168e-01 leta0 = -4.145798519e-08 weta0 = -1.229319511e-06 peta0 = 1.252293151e-13
+ etab = 1.259882392e-01 letab = -1.476656842e-08 wetab = -5.351026606e-07 petab = 4.460436910e-14
+ u0 = 1.229672512e-01 lu0 = -1.308698410e-08 wu0 = -2.468069440e-07 pu0 = 3.387507237e-14
+ ua = 1.413052107e-08 lua = -1.867113527e-15 wua = -4.643578657e-14 pua = 5.667526093e-21
+ ub = -1.190724370e-17 lub = 1.588542695e-24 wub = 4.733095987e-23 pub = -5.407378089e-30
+ uc = 4.521913365e-10 luc = -4.460439081e-17 wuc = -1.185454086e-15 puc = 1.347334502e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.142616724e+04 lvsat = 1.631491388e-02 wvsat = 3.421998280e-01 pvsat = -3.443644759e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 4.486553997e-01 lketa = -6.363754488e-08 wketa = -2.217910757e-06 pketa = 2.857851579e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.240227986e+00 lpclm = -2.160935714e-07 wpclm = -5.013426888e-06 ppclm = 5.232030687e-13
+ pdiblc1 = 6.720608263e-01 lpdiblc1 = -3.545149067e-08 wpdiblc1 = -9.517669383e-07 ppdiblc1 = 1.070859072e-13
+ pdiblc2 = 1.392380302e-02 lpdiblc2 = -4.341878175e-10 wpdiblc2 = -1.666691376e-08 ppdiblc2 = 1.311521616e-15
+ pdiblcb = -7.104703304e-01 lpdiblcb = 7.911613905e-08 wpdiblcb = 1.834050907e-06 ppdiblcb = -2.389807413e-13
+ drout = 4.028640229e+00 ldrout = -3.657242319e-07 wdrout = -1.064867498e-05 pdrout = 1.104718318e-12
+ pscbe1 = 8.524974665e+08 lpscbe1 = -6.014920034e+00 wpscbe1 = -1.844929122e+02 ppscbe1 = 1.816885993e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.873285153e-05 lalpha0 = -1.905465217e-12 walpha0 = -5.649443183e-11 palpha0 = 5.755709209e-18
+ alpha1 = -1.121259363e+00 lalpha1 = 2.008338752e-07 walpha1 = 5.954449113e-06 palpha1 = -6.066452301e-13
+ beta0 = 6.128321571e+01 lbeta0 = -4.831524640e-06 wbeta0 = -1.380693513e-04 pbeta0 = 1.406664358e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.819417563e-01 lkt1 = 3.641104778e-08 wkt1 = 9.997718494e-07 pkt1 = -1.099843761e-13
+ kt2 = -1.041773440e-01 lkt2 = 7.593906249e-09 wkt2 = 2.274487717e-07 pkt2 = -2.293839622e-14
+ at = -2.058297919e+05 lat = 2.666730238e-02 wat = 1.004332286e+00 pat = -1.008449667e-7
+ ute = -1.824424930e+01 lute = 2.061706844e-06 wute = 5.112481916e-05 pute = -6.227657667e-12
+ ua1 = -2.139862697e-08 lua1 = 2.647654757e-15 wua1 = 6.456534336e-14 pua1 = -7.997590684e-21
+ ub1 = 1.277037842e-17 lub1 = -1.566275622e-24 wub1 = -3.643675183e-23 pub1 = 4.731142266e-30
+ uc1 = -3.247285595e-10 luc1 = 4.627513910e-17 wuc1 = 1.425480975e-15 puc1 = -1.397801660e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.27 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.352093468e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.017212582e-07 wvth0 = -4.036764925e-08 pvth0 = 8.054105342e-13
+ k1 = 5.343395989e-01 lk1 = 3.417320482e-07 wk1 = 1.172605686e-08 pk1 = -2.339568910e-13
+ k2 = -3.086853240e-02 lk2 = 5.876787443e-08 wk2 = 1.341677538e-08 pk2 = -2.676899059e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.081482666e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 4.788444739e-08 wvoff = 9.059768345e-09 pvoff = -1.807594199e-13
+ nfactor = 1.475816038e+00 lnfactor = 3.038838997e-05 wnfactor = 3.013720455e-06 pnfactor = -6.012939189e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.505016514e-02 lu0 = -9.409836093e-08 wu0 = -7.994137534e-09 pu0 = 1.594980808e-13
+ ua = -8.705104692e-10 lua = 3.412030810e-15 wua = 2.975976504e-16 pua = -5.937632908e-21
+ ub = 2.071732686e-18 lub = -9.783458446e-24 wub = -9.018512708e-25 pub = 1.799362923e-29
+ uc = 5.003049930e-11 luc = 4.178223299e-16 wuc = -1.875186893e-17 puc = 3.741350573e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.192345324e+00 la0 = 4.453173568e-06 wa0 = 2.928433387e-07 pa0 = -5.842775445e-12
+ ags = 4.539511377e-01 lags = -5.124688067e-07 wags = -9.535313910e-08 pags = 1.902474484e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.255574854e-25 lb0 = 5.253045924e-29
+ b1 = 7.953053588e-24 lb1 = -1.586783788e-28 wb1 = -1.607019458e-29 pb1 = 3.206306099e-34
+ keta = -1.616009329e-02 lketa = 2.095385108e-07 wketa = 1.988543961e-08 pketa = -3.967519248e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.156109759e-01 lpclm = 3.973257005e-06 wpclm = 3.856067524e-07 ppclm = -7.693580037e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 2.922291478e-03 lpdiblc2 = -9.172960639e-09 wpdiblc2 = 9.168527659e-10 ppdiblc2 = -1.829293728e-14
+ pdiblcb = 5.951584812e-01 lpdiblcb = -6.198600671e-05 wpdiblcb = -1.110223025e-22 ppdiblcb = -2.131628207e-26
+ drout = 0.56
+ pscbe1 = 8.968247800e+08 lpscbe1 = -2.061208873e+03 wpscbe1 = -4.586457013e+02 ppscbe1 = 9.150844453e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.835000775e-01 lkt1 = -6.552182248e-07 wkt1 = -8.670546958e-08 pkt1 = 1.729937211e-12
+ kt2 = -4.587846272e-02 lkt2 = 9.610423470e-08 wkt2 = -1.495924815e-09 pkt2 = 2.984651389e-14
+ at = 140000.0
+ ute = -1.641683510e+00 lute = -2.965178519e-06 wute = -5.360945041e-07 pute = 1.069609375e-11
+ ua1 = 6.824511129e-10 lua1 = -7.014505007e-15 wua1 = -8.916098068e-16 pua1 = 1.778929276e-20
+ ub1 = -1.051014948e-18 lub1 = 1.248698345e-23 wub1 = 1.081111207e-24 pub1 = -2.157020215e-29
+ uc1 = 1.297245376e-11 luc1 = 4.379194940e-17 wuc1 = 9.129727533e-18 puc1 = -1.821552373e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.28 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {0.5200869+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.55146741
+ k2 = -0.027923052
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.10574827+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 2.9989
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0303339
+ ua = -6.9949748e-10
+ ub = 1.58138e-18
+ uc = 7.0972e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.415541
+ ags = 0.4282659
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 2.1073e-24
+ b1 = 0.0
+ keta = -0.0056579
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.083531
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0024625373
+ pdiblcb = -2.5116166
+ drout = 0.56
+ pscbe1 = 793515780.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.31634
+ kt2 = -0.041061662
+ at = 140000.0
+ ute = -1.7903
+ ua1 = 3.3088e-10
+ ub1 = -4.2516e-19
+ uc1 = 1.5167332e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.29 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.176593583e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.930352273e-8
+ k1 = 5.483501070e-01 lk1 = 2.478842258e-8
+ k2 = -2.408197285e-02 lk2 = -3.054380430e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.077667525e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.605073263e-8
+ nfactor = 2.730764874e+00 lnfactor = 2.132178613e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.085791942e-02 lu0 = -4.166940074e-9
+ ua = -7.465776512e-10 lua = 3.743759184e-16
+ ub = 1.673557624e-18 lub = -7.329854995e-25
+ uc = 8.117378080e-11 luc = -8.112334692e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.555277536e+00 la0 = -1.111168307e-6
+ ags = 4.221285300e-01 lags = 4.880363581e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.189249708e-24 lb0 = -1.655541632e-29
+ b1 = 0.0
+ keta = -1.056965338e-02 lketa = 3.905767835e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.169121138e-01 lpclm = 3.184275988e-06 ppclm = 8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 1.446243820e-03 lpdiblc2 = 8.081444813e-9
+ pdiblcb = -4.968319824e+00 lpdiblcb = 1.953541169e-5
+ drout = 0.56
+ pscbe1 = 7.871095635e+08 lpscbe1 = 5.094147091e+1
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.141467060e-01 lkt1 = -1.744081253e-8
+ kt2 = -3.997479494e-02 lkt2 = -8.642637524e-9
+ at = 140000.0
+ ute = -1.817271588e+00 lute = 2.144748568e-7
+ ua1 = 3.745936823e-10 lua1 = -3.476059996e-16
+ ub1 = -4.986867121e-19 lub1 = 5.846756647e-25
+ uc1 = 3.327652623e-12 luc1 = 9.414772148e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.30 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.126050219e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.927765852e-8
+ k1 = 5.404459826e-01 lk1 = 5.602458147e-8
+ k2 = -2.340426079e-02 lk2 = -3.322204172e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.064178854e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.072017044e-8
+ nfactor = 3.659602665e+00 lnfactor = -1.538477807e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.984585582e-02 lu0 = -1.673851512e-10
+ ua = -5.156850280e-10 lua = -5.380842521e-16
+ ub = 1.274274859e-18 lub = 8.449324743e-25
+ uc = 5.726534211e-11 luc = 1.335995769e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.029984171e+00 la0 = 9.647285615e-7
+ ags = 2.062494344e-01 lags = 9.019321322e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -2.056599416e-24 lb0 = 8.127436155e-30
+ b1 = 0.0
+ keta = -1.735957830e-03 lketa = 4.147964760e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.740059450e-01 lpclm = 5.866193894e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 2.166173716e-03 lpdiblc2 = 5.236367537e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 8.081380067e+08 lpscbe1 = -3.216043418e+1
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.150856518e-01 lkt1 = -1.373021056e-8
+ kt2 = -4.269599381e-02 lkt2 = 2.111216570e-9
+ at = 1.643009185e+05 lat = -9.603433791e-2
+ ute = -1.936131845e+00 lute = 6.841964476e-7
+ ua1 = 3.247381814e-11 lua1 = 1.004410991e-15
+ ub1 = -2.950781812e-19 lub1 = -2.199610200e-25
+ uc1 = 9.861007087e-12 luc1 = 6.832868211e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.31 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.980184208e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.774896808e-8
+ k1 = 6.287345350e-01 lk1 = -1.163041665e-7
+ k2 = -6.139263891e-02 lk2 = 4.092675175e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.455643000e-01 ldsub = -5.573875314e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-6.965807302e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -6.103060895e-8
+ nfactor = 3.418716155e+00 lnfactor = -1.068296003e-6
+ eta0 = 1.537410312e-01 leta0 = -1.439337178e-7
+ etab = -5.631671063e-02 letab = -2.670815255e-8
+ u0 = 3.390031783e-02 lu0 = -8.081212522e-9
+ ua = -1.383272633e-10 lua = -1.274641703e-15
+ ub = 1.118394756e-18 lub = 1.149191885e-24
+ uc = 5.386395292e-11 luc = 1.999906463e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.420255462e+04 lvsat = -8.202886504e-3
+ a0 = 2.065297727e+00 la0 = -1.056080298e-6
+ ags = 3.146263949e-01 lags = 6.903932022e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.113198831e-24 lb0 = -3.915275817e-30
+ b1 = 0.0
+ keta = 4.960535517e-02 lketa = -9.606416860e-08 wketa = 6.938893904e-24 pketa = 2.428612866e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.374335140e-01 lpclm = 7.156112720e-7
+ pdiblc1 = 1.705248073e-01 lpdiblc1 = 4.283894585e-7
+ pdiblc2 = 6.342319838e-03 lpdiblc2 = -2.914972732e-9
+ pdiblcb = -4.861457464e-02 lpdiblcb = 4.609283956e-8
+ drout = 8.455643000e-01 ldrout = -5.573875314e-7
+ pscbe1 = 1.145718696e+09 lpscbe1 = -6.910777669e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.585827200e-09 lalpha0 = 5.350920302e-14
+ alpha1 = 6.396342990e-01 lalpha1 = 4.106088148e-7
+ beta0 = 1.322319161e+01 lbeta0 = 1.242974195e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.860578468e-01 lkt1 = 1.247990683e-7
+ kt2 = -4.711907459e-02 lkt2 = 1.074454392e-8
+ at = 1.621895531e+05 lat = -9.191320394e-2
+ ute = -1.977870160e+00 lute = 7.656646724e-7
+ ua1 = -4.878066519e-10 lua1 = 2.019936555e-15 pua1 = 8.271806126e-37
+ ub1 = 5.834418662e-19 lub1 = -1.934727609e-24 pub1 = -7.703719778e-46
+ uc1 = 1.020383967e-10 luc1 = -1.115906132e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.32 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.717879852e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.470878628e-9
+ k1 = 4.427124355e-01 lk1 = 6.076673566e-8
+ k2 = 8.470512065e-04 lk2 = -1.831802672e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.968530194e-01 ldsub = 6.010841108e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.286641533e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -4.863842250e-9
+ nfactor = 1.883906055e+00 lnfactor = 3.926605692e-7
+ eta0 = -4.380244824e-01 leta0 = 4.193566311e-07 weta0 = 6.591949209e-23 peta0 = 2.116362641e-28
+ etab = -1.600650675e-01 letab = 7.204793714e-8
+ u0 = 2.820781092e-02 lu0 = -2.662623351e-9
+ ua = -1.374538532e-09 lua = -9.791568438e-17
+ ub = 2.394112859e-18 lub = -6.513993792e-26
+ uc = 7.403259758e-11 luc = 8.009149789e-19
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.028179688e+04 lvsat = 3.360444829e-2
+ a0 = 4.640317362e-01 la0 = 4.681343750e-7
+ ags = 9.093444662e-01 lags = 1.242923697e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -6.554655739e-02 lketa = 1.354674908e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.331358446e+00 lpclm = -4.208631858e-7
+ pdiblc1 = 7.295365653e-01 lpdiblc1 = -1.037232127e-7
+ pdiblc2 = 5.255966467e-03 lpdiblc2 = -1.880893598e-9
+ pdiblcb = 2.222914927e-02 lpdiblcb = -2.134195520e-08 wpdiblcb = -7.806255642e-24 ppdiblcb = 9.974659987e-30
+ drout = -4.087838800e-01 ldrout = 6.366026685e-07 pdrout = -2.220446049e-28
+ pscbe1 = 7.601058167e+07 lpscbe1 = 3.271570623e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -2.816247674e-06 lalpha0 = 2.736703255e-12 walpha0 = -1.058791184e-27 palpha0 = 1.164670302e-33
+ alpha1 = 1.270731402e+00 lalpha1 = -1.901205267e-7
+ beta0 = 1.137577438e+01 lbeta0 = 3.001495554e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.330485209e-01 lkt1 = -2.084760183e-8
+ kt2 = -3.484510072e-02 lkt2 = -9.388186018e-10
+ at = 8.283445085e+04 lat = -1.637658988e-2
+ ute = -1.101602841e+00 lute = -6.843753974e-8
+ ua1 = 2.169780508e-09 lua1 = -5.097701682e-16
+ ub1 = -2.235363667e-18 lub1 = 7.484398209e-25
+ uc1 = -7.594942592e-11 luc1 = 5.783261332e-17 wuc1 = -2.584939414e-32 puc1 = -1.292469707e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.33 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {6.097018043e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.960341312e-8
+ k1 = 4.142983009e-01 lk1 = 7.360654324e-8
+ k2 = -5.463888719e-03 lk2 = -1.546623287e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.331531951e-01 ldsub = 8.889315138e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.348874771e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.051640481e-9
+ nfactor = 2.619917653e+00 lnfactor = 6.007091230e-8
+ eta0 = 0.49
+ etab = -0.000625
+ u0 = 2.626595586e-02 lu0 = -1.785135944e-9
+ ua = -1.186784979e-09 lua = -1.827579476e-16
+ ub = 2.016278705e-18 lub = 1.055961373e-25
+ uc = 7.692988093e-11 luc = -5.083123204e-19 wuc = 1.033975766e-31
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.022314147e+05 lvsat = 5.610593024e-3
+ a0 = 1.5
+ ags = 2.125059674e+00 lags = -4.250662343e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.205412753e-02 lketa = -1.587843621e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.635279131e-01 lpclm = -2.870705689e-8
+ pdiblc1 = 7.782704528e-01 lpdiblc1 = -1.257451305e-7
+ pdiblc2 = -1.078606283e-04 lpdiblc2 = 5.429179532e-10
+ pdiblcb = 1.365048000e-01 lpdiblcb = -7.298095053e-08 wpdiblcb = -5.551115123e-23 ppdiblcb = 2.081668171e-29
+ drout = 1.0
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.191548560e-06 lalpha0 = 2.189428516e-14
+ alpha1 = 0.85
+ beta0 = 1.712245588e+01 lbeta0 = 4.046793707e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.057206144e-01 lkt1 = 1.199153647e-8
+ kt2 = -5.292091023e-02 lkt2 = 7.229296276e-9
+ at = 6.589423514e+04 lat = -8.721628268e-3
+ ute = -2.038377412e+00 lute = 3.548730904e-7
+ ua1 = -4.578267072e-11 lua1 = 4.914007367e-16
+ ub1 = 1.195109989e-19 lub1 = -3.156832979e-25 pub1 = -1.925929944e-46
+ uc1 = 5.305567625e-11 luc1 = -4.623412548e-19
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.34 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {3.974985320e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.323639570e-08 wvth0 = 7.076518912e-07 pvth0 = -1.428614715e-13
+ k1 = 5.374248511e-01 lk1 = 4.874963215e-8
+ k2 = 1.428648426e-02 lk2 = -1.945345792e-08 wk2 = -1.516980086e-07 pk2 = 3.062494567e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 7.898336014e-01 ldsub = -4.367814573e-08 wdsub = 5.680625851e-11 pdsub = -1.146810428e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 1.170767983e-02 lcdscd = -1.273400711e-9
+ cit = 0.0
+ voff = {-1.723984696e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 5.521116205e-09 wvoff = 2.931156942e-07 pvoff = -5.917448947e-14
+ nfactor = 6.799208278e+00 lnfactor = -7.836484583e-07 wnfactor = -8.437914245e-06 pnfactor = 1.703454566e-12
+ eta0 = 1.411859226e+00 leta0 = -1.861058623e-07 weta0 = 1.402907657e-14 peta0 = -2.832203805e-21
+ etab = 1.218543674e-01 letab = -2.472625718e-08 wetab = -8.236907484e-08 petab = 1.662875120e-14
+ u0 = -5.976314886e-03 lu0 = 4.723965916e-09 wu0 = 1.582755753e-08 pu0 = -3.195283143e-15
+ ua = -3.792483549e-09 lua = 3.432830854e-16 wua = -9.446627807e-17 pua = 1.907094668e-23
+ ub = 2.661018075e-18 lub = -2.456449154e-26 wub = 1.374159492e-24 pub = -2.774166925e-31
+ uc = 1.884765684e-10 luc = -2.302746913e-17 wuc = -2.610443066e-16 puc = 5.269988566e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.804983786e+05 lvsat = -1.019001991e-02 wvsat = -1.473627941e-01 pvsat = 2.974974824e-8
+ a0 = 1.5
+ ags = -2.298690174e+00 lags = 4.680048089e-07 wags = 7.771561172e-22 pags = -1.387778781e-29
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.437387113e-01 lketa = -5.726517772e-08 wketa = -7.952531215e-07 pketa = 1.605464954e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.687629139e-02 lpclm = 5.338817915e-08 wpclm = 1.174417648e-06 ppclm = -2.370926092e-13
+ pdiblc1 = -2.243565331e-01 lpdiblc1 = 7.666620805e-8
+ pdiblc2 = -8.392336117e-03 lpdiblc2 = 2.215396149e-9
+ pdiblcb = -4.542925080e-01 lpdiblcb = 4.628980080e-8
+ drout = 1.935739668e+00 ldrout = -1.889080599e-7
+ pscbe1 = 8.161650687e+08 lpscbe1 = -3.263420225e+0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 9.460726714e-06 lalpha0 = -1.243733670e-12
+ alpha1 = 0.85
+ beta0 = 2.683064685e+01 lbeta0 = -1.555219929e-06 wbeta0 = 4.484704620e-06 pbeta0 = -9.053766533e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.995123407e-01 lkt1 = -9.449896030e-09 wkt1 = -1.149924261e-07 pkt1 = 2.321478598e-14
+ kt2 = 5.059333590e-03 lkt2 = -4.475813327e-9
+ at = -1.343167466e+05 lat = 3.169716493e-02 wat = 1.724886392e-01 pat = -3.482217897e-8
+ ute = 1.676002233e+00 lute = -3.949895867e-07 wute = -8.881784197e-22 pute = 1.110223025e-28
+ ua1 = 6.932901369e-09 lua1 = -9.174629760e-16
+ ub1 = -5.498507054e-18 lub1 = 8.184878046e-25 wub1 = -3.081487911e-39 pub1 = 3.851859889e-46
+ uc1 = -1.308925445e-10 luc1 = 3.667330950e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.35 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {1.411423877e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.104810928e-07 wvth0 = -2.068359080e-06 pvth0 = 2.232416315e-13
+ k1 = 0.90707349
+ k2 = -2.706498401e-01 lk2 = 1.812422947e-08 wk2 = 3.582112560e-07 pk2 = -3.662239805e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586906573e-01 ldsub = -6.683115145e-12 wdsub = -1.325479365e-10 pdsub = 1.350411632e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {-1.305340903e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = -1.555803990e-7
+ nfactor = -1.034356669e+01 lnfactor = 1.477157847e-06 wnfactor = 2.711115636e-05 pnfactor = -2.984792415e-12
+ eta0 = 6.941549801e-04 leta0 = -1.650485927e-15 weta0 = -3.273451064e-14 peta0 = 3.335024679e-21
+ etab = -6.563478702e-02 wetab = 4.371998422e-8
+ u0 = 7.272991649e-02 lu0 = -5.655890584e-09 wu0 = -9.505844307e-08 pu0 = 1.142847350e-14
+ ua = -1.399266490e-09 lua = 2.766322641e-17 wua = 4.739867000e-16 pua = -5.589720052e-23
+ ub = 7.092366799e-18 lub = -6.089751926e-25 wub = -1.005987160e-23 pub = 1.230514761e-30
+ uc = 1.386863297e-11 wuc = 1.385574985e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -9.331265129e+03 lvsat = 1.484490334e-02 wvsat = 3.056655796e-01 pvsat = -2.999608672e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.999038997e-01 lketa = 9.355955346e-08 wketa = 1.855590617e-06 pketa = -1.890494276e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.443916633e+00 lpclm = -1.295360881e-07 wpclm = -2.608063331e-06 ppclm = 2.617447647e-13
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 1.903873159e+01 lbeta0 = -5.276143536e-07 wbeta0 = -1.046431078e-05 pbeta0 = 1.066114446e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.711670600e-01 wkt1 = 6.103585679e-8
+ kt2 = -0.028878939
+ at = 2.599024714e+05 lat = -2.029285975e-02 wat = -4.024734915e-01 pat = 4.100440179e-8
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.36 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.152316124e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.687211961e-8
+ k1 = 5.401427619e-01 lk1 = 2.259480306e-7
+ k2 = -2.422864182e-02 lk2 = -7.371043230e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.036646356e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -4.157242546e-08 wvoff = -2.220446049e-22
+ nfactor = 2.967290218e+00 lnfactor = 6.306746162e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.109390912e-02 lu0 = -1.516361142e-8
+ ua = -7.232309792e-10 lua = 4.735279513e-16
+ ub = 1.625411302e-18 lub = -8.785073053e-25
+ uc = 4.075029938e-11 luc = 6.029797744e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.337271930e+00 la0 = 1.561615162e-6
+ ags = 4.067613777e-01 lags = 4.290556690e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.255574854e-25 lb0 = 5.253045924e-29
+ b1 = 0.0
+ keta = -6.318895283e-03 lketa = 1.318809922e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 7.522374929e-02 lpclm = 1.657452776e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 3.376037021e-03 lpdiblc2 = -1.822603774e-8
+ pdiblcb = 5.951584812e-01 lpdiblcb = -6.198600671e-05 wpdiblcb = -5.551115123e-23 ppdiblcb = -4.174438573e-26
+ drout = 0.56
+ pscbe1 = 6.698434685e+08 lpscbe1 = 2.467495241e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.264101520e-01 lkt1 = 2.009184746e-7
+ kt2 = -4.661878793e-02 lkt2 = 1.108751152e-7
+ at = 140000.0
+ ute = -1.906993821e+00 lute = 2.328261231e-6
+ ua1 = 2.411981748e-10 lua1 = 1.789321105e-15
+ ub1 = -5.159787779e-19 lub1 = 1.812005449e-24
+ uc1 = 1.749070723e-11 luc1 = -4.635570604e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.37 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {0.5200869+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.55146741
+ k2 = -0.027923052
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.10574827+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 2.9989
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0303339
+ ua = -6.9949748e-10
+ ub = 1.58138e-18
+ uc = 7.0972e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.415541
+ ags = 0.4282659
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 2.1073e-24
+ b1 = 0.0
+ keta = -0.0056579
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.083531
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0024625373
+ pdiblcb = -2.5116166
+ drout = 0.56
+ pscbe1 = 793515780.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.31634
+ kt2 = -0.041061662
+ at = 140000.0
+ ute = -1.7903
+ ua1 = 3.3088e-10
+ ub1 = -4.2516e-19
+ uc1 = 1.5167332e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.38 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.176593583e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.930352273e-8
+ k1 = 5.483501070e-01 lk1 = 2.478842258e-8
+ k2 = -2.408197285e-02 lk2 = -3.054380430e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.077667525e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.605073263e-8
+ nfactor = 2.730764874e+00 lnfactor = 2.132178613e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.085791942e-02 lu0 = -4.166940074e-9
+ ua = -7.465776512e-10 lua = 3.743759184e-16
+ ub = 1.673557624e-18 lub = -7.329854995e-25
+ uc = 8.117378080e-11 luc = -8.112334692e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.555277536e+00 la0 = -1.111168307e-06 wa0 = -3.552713679e-21
+ ags = 4.221285300e-01 lags = 4.880363581e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.189249708e-24 lb0 = -1.655541632e-29
+ b1 = 0.0
+ keta = -1.056965338e-02 lketa = 3.905767835e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.169121138e-01 lpclm = 3.184275988e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 1.446243820e-03 lpdiblc2 = 8.081444813e-9
+ pdiblcb = -4.968319824e+00 lpdiblcb = 1.953541169e-5
+ drout = 0.56
+ pscbe1 = 7.871095635e+08 lpscbe1 = 5.094147091e+1
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.141467060e-01 lkt1 = -1.744081253e-8
+ kt2 = -3.997479494e-02 lkt2 = -8.642637524e-9
+ at = 140000.0
+ ute = -1.817271588e+00 lute = 2.144748568e-7
+ ua1 = 3.745936823e-10 lua1 = -3.476059996e-16
+ ub1 = -4.986867121e-19 lub1 = 5.846756647e-25
+ uc1 = 3.327652623e-12 luc1 = 9.414772148e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.39 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.126050219e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.927765852e-8
+ k1 = 5.404459826e-01 lk1 = 5.602458147e-8
+ k2 = -2.340426079e-02 lk2 = -3.322204172e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.064178854e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.072017044e-8
+ nfactor = 3.659602665e+00 lnfactor = -1.538477807e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.984585582e-02 lu0 = -1.673851512e-10
+ ua = -5.156850280e-10 lua = -5.380842521e-16
+ ub = 1.274274859e-18 lub = 8.449324743e-25
+ uc = 5.726534211e-11 luc = 1.335995769e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.029984171e+00 la0 = 9.647285615e-7
+ ags = 2.062494344e-01 lags = 9.019321322e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -2.056599416e-24 lb0 = 8.127436155e-30
+ b1 = 0.0
+ keta = -1.735957830e-03 lketa = 4.147964760e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.740059450e-01 lpclm = 5.866193894e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 2.166173716e-03 lpdiblc2 = 5.236367537e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 8.081380067e+08 lpscbe1 = -3.216043418e+01 wpscbe1 = 1.907348633e-12
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.150856518e-01 lkt1 = -1.373021056e-8
+ kt2 = -4.269599381e-02 lkt2 = 2.111216570e-9
+ at = 1.643009184e+05 lat = -9.603433791e-2
+ ute = -1.936131845e+00 lute = 6.841964476e-7
+ ua1 = 3.247381814e-11 lua1 = 1.004410991e-15
+ ub1 = -2.950781812e-19 lub1 = -2.199610200e-25
+ uc1 = 9.861007087e-12 luc1 = 6.832868211e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.40 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.980184208e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.774896808e-8
+ k1 = 6.287345350e-01 lk1 = -1.163041665e-7
+ k2 = -6.139263891e-02 lk2 = 4.092675175e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.455643000e-01 ldsub = -5.573875314e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-6.965807302e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -6.103060895e-8
+ nfactor = 3.418716155e+00 lnfactor = -1.068296003e-6
+ eta0 = 1.537410312e-01 leta0 = -1.439337178e-7
+ etab = -5.631671062e-02 letab = -2.670815255e-8
+ u0 = 3.390031783e-02 lu0 = -8.081212522e-9
+ ua = -1.383272633e-10 lua = -1.274641703e-15
+ ub = 1.118394756e-18 lub = 1.149191885e-24
+ uc = 5.386395292e-11 luc = 1.999906463e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.420255462e+04 lvsat = -8.202886504e-3
+ a0 = 2.065297727e+00 la0 = -1.056080298e-06 wa0 = -3.552713679e-21
+ ags = 3.146263949e-01 lags = 6.903932022e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.113198831e-24 lb0 = -3.915275817e-30
+ b1 = 0.0
+ keta = 4.960535517e-02 lketa = -9.606416860e-08 wketa = 1.040834086e-23 pketa = -5.637851297e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.374335140e-01 lpclm = 7.156112720e-7
+ pdiblc1 = 1.705248073e-01 lpdiblc1 = 4.283894585e-7
+ pdiblc2 = 6.342319838e-03 lpdiblc2 = -2.914972732e-09 wpdiblc2 = -1.387778781e-23
+ pdiblcb = -4.861457464e-02 lpdiblcb = 4.609283956e-8
+ drout = 8.455643000e-01 ldrout = -5.573875314e-7
+ pscbe1 = 1.145718696e+09 lpscbe1 = -6.910777669e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.585827200e-09 lalpha0 = 5.350920302e-14
+ alpha1 = 6.396342990e-01 lalpha1 = 4.106088148e-7
+ beta0 = 1.322319161e+01 lbeta0 = 1.242974195e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.860578468e-01 lkt1 = 1.247990683e-7
+ kt2 = -4.711907459e-02 lkt2 = 1.074454392e-8
+ at = 1.621895531e+05 lat = -9.191320394e-2
+ ute = -1.977870160e+00 lute = 7.656646724e-7
+ ua1 = -4.878066519e-10 lua1 = 2.019936555e-15 pua1 = -1.654361225e-36
+ ub1 = 5.834418662e-19 lub1 = -1.934727609e-24 pub1 = -1.540743956e-45
+ uc1 = 1.020383967e-10 luc1 = -1.115906132e-16 puc1 = -1.033975766e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.41 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.717879852e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.470878628e-9
+ k1 = 4.427124355e-01 lk1 = 6.076673566e-8
+ k2 = 8.470512065e-04 lk2 = -1.831802672e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.968530194e-01 ldsub = 6.010841108e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.286641533e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -4.863842250e-9
+ nfactor = 1.883906055e+00 lnfactor = 3.926605692e-7
+ eta0 = -4.380244824e-01 leta0 = 4.193566311e-07 weta0 = -1.040834086e-22 peta0 = -3.504141421e-28
+ etab = -1.600650675e-01 letab = 7.204793714e-8
+ u0 = 2.820781092e-02 lu0 = -2.662623351e-9
+ ua = -1.374538532e-09 lua = -9.791568438e-17
+ ub = 2.394112859e-18 lub = -6.513993792e-26
+ uc = 7.403259758e-11 luc = 8.009149789e-19
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.028179688e+04 lvsat = 3.360444829e-2
+ a0 = 4.640317362e-01 la0 = 4.681343750e-7
+ ags = 9.093444662e-01 lags = 1.242923697e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -6.554655739e-02 lketa = 1.354674908e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.331358446e+00 lpclm = -4.208631858e-7
+ pdiblc1 = 7.295365653e-01 lpdiblc1 = -1.037232127e-7
+ pdiblc2 = 5.255966467e-03 lpdiblc2 = -1.880893598e-9
+ pdiblcb = 2.222914927e-02 lpdiblcb = -2.134195520e-08 wpdiblcb = 3.469446952e-24 ppdiblcb = -1.170938346e-29
+ drout = -4.087838800e-01 ldrout = 6.366026685e-07 pdrout = 4.440892099e-28
+ pscbe1 = 7.601058167e+07 lpscbe1 = 3.271570623e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -2.816247674e-06 lalpha0 = 2.736703255e-12 walpha0 = -8.470329473e-28 palpha0 = 1.270549421e-33
+ alpha1 = 1.270731402e+00 lalpha1 = -1.901205267e-7
+ beta0 = 1.137577438e+01 lbeta0 = 3.001495554e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.330485209e-01 lkt1 = -2.084760183e-8
+ kt2 = -3.484510072e-02 lkt2 = -9.388186018e-10
+ at = 8.283445085e+04 lat = -1.637658988e-2
+ ute = -1.101602841e+00 lute = -6.843753974e-8
+ ua1 = 2.169780508e-09 lua1 = -5.097701682e-16
+ ub1 = -2.235363667e-18 lub1 = 7.484398209e-25 pub1 = -1.540743956e-45
+ uc1 = -7.594942592e-11 luc1 = 5.783261332e-17 puc1 = -2.584939414e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.42 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {6.097018043e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.960341312e-8
+ k1 = 4.142983009e-01 lk1 = 7.360654324e-8
+ k2 = -5.463888719e-03 lk2 = -1.546623287e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.331531951e-01 ldsub = 8.889315138e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.348874771e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.051640481e-9
+ nfactor = 2.619917653e+00 lnfactor = 6.007091230e-8
+ eta0 = 0.49
+ etab = -0.000625
+ u0 = 2.626595586e-02 lu0 = -1.785135944e-9
+ ua = -1.186784979e-09 lua = -1.827579476e-16
+ ub = 2.016278705e-18 lub = 1.055961373e-25
+ uc = 7.692988093e-11 luc = -5.083123204e-19
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.022314147e+05 lvsat = 5.610593024e-3
+ a0 = 1.5
+ ags = 2.125059674e+00 lags = -4.250662343e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.205412753e-02 lketa = -1.587843621e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.635279131e-01 lpclm = -2.870705689e-8
+ pdiblc1 = 7.782704528e-01 lpdiblc1 = -1.257451305e-7
+ pdiblc2 = -1.078606283e-04 lpdiblc2 = 5.429179532e-10
+ pdiblcb = 1.365048000e-01 lpdiblcb = -7.298095053e-08 wpdiblcb = 5.551115123e-23 ppdiblcb = -2.775557562e-29
+ drout = 1.0
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.191548560e-06 lalpha0 = 2.189428516e-14
+ alpha1 = 0.85
+ beta0 = 1.712245588e+01 lbeta0 = 4.046793707e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.057206144e-01 lkt1 = 1.199153647e-8
+ kt2 = -5.292091023e-02 lkt2 = 7.229296276e-9
+ at = 6.589423514e+04 lat = -8.721628268e-3
+ ute = -2.038377412e+00 lute = 3.548730904e-07 wute = -3.552713679e-21
+ ua1 = -4.578267072e-11 lua1 = 4.914007367e-16
+ ub1 = 1.195109989e-19 lub1 = -3.156832979e-25
+ uc1 = 5.305567625e-11 luc1 = -4.623412548e-19
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.43 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {6.662796355e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.102540225e-08 wvth0 = 1.645441925e-07 pvth0 = -3.321834613e-14
+ k1 = 5.374248511e-01 lk1 = 4.874963215e-8
+ k2 = -9.958667004e-02 lk2 = 3.535368344e-09 wk2 = 7.839773097e-08 pk2 = -1.582701233e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 7.898617145e-01 ldsub = -4.368382123e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 1.170767983e-02 lcdscd = -1.273400711e-9
+ cit = 0.0
+ voff = {-2.733707583e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.376402303e-8
+ nfactor = 2.447108696e+00 lnfactor = 9.495775730e-08 wnfactor = 3.560774361e-07 pnfactor = -7.188526889e-14
+ eta0 = 1.411859233e+00 leta0 = -1.861058637e-7
+ etab = 8.109035161e-02 letab = -1.649677690e-08 wetab = -3.122502257e-23 petab = -9.540979118e-30
+ u0 = -4.287039806e-03 lu0 = 4.382933374e-09 wu0 = 1.241415425e-08 pu0 = -2.506181874e-15
+ ua = -3.804200505e-09 lua = 3.456485162e-16 wua = -7.079062211e-17 pua = 1.429128158e-23
+ ub = 2.634767189e-18 lub = -1.926493632e-26 wub = 1.427202874e-24 pub = -2.881251434e-31
+ uc = -1.223104284e-10 luc = 3.971452056e-17 wuc = 3.669418443e-16 puc = -7.407858647e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.771364931e+05 lvsat = -9.511319092e-03 wvsat = -1.405696606e-01 pvsat = 2.837834365e-8
+ a0 = 1.5
+ ags = -2.298690174e+00 lags = 4.680048089e-07 wags = 9.992007222e-22 pags = -1.665334537e-28
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.342389045e-01 lketa = 5.941752133e-08 wketa = 3.726269443e-07 pketa = -7.522630013e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.153354978e-01 lpclm = -3.916602391e-08 wpclm = 2.480403049e-07 ppclm = -5.007462480e-14
+ pdiblc1 = -2.243565331e-01 lpdiblc1 = 7.666620805e-8
+ pdiblc2 = -8.392336117e-03 lpdiblc2 = 2.215396149e-9
+ pdiblcb = -4.542925080e-01 lpdiblcb = 4.628980080e-08 wpdiblcb = 8.881784197e-22
+ drout = 1.935739668e+00 ldrout = -1.889080599e-07 wdrout = 3.552713679e-21
+ pscbe1 = 8.161650687e+08 lpscbe1 = -3.263420225e+0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 9.460726714e-06 lalpha0 = -1.243733670e-12
+ alpha1 = 0.85
+ beta0 = 2.864960137e+01 lbeta0 = -1.922432287e-06 wbeta0 = 8.092669003e-07 pbeta0 = -1.633756111e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.617054272e-02 lkt1 = -3.838788156e-08 wkt1 = -4.046334502e-07 pkt1 = 8.168780555e-14
+ kt2 = 5.059333590e-03 lkt2 = -4.475813327e-9
+ at = -4.895303898e+04 lat = 1.446385428e-2
+ ute = 1.676002233e+00 lute = -3.949895867e-07 pute = 2.220446049e-28
+ ua1 = 6.932901369e-09 lua1 = -9.174629760e-16
+ ub1 = -5.498507054e-18 lub1 = 8.184878046e-25
+ uc1 = -1.308925445e-10 luc1 = 3.667330950e-17 puc1 = -2.584939414e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.44 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.310266252e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = -8.733701955e-8
+ k1 = 0.90707349
+ k2 = -7.277940937e-02 wk2 = -4.161206821e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.45862506
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 3.167134760e+00 wnfactor = -1.889993292e-7
+ eta0 = 0.00069413878
+ etab = -0.043998
+ u0 = 2.894696186e-02 wu0 = -6.589203885e-9
+ ua = -1.183288348e-09 wua = 3.757435527e-17
+ ub = 2.488689010e-18 wub = -7.575329362e-25
+ uc = 1.788286331e-10 wuc = -1.947659564e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.050160277e+05 wvsat = 7.461178063e-2
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.163000005e-01 wketa = -1.977835025e-7
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.183554635e-01 wpclm = -1.316552145e-7
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 1.407257900e+01 wbeta0 = -4.295439299e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.472502400e-01 wkt1 = 2.147719650e-7
+ kt2 = -0.028878939
+ at = 60720.487
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.45 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.046439939e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.922532212e-08 wvth0 = 1.800564292e-08 pvth0 = 2.144453445e-13
+ k1 = 4.463345813e-01 lk1 = 6.839831817e-06 wk1 = 1.595331939e-07 pk1 = -1.124778241e-11
+ k2 = 8.170793039e-03 lk2 = -2.410917766e-06 wk2 = -5.509951570e-08 pk2 = 3.974729583e-12
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.016224261e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.625656350e-07 wvoff = -3.473046787e-09 pvoff = -5.172269181e-13
+ nfactor = 2.591192879e+00 lnfactor = 3.051173988e-05 wnfactor = 6.396031696e-07 pnfactor = -5.081669577e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.242139722e-02 lu0 = 3.754040671e-08 wu0 = -2.257568748e-09 pu0 = -8.963013978e-14
+ ua = -7.654241679e-10 lua = -1.098493663e-15 wua = 7.175508696e-17 pua = 2.673430262e-21
+ ub = 1.703258241e-18 lub = 2.081096182e-24 wub = -1.323889943e-25 pub = -5.033196398e-30
+ uc = -8.575107727e-11 luc = 5.875053767e-15 wuc = 2.151322892e-16 puc = -8.965857737e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.070887868e+00 la0 = 9.095036609e-06 wa0 = 4.530212613e-07 pa0 = -1.281157758e-11
+ ags = 2.660327294e-01 lags = 9.249552716e-06 wags = 2.393276427e-07 pags = -1.500041953e-11
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.015595577e-23 lb0 = 3.728742072e-28 wb0 = 1.637776350e-29 pb0 = -5.447868288e-34
+ b1 = 0.0
+ keta = -5.197856155e-03 lketa = -2.600983866e-07 wketa = -1.906475013e-09 pketa = 4.647597429e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.989391336e-02 lpclm = 6.711231498e-07 wpclm = 4.307672954e-08 ppclm = -8.594617816e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 6.684473099e-03 lpdiblc2 = -1.260805468e-07 wpdiblc2 = -5.626432263e-09 ppdiblc2 = 1.834208295e-13
+ pdiblcb = 1.029096104e+01 lpdiblcb = -2.732643605e-04 wpdiblcb = -1.648899210e-05 ppdiblcb = 3.593067294e-10
+ drout = 0.56
+ pscbe1 = 2.684154712e+08 lpscbe1 = 1.242360350e+04 wpscbe1 = 6.826812980e+02 ppscbe1 = -1.693167630e-2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.389710282e-01 lkt1 = -1.000009542e-06 wkt1 = 2.136142804e-08 pkt1 = 2.042336614e-12
+ kt2 = -4.803101803e-02 lkt2 = -1.103519029e-06 wkt2 = 2.401683697e-09 pkt2 = 2.065237542e-12
+ at = 140000.0
+ ute = -1.880607096e+00 lute = -2.877425423e-05 wute = -4.487410903e-08 pute = 5.289393308e-11
+ ua1 = 7.454714832e-10 lua1 = -7.048982370e-14 wua1 = -8.575833251e-16 pua1 = 1.229202266e-19
+ ub1 = -1.185971500e-18 lub1 = 4.662562249e-23 wub1 = 1.139411064e-24 pub1 = -7.621147117e-29
+ uc1 = -5.520219894e-12 luc1 = 2.820370441e-15 wuc1 = 3.913311901e-17 puc1 = -4.875246221e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.46 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.031792036e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = 2.875376961e-8
+ k1 = 7.891509712e-01 wk1 = -4.042122700e-7
+ k2 = -1.126658221e-01 wk2 = 1.441162666e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-8.846248221e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = -2.939676386e-8
+ nfactor = 4.120459211e+00 wnfactor = -1.907359484e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.430294446e-02 wu0 = -6.749884023e-9
+ ua = -8.204813158e-10 wua = 2.057489827e-16
+ ub = 1.807564004e-18 wub = -3.846557554e-25
+ uc = 2.087100698e-10 wuc = -2.342417692e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.526736447e+00 wa0 = -1.891025356e-7
+ ags = 7.296257468e-01 wags = -5.125021990e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 8.532718604e-24 wb0 = -1.092727249e-29
+ b1 = 0.0
+ keta = -1.823414013e-02 wketa = 2.138755641e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.083531
+ pdiblc1 = 0.39
+ pdiblc2 = 3.652420048e-04 wpdiblc2 = 3.566727492e-9
+ pdiblcb = -3.405209289e+00 wpdiblcb = 1.519672322e-6
+ drout = 0.56
+ pscbe1 = 8.910937792e+08 wpscbe1 = -1.659442679e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.890920941e-01 wkt1 = 1.237245393e-7
+ kt2 = -1.033400402e-01 wkt2 = 1.059126029e-7
+ at = 140000.0
+ ute = -3.322789627e+00 wute = 2.606200899e-6
+ ua1 = -2.787519902e-09 wua1 = 5.303250663e-15
+ ub1 = 1.150932097e-18 wub1 = -2.680352655e-24
+ uc1 = 1.358384039e-10 wuc1 = -2.052170864e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.47 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.918224778e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.030733221e-08 wvth0 = 4.393902584e-08 pvth0 = -1.207513505e-13
+ k1 = 8.269486171e-01 lk1 = -3.005623821e-07 wk1 = -4.737935414e-07 pk1 = 5.533019897e-13
+ k2 = -1.207846379e-01 lk2 = 6.455985656e-08 wk2 = 1.644556466e-07 pk2 = -1.617363290e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-8.034677303e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -6.453515364e-08 wvoff = -4.663129453e-08 pvoff = 1.370469370e-13
+ nfactor = 3.781019545e+00 lnfactor = 2.699183832e-06 wnfactor = -1.786096701e-06 pnfactor = -9.642672200e-13
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.354818157e-02 lu0 = 6.001784707e-09 wu0 = -4.575145900e-09 pu0 = -1.729325876e-14
+ ua = -1.122191356e-09 lua = 2.399162336e-15 wua = 6.387806861e-16 pua = -3.443416575e-21
+ ub = 2.179718138e-18 lub = -2.959325385e-24 wub = -8.607927664e-25 pub = 3.786184851e-30
+ uc = 2.487470922e-10 luc = -3.183696372e-16 wuc = -2.849805357e-16 puc = 4.034686332e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.736298414e+00 la0 = -1.666411821e-06 wa0 = -3.078498971e-07 pa0 = 9.442648878e-13
+ ags = 6.749425468e-01 lags = 4.348342995e-07 wags = -4.299436069e-07 pags = -6.564960996e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.696279074e-23 lb0 = -6.703493042e-29 wb0 = -2.172309263e-29 pb0 = 8.584707701e-35
+ b1 = 0.0
+ keta = -4.101616908e-03 lketa = -1.123801429e-07 wketa = -1.099974980e-08 pketa = 2.575400048e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.834307373e-01 lpclm = 2.122847967e-06 wpclm = -2.270027002e-07 ppclm = 1.805098459e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -3.164631714e-03 lpdiblc2 = 2.806913576e-08 wpdiblc2 = 7.841402481e-09 ppdiblc2 = -3.399170683e-14
+ pdiblcb = -6.744755505e+00 lpdiblcb = 2.655567411e-05 wpdiblcb = 3.021063365e-06 ppdiblcb = -1.193888291e-11
+ drout = 0.56
+ pscbe1 = 8.160956676e+08 lpscbe1 = 5.963760582e+02 wpscbe1 = -4.929469617e+01 ppscbe1 = -9.275835130e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.839164810e-01 lkt1 = -4.115585972e-08 wkt1 = 1.186527119e-07 pkt1 = 4.033056814e-14
+ kt2 = -9.912512098e-02 lkt2 = -3.351653607e-08 wkt2 = 1.005929373e-07 pkt2 = 4.230134783e-14
+ at = 140000.0
+ ute = -2.822884827e+00 lute = -3.975183481e-06 wute = 1.710178054e-06 pute = 7.125067038e-12
+ ua1 = -2.303549787e-09 lua1 = -3.848472769e-15 wua1 = 4.554536484e-15 pua1 = 5.953686055e-21
+ ub1 = 8.345060618e-19 lub1 = 2.516182178e-24 wub1 = -2.267270293e-24 pub1 = -3.284781785e-30
+ uc1 = 1.063448109e-10 luc1 = 2.345295422e-16 wuc1 = -1.751942759e-16 puc1 = -2.387378165e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.48 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.283092312e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -5.388397538e-08 wvth0 = -2.670708074e-08 pvth0 = 1.584336558e-13
+ k1 = 8.398052416e-01 lk1 = -3.513702322e-07 wk1 = -5.090999353e-07 pk1 = 6.928286568e-13
+ k2 = -1.394063219e-01 lk2 = 1.381505361e-07 wk2 = 1.972768172e-07 pk2 = -2.914416897e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.666941931e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.766995752e-07 wvoff = 1.025078177e-07 pvoff = -4.523330871e-13
+ nfactor = 4.876145054e+00 lnfactor = -1.628621860e-06 wnfactor = -2.068890915e-06 pnfactor = 1.533018613e-13
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.251245339e-02 lu0 = 1.009485921e-08 wu0 = -4.534901168e-09 pu0 = -1.745230115e-14
+ ua = -1.334666642e-09 lua = 3.238839383e-15 wua = 1.392786341e-15 pua = -6.423157195e-21
+ ub = 2.288211241e-18 lub = -3.388077216e-24 wub = -1.724332657e-24 pub = 7.198791736e-30
+ uc = 2.399518433e-10 luc = -2.836118602e-16 wuc = -3.106825098e-16 puc = 5.050397765e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = -1.475991584e-02 la0 = 5.253562321e-06 wa0 = 1.776725226e-06 pa0 = -7.293727935e-12
+ ags = 2.069154692e-01 lags = 2.284421615e-06 wags = -1.132680112e-09 pags = -2.351105854e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -8.327425661e-24 lb0 = 3.290899525e-29 wb0 = 1.066436778e-29 pb0 = -4.214431240e-35
+ b1 = 0.0
+ keta = -9.214740762e-02 lketa = 2.355663445e-07 wketa = 1.537566047e-07 pketa = -3.935575020e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.648479260e-01 lpclm = -4.388406556e-08 wpclm = 1.856376202e-07 ppclm = 1.743930167e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 4.382386258e-03 lpdiblc2 = -1.755781171e-09 wpdiblc2 = -3.768961967e-09 ppdiblc2 = 1.189107184e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 1.162943907e+09 lpscbe1 = -7.743269107e+02 wpscbe1 = -6.033942685e+02 ppscbe1 = 1.262152059e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.742218610e-01 lkt1 = -7.946784418e-08 wkt1 = 1.005689297e-07 pkt1 = 1.117955233e-13
+ kt2 = -1.008433599e-01 lkt2 = -2.672626044e-08 wkt2 = 9.888727145e-08 pkt2 = 4.904193620e-14
+ at = 1.526954411e+05 lat = -5.017087259e-02 wat = 1.973664610e-02 pat = -7.799687674e-8
+ ute = -2.556793238e+00 lute = -5.026745773e-06 wute = 1.055516627e-06 pute = 9.712211091e-12
+ ua1 = 2.106856118e-09 lua1 = -2.127787207e-14 wua1 = -3.527760919e-15 pua1 = 3.789396360e-20
+ ub1 = -3.623872137e-18 lub1 = 2.013516227e-23 wub1 = 5.661053523e-24 pub1 = -3.461657404e-29
+ uc1 = 6.016646178e-11 luc1 = 4.170208827e-16 wuc1 = -8.555106602e-17 puc1 = -5.929971144e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.49 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.371360412e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.240752418e-07 wvth0 = 1.035385231e-07 pvth0 = -9.579026361e-14
+ k1 = 7.264654260e-01 lk1 = -1.301443997e-07 wk1 = -1.662042806e-07 pk1 = 2.353714356e-14
+ k2 = -9.744117932e-02 lk2 = 5.623957154e-08 wk2 = 6.130530139e-08 pk2 = -2.604147135e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.455643000e-01 ldsub = -5.573875314e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {2.768516321e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.027057972e-07 wvoff = -1.655450225e-07 pvoff = 7.087415877e-14
+ nfactor = 5.044109474e+00 lnfactor = -1.956468421e-06 wnfactor = -2.764195892e-06 pnfactor = 1.510454435e-12
+ eta0 = 1.537411763e-01 leta0 = -1.439340010e-07 weta0 = -2.467959727e-13 peta0 = 4.817163701e-19
+ etab = -5.631671062e-02 letab = -2.670815255e-8
+ u0 = 4.966215914e-02 lu0 = -2.337932560e-08 wu0 = -2.680509171e-08 pu0 = 2.601646064e-14
+ ua = 2.295668253e-09 lua = -3.847142323e-15 wua = -4.139330663e-15 pua = 4.374876875e-21
+ ub = -1.489682992e-18 lub = 3.985922757e-24 wub = 4.435380478e-24 pub = -4.824235296e-30
+ uc = 9.974607936e-11 luc = -9.946893485e-18 wuc = -7.802861246e-17 puc = 5.092705464e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.260406942e+05 lvsat = -8.986595616e-02 wvsat = -7.115127893e-02 pvsat = 1.388788295e-7
+ a0 = 3.915454724e+00 la0 = -2.417748960e-06 wa0 = -3.146436193e-06 pa0 = 2.315697300e-12
+ ags = 2.354306315e-01 lags = 2.228763411e-06 wags = 1.346828495e-07 pags = -2.616201606e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.665485132e-23 lb0 = -1.585343653e-29 wb0 = -2.132873556e-29 pb0 = 2.030241813e-35
+ b1 = 0.0
+ keta = 2.811759188e-01 lketa = -4.931163632e-07 wketa = -3.938163108e-07 pketa = 6.752396677e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.612977447e-01 lpclm = 2.154218272e-06 wpclm = 1.528411138e-06 ppclm = -2.446541100e-12
+ pdiblc1 = -6.475620940e-01 lpdiblc1 = 2.025197738e-06 wpdiblc1 = 1.391264763e-06 ppdiblc1 = -2.715583257e-12
+ pdiblc2 = 1.100942146e-02 lpdiblc2 = -1.469096526e-08 wpdiblc2 = -7.937022360e-09 ppdiblc2 = 2.002662973e-14
+ pdiblcb = -1.913572701e-01 lpdiblcb = 3.247095948e-07 wpdiblcb = 2.427527957e-07 ppdiblcb = -4.738245697e-13
+ drout = 1.244063683e+00 ldrout = -1.335210906e-06 wdrout = -6.777008033e-07 pdrout = 1.322791322e-12
+ pscbe1 = 2.199857802e+09 lpscbe1 = -2.798259440e+03 wpscbe1 = -1.792702697e+03 ppscbe1 = 3.583540584e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -8.448626343e-08 lalpha0 = 2.234635623e-13 walpha0 = 1.480775836e-13 palpha0 = -2.890298220e-19
+ alpha1 = -4.458644308e-01 lalpha1 = 2.529373161e-06 walpha1 = 1.846033876e-06 palpha1 = -3.603238448e-12
+ beta0 = 1.128148399e+01 lbeta0 = 5.032956408e-06 wbeta0 = 3.302130115e-06 pbeta0 = -6.445365031e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.721273846e-01 lkt1 = 3.068201871e-07 wkt1 = 3.164358102e-07 pkt1 = -3.095509394e-13
+ kt2 = -1.906010285e-01 lkt2 = 1.484700275e-07 wkt2 = 2.440100022e-07 pkt2 = -2.342203647e-13
+ at = 2.436952724e+05 lat = -2.277917142e-01 wat = -1.386112344e-01 pat = 2.310793427e-7
+ ute = -8.532535100e+00 lute = 6.637191227e-06 wute = 1.114707295e-05 pute = -9.985305948e-12
+ ua1 = -1.984710257e-08 lua1 = 2.157364277e-14 wua1 = 3.292303814e-14 pua1 = -3.325365851e-20
+ ub1 = 1.641876322e-17 lub1 = -1.898567687e-23 wub1 = -2.693005422e-23 pub1 = 2.899738994e-29
+ uc1 = 6.453970251e-10 luc1 = -7.252795345e-16 wuc1 = -9.240530710e-16 puc1 = 1.043659017e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.50 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.669403964e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.169424222e-10 wvth0 = 8.243964686e-09 pvth0 = -5.081184088e-15
+ k1 = 5.633377937e-01 lk1 = 2.513369407e-08 wk1 = -2.051393442e-07 pk1 = 6.059869079e-14
+ k2 = -2.280293751e-02 lk2 = -1.480715271e-08 wk2 = 4.021992761e-08 pk2 = -5.970704681e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.513422935e-01 ldsub = 1.034292063e-07 wdsub = 7.739699676e-08 pdsub = -7.367273068e-14
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-4.326375067e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -3.517087412e-08 wvoff = -1.452346575e-07 pvoff = 5.154110823e-14
+ nfactor = 4.634141424e+00 lnfactor = -1.566227623e-06 wnfactor = -4.677138275e-06 pnfactor = 3.331347944e-12
+ eta0 = -4.380247727e-01 leta0 = 4.193567623e-07 weta0 = 4.935919454e-13 peta0 = -2.230448218e-19
+ etab = -1.592039168e-01 letab = 7.122822415e-08 wetab = -1.464500433e-09 petab = 1.394030137e-15
+ u0 = 2.692835647e-02 lu0 = -1.739450781e-09 wu0 = 2.175881174e-09 pu0 = -1.569976814e-15
+ ua = -1.582197262e-09 lua = -1.558758191e-16 wua = 3.531510806e-16 pua = 9.856885987e-23
+ ub = 2.597637688e-18 lub = 9.527986099e-26 wub = -3.461208369e-25 pub = -2.728150434e-31
+ uc = 1.062704388e-10 luc = -1.615730730e-17 wuc = -5.482470444e-17 puc = 2.883969547e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -6.197191399e+04 lvsat = 8.909967330e-02 wvsat = 1.738959328e-01 pvsat = -9.437695549e-8
+ a0 = 1.262952997e+00 la0 = 1.071170370e-07 wa0 = -1.358671061e-06 pa0 = 6.139576376e-13
+ ags = 3.589508145e+00 lags = -9.639192459e-07 wags = -4.557972117e-06 pags = 1.850647496e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -4.079831376e-01 lketa = 1.628810486e-07 wketa = 5.823586062e-07 pketa = -2.539626884e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.773170251e+00 lpclm = -1.210174658e-06 wpclm = -2.451991294e-06 ppclm = 1.342328347e-12
+ pdiblc1 = 1.379504193e+00 lpdiblc1 = 9.567185343e-08 wpdiblc1 = -1.105355746e-06 ppdiblc1 = -3.390976300e-13
+ pdiblc2 = -7.999467485e-03 lpdiblc2 = 3.403234953e-09 wpdiblc2 = 2.254261515e-08 ppdiblc2 = -8.986358106e-15
+ pdiblcb = 3.077145403e-01 lpdiblcb = -1.503473792e-07 wpdiblcb = -4.855055915e-07 ppdiblcb = 2.193907522e-13
+ drout = -1.205782647e+00 ldrout = 9.967512681e-07 wdrout = 1.355401607e-06 pdrout = -6.124802333e-13
+ pscbe1 = -2.131522792e+09 lpscbe1 = 1.324699451e+03 wpscbe1 = 3.754201896e+03 ppscbe1 = -1.696452507e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.148784346e-05 lalpha0 = 1.107810261e-11 walpha0 = 1.474719328e-11 palpha0 = -1.418565067e-17
+ alpha1 = 3.441728862e+00 lalpha1 = -1.171153030e-06 walpha1 = -3.692067752e-06 palpha1 = 1.668375268e-12
+ beta0 = 3.801062902e+00 lbeta0 = 1.215342711e-05 wbeta0 = 1.288179673e-05 pbeta0 = -1.556406767e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.000322750e-01 lkt1 = -4.737007786e-08 wkt1 = -5.614848424e-08 pkt1 = 4.510497145e-14
+ kt2 = -3.097212644e-02 lkt2 = -3.477691373e-09 wkt2 = -6.586503998e-09 pkt2 = 4.317688280e-15
+ at = -2.400858317e+04 lat = 2.703049951e-02 wat = 1.817006826e-01 pat = -7.381948525e-8
+ ute = -1.762371008e+00 lute = 1.928006612e-07 wute = 1.123723490e-06 pute = -4.442700441e-13
+ ua1 = 4.564833092e-09 lua1 = -1.663614957e-15 wua1 = -4.073103065e-15 pua1 = 1.962265370e-21
+ ub1 = -6.467945166e-18 lub1 = 2.799745996e-24 wub1 = 7.198063539e-24 pub1 = -3.488516924e-30
+ uc1 = -3.042591023e-10 luc1 = 1.786800897e-16 wuc1 = 3.882707415e-16 puc1 = -2.055170855e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.51 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.800668252e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -5.414641357e-09 wvth0 = 5.039819382e-08 pvth0 = -2.412987930e-14
+ k1 = 8.053886150e-01 lk1 = -8.424447309e-08 wk1 = -6.651007031e-07 pk1 = 2.684464896e-13
+ k2 = -1.583737549e-01 lk2 = 4.645472381e-08 wk2 = 2.600434115e-07 pk2 = -1.053047604e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -5.860802927e-02 ldsub = 1.983017681e-07 wdsub = 3.261152745e-07 pdsub = -1.860637947e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = -2.843581713e-03 lcdscd = 3.725117948e-09 wcdscd = 1.401929886e-08 pcdscd = -6.335054787e-15
+ cit = 0.0
+ voff = {-1.840647861e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.845443856e-08 wvoff = 8.363250538e-08 pvoff = -5.187961421e-14
+ nfactor = -5.889213915e-01 lnfactor = 7.939752252e-07 wnfactor = 5.457054362e-06 pnfactor = -1.248101159e-12
+ eta0 = -7.147887813e-01 leta0 = 5.444211593e-07 weta0 = 2.048902355e-06 peta0 = -9.258600450e-13
+ etab = -1.091420653e-01 letab = 4.860622465e-08 wetab = 1.845475938e-07 petab = -8.266130104e-14
+ u0 = 5.570535131e-02 lu0 = -1.474322799e-08 wu0 = -5.006557797e-08 pu0 = 2.203694599e-14
+ ua = 4.460266351e-10 lua = -1.072391662e-15 wua = -2.776811682e-15 pua = 1.512939563e-21
+ ub = 2.313507692e-18 lub = 2.236728076e-25 wub = -5.054771266e-25 pub = -2.008049639e-31
+ uc = 1.120524070e-10 luc = -1.877006886e-17 wuc = -5.973049174e-17 puc = 3.105652754e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.599730724e+05 lvsat = -1.119304909e-02 wvsat = -9.819731074e-02 pvsat = 2.857681150e-8
+ a0 = 1.5
+ ags = 5.646384181e+00 lags = -1.893382446e-06 wags = -5.988477139e-06 pags = 2.497065536e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.601185496e-01 lketa = 5.087575068e-08 wketa = 2.177904542e-07 pketa = -8.922126730e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.913835700e-01 lpclm = 1.746389874e-07 wpclm = 1.283826625e-06 ppclm = -3.458167900e-13
+ pdiblc1 = 3.246994879e+00 lpdiblc1 = -7.482117054e-07 wpdiblc1 = -4.198391759e-06 ppdiblc1 = 1.058586576e-12
+ pdiblc2 = 1.141089214e-02 lpdiblc2 = -5.367937763e-09 wpdiblc2 = -1.958915955e-08 ppdiblc2 = 1.005219038e-14
+ pdiblcb = 4.361699030e-01 lpdiblcb = -2.083939169e-07 wpdiblcb = -5.096200635e-07 ppdiblcb = 2.302876239e-13
+ drout = -2.229292901e-01 ldrout = 5.526185105e-07 wdrout = 2.079752684e-06 pdrout = -9.398007228e-13
+ pscbe1 = 7.788736797e+08 lpscbe1 = 9.546582739e+00 wpscbe1 = 3.592809633e+01 ppscbe1 = -1.623522410e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.281081873e-05 lalpha0 = 9.799884539e-14 walpha0 = -1.635883866e-11 palpha0 = -1.294258505e-19
+ alpha1 = 0.85
+ beta0 = 2.820271850e+01 lbeta0 = 1.126782581e-06 wbeta0 = -1.884344917e-05 pbeta0 = -1.228031827e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.389331836e-01 lkt1 = 1.539660359e-08 wkt1 = 5.648235785e-08 pkt1 = -5.790766104e-15
+ kt2 = -8.505086596e-02 lkt2 = 2.095946352e-08 wkt2 = 5.464123086e-08 pkt2 = -2.334996178e-14
+ at = 6.124382814e+04 lat = -1.149344536e-02 wat = 7.908630971e-03 pat = 4.713840850e-9
+ ute = -4.744812944e+00 lute = 1.540509506e-06 wute = 4.602650871e-06 pute = -2.016331228e-12
+ ua1 = -6.271403471e-09 lua1 = 3.233074458e-15 wua1 = 1.058748995e-14 pua1 = -4.662578063e-21
+ ub1 = 5.972866688e-18 lub1 = -2.822020505e-24 wub1 = -9.954403992e-24 pub1 = 4.262357257e-30
+ uc1 = 3.611814308e-10 luc1 = -1.220198438e-16 wuc1 = -5.240085183e-16 puc1 = 2.067245787e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.52 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {9.150124452e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.303379808e-08 wvth0 = -2.584587832e-07 pvth0 = 3.822247608e-14
+ k1 = -5.896796149e-01 lk1 = 1.973932962e-07 wk1 = 1.916789922e-06 pk1 = -2.527881717e-13
+ k2 = 4.369275373e-01 lk2 = -7.372529636e-08 wk2 = -8.340154985e-07 pk2 = 1.155649464e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.799799843e+00 ldsub = -1.768754716e-07 wdsub = -1.717533100e-06 pdsub = 2.265099828e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 4.114904309e-02 lcdscd = -5.156157140e-09 wcdscd = -5.006892449e-08 pcdscd = 6.603139830e-15
+ cit = 0.0
+ voff = {2.666359916e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -6.253348514e-08 wvoff = -4.999400056e-07 pvoff = 6.593258788e-14
+ nfactor = 3.604610684e+00 lnfactor = -5.261922369e-08 wnfactor = -1.612407483e-06 pnfactor = 1.790888674e-13
+ eta0 = 5.714676309e+00 leta0 = -7.535656826e-07 weta0 = -7.317508410e-06 peta0 = 9.650403266e-13
+ etab = 4.625002228e-01 letab = -6.679749212e-08 wetab = -6.486378321e-07 petab = 8.554300593e-14
+ u0 = -1.022338346e-01 lu0 = 1.714169281e-08 wu0 = 1.789856078e-07 pu0 = -2.420413644e-14
+ ua = -1.172134803e-08 lua = 1.383970103e-15 wua = 1.339336381e-14 pua = -1.751511635e-21
+ ub = 6.162215032e-18 lub = -5.533080790e-25 wub = -4.571687807e-24 pub = 6.200857145e-31
+ uc = 2.991297838e-11 luc = -2.187678870e-18 wuc = 1.080658476e-16 puc = -2.818365238e-24
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.304865919e+04 lvsat = 2.575556110e-02 wvsat = 1.998716153e-01 pvsat = -3.159764134e-8
+ a0 = 1.5
+ ags = -1.311908588e+01 lags = 1.895009415e-06 wags = 1.840151118e-05 pags = -2.426809697e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.650122539e-01 lketa = -3.495008106e-08 wketa = -6.464787518e-07 pketa = 8.525826426e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.388955325e+00 lpclm = -1.645895091e-07 wpclm = -1.237665529e-06 ppclm = 1.632245676e-13
+ pdiblc1 = -1.996899662e+00 lpdiblc1 = 3.104309684e-07 wpdiblc1 = 3.014443566e-06 ppdiblc1 = -3.975478319e-13
+ pdiblc2 = -5.961288454e-02 lpdiblc2 = 8.970413296e-09 wpdiblc2 = 8.710730370e-08 ppdiblc2 = -1.148779832e-14
+ pdiblcb = -1.524525019e+00 lpdiblcb = 1.874331345e-07 wpdiblcb = 1.820071655e-06 ppdiblcb = -2.400328700e-13
+ drout = 6.303344275e+00 ldrout = -7.649121231e-07 wdrout = -7.427688159e-06 pdrout = 9.795709421e-13
+ pscbe1 = 8.916162125e+08 lpscbe1 = -1.321399253e+01 wpscbe1 = -1.283146297e+02 ppscbe1 = 1.692226168e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.829004730e-05 lalpha0 = -5.045773298e-12 walpha0 = -4.902806513e-11 palpha0 = 6.465870257e-18
+ alpha1 = 0.85
+ beta0 = 7.156919742e+01 lbeta0 = -7.628085550e-06 wbeta0 = -7.218117157e-05 pbeta0 = 9.539840908e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.412434727e-01 lkt1 = 1.586300707e-08 wkt1 = 8.017069688e-08 pkt1 = -1.057299168e-14
+ kt2 = 1.085413286e-01 lkt2 = -1.812312231e-08 wkt2 = -1.759847921e-07 pkt2 = 2.320905037e-14
+ at = -2.168541226e+05 lat = 4.464924703e-02 wat = 2.855379557e-01 pat = -5.133424485e-8
+ ute = 1.080826657e+01 lute = -1.599361740e-06 wute = -1.553062097e-05 pute = 2.048193824e-12
+ ua1 = 2.814488948e-08 lua1 = -3.714921181e-15 wua1 = -3.607378577e-14 pua1 = 4.757446941e-21
+ ub1 = -2.442216287e-17 lub1 = 3.314158457e-24 wub1 = 3.218217464e-23 pub1 = -4.244217373e-30
+ uc1 = -9.787892177e-10 luc1 = 1.484947707e-16 wuc1 = 1.441960215e-15 puc1 = -1.901671551e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.53 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {3.612268501e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = 3.136671157e-8
+ k1 = 0.90707349
+ k2 = -1.221014082e-01 wk2 = 4.226650125e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.45862506
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 3.205620505e+00 wnfactor = -2.544494192e-7
+ eta0 = 0.00069413878
+ etab = -0.043998
+ u0 = 2.774465211e-02 wu0 = -4.544517445e-9
+ ua = -1.227265464e-09 wua = 1.123632457e-16
+ ub = 1.966704845e-18 wub = 1.301700381e-25
+ uc = 1.332469903e-11 wuc = 8.669532994e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.722452884e+05 wvsat = -3.972045142e-2
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 0.0
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.14094
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 1.372852629e+01 wbeta0 = 1.555631257e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.22096074
+ kt2 = -0.028878939
+ at = 1.217029632e+05 wat = -1.037087504e-1
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.54 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {6.595471608e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.671859353e-06 wvth0 = -1.803683096e-07 pvth0 = 3.598687049e-12
+ k1 = 4.897860421e-01 lk1 = -3.246183422e-07 wk1 = 1.038878628e-07 pk1 = -2.072758275e-12
+ k2 = 2.727454267e-02 lk2 = -5.467832096e-07 wk2 = -7.956438880e-08 pk2 = 1.587459217e-12
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-9.192806945e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -3.888482053e-07 wvoff = -1.588795016e-08 pvoff = 3.169944910e-13
+ nfactor = 4.162176543e+00 lnfactor = -3.054845554e-05 wnfactor = -1.372248782e-06 pnfactor = 2.737894440e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 5.323357313e-02 lu0 = -4.828629167e-07 wu0 = -2.891030721e-08 pu0 = 5.768150092e-13
+ ua = 1.024091129e-09 lua = -3.359717951e-14 wua = -2.219955467e-15 pua = 4.429228731e-20
+ ub = 3.707087092e-19 lub = 2.267513899e-23 wub = 1.574116577e-24 pub = -3.140658663e-29
+ uc = 1.922710631e-10 luc = -3.321430793e-15 wuc = -1.409117605e-16 puc = 2.811454676e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.684286442e+00 la0 = -6.089582276e-06 wa0 = -3.325165817e-07 pa0 = 6.634331269e-12
+ ags = 8.618832808e-01 lags = -1.062342454e-05 wags = -5.237376406e-07 pags = 1.044955108e-11
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -4.486854253e-07 lb0 = 8.952118211e-12 wb0 = 5.746009135e-13 pb0 = -1.146436905e-17
+ b1 = -7.895301885e-09 lb1 = 1.575261237e-13 wb1 = 1.011097624e-14 pb1 = -2.017329948e-19
+ keta = -1.213695165e-02 lketa = 2.115616446e-07 wketa = 6.979952726e-09 pketa = -1.392631862e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.104469165e-01 lpclm = -6.522587463e-06 wpclm = -4.186589840e-07 ppclm = 8.353034228e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 9.658615594e-03 lpdiblc2 = -1.298516877e-07 wpdiblc2 = -9.435214315e-09 ppdiblc2 = 1.882502732e-13
+ pdiblcb = -1.478037615e+01 lpdiblcb = 2.506320366e-04 wpdiblcb = 1.561816460e-05 ppdiblcb = -3.116117615e-10
+ drout = 0.56
+ pscbe1 = 3.589796013e+09 lpscbe1 = -5.642955015e+04 wpscbe1 = -3.570784908e+03 ppscbe1 = 7.124387557e-2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.692301717e-01 lkt1 = 3.526498393e-06 wkt1 = 1.881754555e-07 pkt1 = -3.754454295e-12
+ kt2 = -1.027721283e-01 lkt2 = 1.638757208e-06 wkt2 = 7.250490117e-08 pkt2 = -1.446609160e-12
+ at = -3.165832151e+04 lat = 3.424906403e+00 wat = 2.198311396e-01 pat = -4.386044737e-6
+ ute = -5.225710583e+00 lute = 7.857071854e-05 wute = 4.238972460e-06 pute = -8.457547409e-11
+ ua1 = -3.799346932e-09 lua1 = 1.028109840e-13 wua1 = 4.962656572e-15 pua1 = -9.901433336e-20
+ ub1 = 4.115258733e-19 lub1 = -2.700658427e-23 wub1 = -9.063951930e-25 pub1 = 1.808428903e-29
+ uc1 = -6.643697292e-11 luc1 = 8.385506217e-16 wuc1 = 1.171450623e-16 puc1 = -2.337264342e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.55 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {0.525632+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.47351598
+ k2 = -0.0001305531
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.11141737+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 2.63107
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0290322
+ ua = -6.5981925e-10
+ ub = 1.5072e-18
+ uc = 2.5799e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.379073
+ ags = 0.329431
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.0015333577
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.083531
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0031503727
+ pdiblcb = -2.2185512
+ drout = 0.56
+ pscbe1 = 761513800.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.29248
+ kt2 = -0.020636654
+ at = 140000.0
+ ute = -1.2877
+ ua1 = 1.3536e-9
+ ub1 = -9.4206e-19
+ uc1 = -2.4408323e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.56 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.261329009e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.983104483e-9
+ k1 = 4.569800848e-01 lk1 = 1.314914708e-7
+ k2 = 7.632929869e-03 lk2 = -6.173429272e-08 wk2 = -8.673617380e-25 pk2 = -2.775557562e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.167594931e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 4.247992715e-8
+ nfactor = 2.386320130e+00 lnfactor = 1.946221841e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.997561279e-02 lu0 = -7.501906254e-9
+ ua = -6.233902280e-10 lua = -2.896792476e-16
+ ub = 1.507555669e-18 lub = -2.828239869e-27
+ uc = 2.621592345e-11 luc = -3.315325625e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.495909374e+00 la0 = -9.290689409e-7
+ ags = 3.392148694e-01 lags = -7.780016508e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.269093046e-02 lketa = 8.872369085e-08 wketa = -1.734723476e-24 pketa = -2.081668171e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.606890755e-01 lpclm = 3.532385178e-06 wpclm = -1.110223025e-22
+ pdiblc1 = 0.39
+ pdiblc2 = 2.958440708e-03 lpdiblc2 = 1.526220364e-9
+ pdiblcb = -4.385714527e+00 lpdiblcb = 1.723302489e-5
+ drout = 0.56
+ pscbe1 = 7.776031919e+08 lpscbe1 = -1.279409298e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.912647966e-01 lkt1 = -9.663152887e-9
+ kt2 = -2.057567252e-02 lkt2 = -4.849174381e-10
+ at = 140000.0
+ ute = -1.487467585e+00 lute = 1.588528060e-6
+ ua1 = 1.252925832e-09 lua1 = 8.005490075e-16
+ ub1 = -9.359247047e-19 lub1 = -4.878713775e-26
+ uc1 = -3.045817068e-11 luc1 = 4.810766883e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.57 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.074546213e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.983123382e-8
+ k1 = 4.422672016e-01 lk1 = 1.896350346e-7
+ k2 = 1.464013110e-02 lk2 = -8.942591814e-08 pk2 = 2.775557562e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-8.664948260e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.651125123e-8
+ nfactor = 3.260621691e+00 lnfactor = -1.508913887e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.897131030e-02 lu0 = -3.533022299e-9
+ ua = -2.470893049e-10 lua = -1.776775716e-15
+ ub = 9.417411723e-19 lub = 2.233203320e-24
+ uc = -2.649083338e-12 luc = 1.107557462e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.372621647e+00 la0 = -4.418505176e-7
+ ags = 2.060309996e-01 lags = 4.485266396e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.791565865e-02 lketa = -7.174871712e-08 pketa = -2.775557562e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.098057438e-01 lpclm = 9.229324121e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 1.439337851e-03 lpdiblc2 = 7.529534081e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.917747749e+08 lpscbe1 = 2.112427606e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.956911592e-01 lkt1 = 7.829305460e-9
+ kt2 = -2.362580522e-02 lkt2 = 1.156884401e-8
+ at = 1.681070864e+05 lat = -1.110758607e-1
+ ute = -1.732577830e+00 lute = 2.557174581e-6
+ ua1 = -6.478469656e-10 lua1 = 8.312176910e-15
+ ub1 = 7.966432982e-19 lub1 = -6.895689710e-24 pub1 = -3.081487911e-45
+ uc1 = -6.637324182e-12 luc1 = -4.602948185e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.58 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.179855929e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.927603051e-8
+ k1 = 5.966824121e-01 lk1 = -1.117650811e-7
+ k2 = -4.957004899e-02 lk2 = 3.590471238e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.455643000e-01 ldsub = -5.573875314e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.015830594e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -4.736268633e-8
+ nfactor = 2.885647174e+00 lnfactor = -7.770082518e-7
+ eta0 = 1.537409836e-01 leta0 = -1.439336249e-7
+ etab = -5.631671062e-02 letab = -2.670815255e-8
+ u0 = 2.873101599e-02 lu0 = -3.063996420e-9
+ ua = -9.365879010e-10 lua = -4.309565068e-16
+ ub = 1.973747937e-18 lub = 2.188489244e-25
+ uc = 3.881630995e-11 luc = 2.982023293e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.048119000e+04 lvsat = 1.857958438e-2
+ a0 = 1.458514562e+00 la0 = -6.095032656e-7
+ ags = 3.405996804e-01 lags = 1.858645883e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.634123739e-02 lketa = 3.415428738e-08 wketa = -1.387778781e-23 pketa = -1.387778781e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.321841752e-01 lpclm = 2.438013063e-7
+ pdiblc1 = 4.388270976e-01 lpdiblc1 = -9.530468411e-08 wpdiblc1 = -4.440892099e-22
+ pdiblc2 = 4.811682871e-03 lpdiblc2 = 9.471179099e-10
+ pdiblcb = -1.800242252e-03 lpdiblcb = -4.528316635e-8
+ drout = 7.148712196e-01 ldrout = -3.022901909e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.114225720e-08 lalpha0 = -2.229550126e-15
+ alpha1 = 9.956377930e-01 lalpha1 = -2.842676410e-7
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.250339102e-01 lkt1 = 6.510286367e-8
+ kt2 = -6.229275676e-05 lkt2 = -3.442432826e-8
+ at = 1.354586873e+05 lat = -4.735007080e-2
+ ute = 1.718178647e-01 lute = -1.159979192e-6
+ ua1 = 5.861327436e-09 lua1 = -4.392956931e-15
+ ub1 = -4.609958711e-18 lub1 = 3.657354026e-24 wub1 = -3.081487911e-39
+ uc1 = -7.616316627e-11 luc1 = 8.967668832e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.59 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.733778153e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.450773586e-9
+ k1 = 4.031517729e-01 lk1 = 7.245305732e-8
+ k2 = 8.603374070e-03 lk2 = -1.946946373e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.117788567e-01 ldsub = 4.590079015e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.566723314e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 5.075744911e-9
+ nfactor = 9.819304253e-01 lnfactor = 1.035103551e-6
+ eta0 = -4.380243872e-01 leta0 = 4.193565881e-07 weta0 = -7.979727989e-23 peta0 = 3.469446952e-29
+ etab = -1.603474931e-01 letab = 7.231677273e-8
+ u0 = 2.862742473e-02 lu0 = -2.965389860e-9
+ ua = -1.306434138e-09 lua = -7.890690076e-17
+ ub = 2.327364231e-18 lub = -1.177517074e-25
+ uc = 6.345977625e-11 luc = 6.362585589e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.381723763e+04 lvsat = 1.540406403e-2
+ a0 = 2.020150684e-01 la0 = 5.865347289e-7
+ ags = 3.034976292e-02 lags = 4.811855900e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 4.675999412e-02 lketa = -3.542938598e-08 wketa = 1.387778781e-23 pketa = 6.938893904e-30
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 8.584974222e-01 lpclm = -1.619981737e-7
+ pdiblc1 = 5.163711879e-01 lpdiblc1 = -1.691174303e-7
+ pdiblc2 = 9.603259256e-03 lpdiblc2 = -3.613892611e-9
+ pdiblcb = -7.139951550e-02 lpdiblcb = 2.096705946e-08 wpdiblcb = 5.551115123e-23
+ drout = -1.473977191e-01 ldrout = 5.184872287e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.771548560e-08 lalpha0 = 1.032328652e-15
+ alpha1 = 5.587244140e-01 lalpha1 = 1.316219031e-7
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.438766302e-01 lkt1 = -1.214920922e-8
+ kt2 = -3.611529325e-02 lkt2 = -1.061620977e-10
+ at = 1.178750201e+05 lat = -3.061251210e-2
+ ute = -8.848952854e-01 lute = -1.541140217e-7
+ ua1 = 1.384291714e-09 lua1 = -1.313516911e-16
+ ub1 = -8.472332519e-19 lub1 = 7.568715372e-26
+ uc1 = -1.072283955e-12 luc1 = 1.819910418e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.60 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {6.194209830e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.425680624e-8
+ k1 = 2.860351215e-01 lk1 = 1.253758469e-7
+ k2 = 4.468490015e-02 lk2 = -3.577401981e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.960437946e-01 ldsub = 5.301116574e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.103590352e-03 lcdscd = -1.221701112e-9
+ cit = 0.0
+ voff = {-1.187591359e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.205650776e-8
+ nfactor = 3.672298352e+00 lnfactor = -1.806225979e-7
+ eta0 = 8.851262253e-01 leta0 = -1.785500338e-7
+ etab = 3.496458970e-02 letab = -1.594104657e-08 wetab = -4.770489559e-24 petab = -5.095750211e-30
+ u0 = 1.661092140e-02 lu0 = 2.464639680e-9
+ ua = -1.722286886e-09 lua = 1.090090550e-16 wua = 1.654361225e-30
+ ub = 1.918798574e-18 lub = 6.687135026e-26
+ uc = 6.541098952e-11 luc = 5.480869385e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.329428353e+04 lvsat = 1.112156705e-2
+ a0 = 1.5
+ ags = 9.701952848e-01 lags = 5.648725571e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 9.946273253e-03 lketa = -1.879396498e-08 pketa = -6.938893904e-30
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 7.111109993e-01 lpclm = -9.539704948e-8
+ pdiblc1 = -3.137998472e-02 lpdiblc1 = 7.840091731e-8
+ pdiblc2 = -3.885586127e-03 lpdiblc2 = 2.481460330e-9
+ pdiblcb = 3.822571337e-02 lpdiblcb = -2.857049858e-08 ppdiblcb = 6.938893904e-30
+ drout = 1.401075642e+00 ldrout = -1.812384623e-7
+ pscbe1 = 8.069286528e+08 lpscbe1 = -3.130926566e+0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.678320160e-08 lalpha0 = -3.065199922e-15
+ alpha1 = 0.85
+ beta0 = 1.348853896e+01 lbeta0 = 1.678561862e-07 wbeta0 = 1.421085472e-20
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.948281184e-01 lkt1 = 1.087480021e-8
+ kt2 = -4.238347137e-02 lkt2 = 2.726308500e-9
+ at = 6.741939690e+04 lat = -7.812574629e-3
+ ute = -1.150766511e+00 lute = -3.397186617e-8
+ ua1 = 1.995991029e-09 lua1 = -4.077669889e-16
+ ub1 = -1.800173492e-18 lub1 = 5.063027425e-25
+ uc1 = -4.799819162e-11 luc1 = 3.940403026e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.61 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {1.111546436e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.236075849e-07 wvth0 = -5.101465013e-07 pvth0 = 1.029888858e-13
+ k1 = 0.90707349
+ k2 = -3.911422109e-01 lk2 = 5.221119318e-08 wk2 = 2.264371192e-07 pk2 = -4.571335207e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586393070e-01 ldsub = -1.878912639e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {-1.237493850e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.104907129e-8
+ nfactor = -4.684159752e+00 lnfactor = 1.506387520e-06 wnfactor = 9.002457177e-06 pnfactor = -1.817425057e-12
+ eta0 = 6.941422985e-04 leta0 = -4.640229594e-16
+ etab = -0.043998
+ u0 = 5.480530824e-02 lu0 = -5.246081330e-09 wu0 = -2.212374380e-08 pu0 = 4.466363522e-15
+ ua = -1.493330234e-09 lua = 6.278705698e-17 wua = 2.950369207e-16 pua = -5.956234859e-23
+ ub = 4.009202378e-18 lub = -3.551414601e-25 wub = -1.814470906e-24 pub = 3.663072010e-31
+ uc = 3.300159011e-10 luc = -4.793783477e-17 wuc = -2.762555585e-16 puc = 5.577074841e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.801864384e+05 lvsat = -8.439118071e-03 wvsat = -6.039775428e-02 pvsat = 1.219315903e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.282328101e-01 lketa = 8.985416655e-08 wketa = 3.693762611e-07 pketa = -7.457004896e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.390826769e-01 lpclm = -2.029159973e-08 wpclm = 1.068349801e-07 ppclm = -2.156795262e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.634970560e-08 lalpha0 = 1.573656452e-14 walpha0 = 7.955796392e-14 palpha0 = -1.606124131e-20
+ alpha1 = 0.85
+ beta0 = 1.690650061e+01 lbeta0 = -5.221653288e-07 wbeta0 = -2.178372822e-06 pbeta0 = 4.397720836e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.265552771e-01 lkt1 = 3.746801075e-08 wkt1 = 1.894237236e-07 pkt1 = -3.824105075e-14
+ kt2 = -0.028878939
+ at = 1.540265670e+05 lat = -2.529691673e-02 wat = -1.894237236e-01 pat = 3.824105075e-8
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.62 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {-5.784099618e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.926555485e-08 wvth0 = 1.234695681e-06 pvth0 = -1.271226460e-13
+ k1 = 0.90707349
+ k2 = 3.004923798e-01 lk2 = -3.900226827e-08 wk2 = -4.989206267e-07 pk2 = 4.994755282e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.45862506
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 2.607607110e+01 lnfactor = -2.550302484e-06 wnfactor = -2.954308030e-05 pnfactor = 3.265998971e-12
+ eta0 = 0.00069413878
+ etab = -0.043998
+ u0 = -1.826148739e-02 lu0 = 4.390040744e-09 wu0 = 5.437241699e-08 pu0 = -5.622026659e-15
+ ua = -7.048125619e-10 lua = -4.120344209e-17 wua = -5.567066590e-16 pua = 5.276644644e-23
+ ub = -1.932200094e-18 lub = 4.284166394e-25 wub = 5.123232468e-24 pub = -5.486440577e-31
+ uc = -4.223203366e-10 luc = 5.128102060e-17 wuc = 6.445963032e-16 puc = -6.567211597e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.001453269e+05 lvsat = 2.116783763e-03 wvsat = 5.261306650e-02 pvsat = -2.710821024e-9
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.730098440e-01 lketa = -6.856691591e-08 wketa = -8.618779425e-07 pketa = 8.780898666e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.852197268e-01 wpclm = -5.670603505e-8
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.749559664e-07 lalpha0 = -1.476825881e-14 walpha0 = -1.856352492e-13 palpha0 = 1.891270482e-20
+ alpha1 = 0.85
+ beta0 = 9.880967587e+00 lbeta0 = 4.043689913e-07 wbeta0 = 5.082869917e-06 pbeta0 = -5.178478700e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 1.241725133e-01 lkt1 = -3.516252098e-08 wkt1 = -4.419886885e-07 pkt1 = 4.503024957e-14
+ kt2 = -0.028878939
+ at = -3.044127663e+05 lat = 3.516252098e-02 wat = 4.419886885e-01 pat = -4.503024957e-8
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.63 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.368623031e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.448136835e-06 wvth0 = 4.691098210e-08 pvth0 = -4.688840901e-12
+ k1 = 7.183346898e-01 lk1 = -1.502546339e-05 wk1 = -1.293762006e-07 pk1 = 1.293139461e-11
+ k2 = -1.049588928e-01 lk2 = 6.433717352e-06 wk2 = 5.539728694e-08 pk2 = -5.537063032e-12
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.032831597e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -4.992276900e-07 wvoff = -4.298581688e-09 pvoff = 4.296513253e-13
+ nfactor = 3.018021011e+00 lnfactor = -2.374866795e-05 wnfactor = -2.044870331e-07 pnfactor = 2.043886360e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.047911880e-02 lu0 = 5.249354044e-07 wu0 = 4.519937018e-09 pu0 = -4.517762070e-13
+ ua = -1.678365121e-09 lua = 6.251206748e-14 wua = 5.382578609e-16 pua = -5.379988566e-20
+ ub = 2.348724528e-18 lub = -5.164758856e-23 wub = -4.447096642e-25 pub = 4.444956744e-29
+ uc = 8.471089878e-11 luc = -3.615649226e-15 wuc = -3.113241486e-17 puc = 3.111743425e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.336393094e+00 la0 = 2.619429576e-06 wa0 = 2.255450215e-08 pa0 = -2.254364915e-12
+ ags = 3.694578240e-01 lags = -2.456599740e-06 wags = -2.115246183e-08 pags = 2.114228348e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 2.370259543e-07 lb0 = -1.454719209e-11 wb0 = -1.252580632e-13 pb0 = 1.251977903e-17
+ b1 = 4.170831852e-09 lb1 = -2.559799509e-13 wb1 = -2.204105965e-15 pb1 = 2.203045371e-19
+ keta = -9.340369107e-03 lketa = 4.791462394e-07 wketa = 4.125671095e-09 pketa = -4.123685863e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -8.916807315e-02 lpclm = 1.059920463e-05 wpclm = 9.126406213e-08 ppclm = -9.122014677e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -2.523816917e-03 lpdiblc2 = 3.482467841e-07 wpdiblc2 = 2.998566143e-09 ppdiblc2 = -2.997123263e-13
+ pdiblcb = 3.464722011e+00 lpdiblcb = -3.488042791e-04 wpdiblcb = -3.003366434e-06 ppdiblcb = 3.001921244e-10
+ drout = 0.56
+ pscbe1 = -6.285401485e+08 lpscbe1 = 8.531294335e+04 wpscbe1 = 7.345839651e+02 ppscbe1 = -7.342304906e-2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.766755061e-01 lkt1 = -9.699824207e-07 wkt1 = -8.351998004e-09 pkt1 = 8.347979107e-13
+ kt2 = -4.364716027e-02 lkt2 = 1.412243043e-06 wkt2 = 1.216006685e-08 pkt2 = -1.215421555e-12
+ at = 2.306815224e+05 lat = -5.565472905e+00 wat = -4.792130003e-02 pat = 4.789824078e-6
+ ute = -8.412878195e-01 lute = -2.739802805e-05 wute = -2.359097141e-07 pute = 2.357961967e-11
+ ua1 = 7.509565108e-10 lua1 = 3.698654279e-14 wua1 = 3.184712682e-16 pua1 = -3.183180230e-20
+ ub1 = 2.328366995e-20 lub1 = -5.924684428e-23 wub1 = -5.101427765e-25 pub1 = 5.098973009e-29
+ uc1 = 1.264512325e-10 luc1 = -9.258829650e-15 wuc1 = -7.972281261e-17 puc1 = 7.968445079e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.64 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {8.320498673e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.436598417e-06 wvth0 = -3.127398807e-07 pvth0 = 2.486870315e-12
+ k1 = -3.715564891e-01 lk1 = 6.719915711e-06 wk1 = 8.625080043e-07 pk1 = -6.858561012e-12
+ k2 = 3.617190129e-01 lk2 = -2.877384689e-06 wk2 = -3.693152463e-07 pk2 = 2.936750890e-12
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.394952779e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.232721820e-07 wvoff = 2.865721125e-08 pvoff = -2.278787337e-13
+ nfactor = 1.295381047e+00 lnfactor = 1.062123961e-05 wnfactor = 1.363246887e-06 pnfactor = -1.084037702e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 5.855597885e-02 lu0 = -2.347695761e-07 wu0 = -3.013291346e-08 pu0 = 2.396133420e-13
+ ua = 2.856027538e-09 lua = -2.795759528e-14 wua = -3.588385739e-15 pua = 2.853441638e-20
+ ub = -1.397599276e-18 lub = 2.309861817e-23 wub = 2.964731095e-24 pub = -2.357518886e-29
+ uc = -1.775548360e-10 luc = 1.617045505e-15 wuc = 2.075494324e-16 puc = -1.650408388e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.526396764e+00 la0 = -1.171501038e-06 wa0 = -1.503633477e-07 pa0 = 1.195671448e-12
+ ags = 1.912652241e-01 lags = 1.098677808e-06 wags = 1.410164122e-07 pags = -1.121345729e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -8.181732050e-07 lb0 = 6.506015964e-12 wb0 = 8.350537546e-13 pb0 = -6.640248085e-18
+ b1 = -1.439700085e-08 lb1 = 1.144832375e-13 wb1 = 1.469403977e-14 pb1 = -1.168452556e-19
+ keta = 2.541511537e-02 lketa = -2.142910510e-07 wketa = -2.750447396e-08 pketa = 2.187123039e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.796587727e-01 lpclm = -4.740337109e-06 wpclm = -6.084270809e-07 ppclm = 4.838139744e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 2.273670838e-02 lpdiblc2 = -1.557482105e-07 wpdiblc2 = -1.999044096e-08 ppdiblc2 = 1.589616076e-13
+ pdiblcb = -2.183624190e+01 lpdiblcb = 1.559975419e-04 wpdiblcb = 2.002244289e-05 ppdiblcb = -1.592160832e-10
+ drout = 0.56
+ pscbe1 = 5.559743166e+09 lpscbe1 = -3.815494893e+04 wpscbe1 = -4.897226434e+03 ppscbe1 = 3.894216183e-2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.470344199e-01 lkt1 = 4.338102551e-07 wkt1 = 5.567998670e-08 pkt1 = -4.427606283e-13
+ kt2 = 5.879169268e-02 lkt2 = -6.316047608e-07 wkt2 = -8.106711233e-08 pkt2 = 6.446360303e-13
+ at = -1.730171634e+05 lat = 2.489075234e+00 wat = 3.194753335e-01 pat = -2.540429834e-6
+ ute = -2.828638779e+00 lute = 1.225336180e-05 wute = 1.572731428e-06 pute = -1.250617316e-11
+ ua1 = 3.433822634e-09 lua1 = -1.654168284e-14 wua1 = -2.123141788e-15 pua1 = 1.688297084e-20
+ ub1 = -4.274261854e-18 lub1 = 2.649727261e-23 wub1 = 3.400951843e-24 pub1 = -2.704396434e-29
+ uc1 = -5.451498022e-10 luc1 = 4.140874274e-15 wuc1 = 5.314854174e-16 puc1 = -4.226308792e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.65 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.261329009e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.983104483e-9
+ k1 = 4.569800848e-01 lk1 = 1.314914708e-7
+ k2 = 7.632929869e-03 lk2 = -6.173429272e-08 wk2 = -1.734723476e-24 pk2 = -7.806255642e-30
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.167594931e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 4.247992715e-8
+ nfactor = 2.386320130e+00 lnfactor = 1.946221841e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.997561279e-02 lu0 = -7.501906254e-9
+ ua = -6.233902280e-10 lua = -2.896792476e-16
+ ub = 1.507555669e-18 lub = -2.828239869e-27
+ uc = 2.621592345e-11 luc = -3.315325625e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.495909374e+00 la0 = -9.290689409e-07 wa0 = 1.776356839e-21
+ ags = 3.392148694e-01 lags = -7.780016508e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.269093046e-02 lketa = 8.872369085e-08 pketa = 2.775557562e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.606890755e-01 lpclm = 3.532385178e-06 wpclm = -1.110223025e-22 ppclm = -4.440892099e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 2.958440708e-03 lpdiblc2 = 1.526220364e-9
+ pdiblcb = -4.385714527e+00 lpdiblcb = 1.723302489e-5
+ drout = 0.56
+ pscbe1 = 7.776031919e+08 lpscbe1 = -1.279409298e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.912647966e-01 lkt1 = -9.663152887e-9
+ kt2 = -2.057567252e-02 lkt2 = -4.849174381e-10
+ at = 140000.0
+ ute = -1.487467585e+00 lute = 1.588528060e-6
+ ua1 = 1.252925832e-09 lua1 = 8.005490075e-16
+ ub1 = -9.359247047e-19 lub1 = -4.878713775e-26
+ uc1 = -3.045817068e-11 luc1 = 4.810766883e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.66 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.074546213e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.983123382e-8
+ k1 = 4.422672016e-01 lk1 = 1.896350346e-7
+ k2 = 1.464013110e-02 lk2 = -8.942591814e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-8.664948260e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.651125123e-8
+ nfactor = 3.260621691e+00 lnfactor = -1.508913887e-06 wnfactor = 3.552713679e-21
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.897131030e-02 lu0 = -3.533022299e-9
+ ua = -2.470893049e-10 lua = -1.776775716e-15
+ ub = 9.417411723e-19 lub = 2.233203320e-24
+ uc = -2.649083339e-12 luc = 1.107557462e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.372621647e+00 la0 = -4.418505176e-7
+ ags = 2.060309996e-01 lags = 4.485266396e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.791565865e-02 lketa = -7.174871712e-08 wketa = 1.387778781e-23
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.098057438e-01 lpclm = 9.229324121e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 1.439337851e-03 lpdiblc2 = 7.529534081e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.917747749e+08 lpscbe1 = 2.112427606e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.956911592e-01 lkt1 = 7.829305460e-9
+ kt2 = -2.362580522e-02 lkt2 = 1.156884401e-8
+ at = 1.681070864e+05 lat = -1.110758607e-1
+ ute = -1.732577830e+00 lute = 2.557174581e-06 wute = -1.776356839e-21
+ ua1 = -6.478469656e-10 lua1 = 8.312176910e-15
+ ub1 = 7.966432982e-19 lub1 = -6.895689710e-24
+ uc1 = -6.637324182e-12 luc1 = -4.602948185e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.67 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.179855929e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.927603051e-8
+ k1 = 5.966824121e-01 lk1 = -1.117650811e-7
+ k2 = -4.957004899e-02 lk2 = 3.590471238e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.455643000e-01 ldsub = -5.573875314e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.015830594e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -4.736268633e-8
+ nfactor = 2.885647174e+00 lnfactor = -7.770082518e-7
+ eta0 = 1.537409836e-01 leta0 = -1.439336249e-7
+ etab = -5.631671062e-02 letab = -2.670815255e-8
+ u0 = 2.873101599e-02 lu0 = -3.063996420e-9
+ ua = -9.365879010e-10 lua = -4.309565068e-16
+ ub = 1.973747937e-18 lub = 2.188489244e-25
+ uc = 3.881630995e-11 luc = 2.982023293e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.048119000e+04 lvsat = 1.857958438e-2
+ a0 = 1.458514562e+00 la0 = -6.095032656e-07 wa0 = -1.776356839e-21
+ ags = 3.405996804e-01 lags = 1.858645883e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.634123739e-02 lketa = 3.415428738e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.321841752e-01 lpclm = 2.438013063e-7
+ pdiblc1 = 4.388270976e-01 lpdiblc1 = -9.530468411e-8
+ pdiblc2 = 4.811682871e-03 lpdiblc2 = 9.471179099e-10
+ pdiblcb = -1.800242252e-03 lpdiblcb = -4.528316635e-8
+ drout = 7.148712196e-01 ldrout = -3.022901909e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.114225720e-08 lalpha0 = -2.229550126e-15
+ alpha1 = 9.956377930e-01 lalpha1 = -2.842676410e-7
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.250339102e-01 lkt1 = 6.510286367e-8
+ kt2 = -6.229275676e-05 lkt2 = -3.442432826e-8
+ at = 1.354586873e+05 lat = -4.735007080e-2
+ ute = 1.718178647e-01 lute = -1.159979192e-6
+ ua1 = 5.861327436e-09 lua1 = -4.392956931e-15
+ ub1 = -4.609958711e-18 lub1 = 3.657354026e-24
+ uc1 = -7.616316627e-11 luc1 = 8.967668832e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.68 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.733778153e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.450773586e-9
+ k1 = 4.031517729e-01 lk1 = 7.245305732e-8
+ k2 = 8.603374070e-03 lk2 = -1.946946373e-08 pk2 = 6.938893904e-30
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.117788567e-01 ldsub = 4.590079015e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.566723314e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 5.075744911e-9
+ nfactor = 9.819304253e-01 lnfactor = 1.035103551e-6
+ eta0 = -4.380243872e-01 leta0 = 4.193565881e-07 weta0 = -1.838806885e-22 peta0 = 1.561251128e-28
+ etab = -1.603474931e-01 letab = 7.231677273e-8
+ u0 = 2.862742473e-02 lu0 = -2.965389860e-9
+ ua = -1.306434138e-09 lua = -7.890690076e-17
+ ub = 2.327364231e-18 lub = -1.177517074e-25
+ uc = 6.345977625e-11 luc = 6.362585589e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.381723763e+04 lvsat = 1.540406403e-2
+ a0 = 2.020150684e-01 la0 = 5.865347289e-7
+ ags = 3.034976292e-02 lags = 4.811855900e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 4.675999412e-02 lketa = -3.542938598e-08 wketa = -1.387778781e-23 pketa = -6.938893904e-30
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 8.584974222e-01 lpclm = -1.619981737e-7
+ pdiblc1 = 5.163711879e-01 lpdiblc1 = -1.691174303e-7
+ pdiblc2 = 9.603259256e-03 lpdiblc2 = -3.613892611e-09 wpdiblc2 = 6.938893904e-24
+ pdiblcb = -7.139951550e-02 lpdiblcb = 2.096705946e-8
+ drout = -1.473977191e-01 ldrout = 5.184872287e-07 pdrout = 2.220446049e-28
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.771548560e-08 lalpha0 = 1.032328652e-15
+ alpha1 = 5.587244140e-01 lalpha1 = 1.316219031e-7
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.438766302e-01 lkt1 = -1.214920922e-8
+ kt2 = -3.611529325e-02 lkt2 = -1.061620977e-10
+ at = 1.178750201e+05 lat = -3.061251210e-2
+ ute = -8.848952854e-01 lute = -1.541140217e-7
+ ua1 = 1.384291714e-09 lua1 = -1.313516911e-16
+ ub1 = -8.472332519e-19 lub1 = 7.568715372e-26
+ uc1 = -1.072283955e-12 luc1 = 1.819910418e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.69 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {6.194209830e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.425680624e-8
+ k1 = 2.860351215e-01 lk1 = 1.253758469e-7
+ k2 = 4.468490015e-02 lk2 = -3.577401981e-08 pk2 = -1.387778781e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.960437946e-01 ldsub = 5.301116574e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.103590352e-03 lcdscd = -1.221701112e-9
+ cit = 0.0
+ voff = {-1.187591359e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.205650776e-8
+ nfactor = 3.672298352e+00 lnfactor = -1.806225979e-7
+ eta0 = 8.851262253e-01 leta0 = -1.785500338e-7
+ etab = 3.496458970e-02 letab = -1.594104657e-08 wetab = -1.257674520e-23 petab = 2.059984128e-30
+ u0 = 1.661092140e-02 lu0 = 2.464639680e-9
+ ua = -1.722286886e-09 lua = 1.090090550e-16
+ ub = 1.918798574e-18 lub = 6.687135026e-26
+ uc = 6.541098952e-11 luc = 5.480869385e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.329428353e+04 lvsat = 1.112156705e-2
+ a0 = 1.5
+ ags = 9.701952848e-01 lags = 5.648725571e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 9.946273253e-03 lketa = -1.879396498e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 7.111109993e-01 lpclm = -9.539704948e-8
+ pdiblc1 = -3.137998472e-02 lpdiblc1 = 7.840091731e-8
+ pdiblc2 = -3.885586127e-03 lpdiblc2 = 2.481460330e-09 ppdiblc2 = 4.336808690e-31
+ pdiblcb = 3.822571337e-02 lpdiblcb = -2.857049858e-8
+ drout = 1.401075642e+00 ldrout = -1.812384623e-7
+ pscbe1 = 8.069286528e+08 lpscbe1 = -3.130926566e+00 wpscbe1 = -9.536743164e-13
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.678320160e-08 lalpha0 = -3.065199922e-15
+ alpha1 = 0.85
+ beta0 = 1.348853896e+01 lbeta0 = 1.678561862e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.948281184e-01 lkt1 = 1.087480021e-8
+ kt2 = -4.238347137e-02 lkt2 = 2.726308500e-9
+ at = 6.741939690e+04 lat = -7.812574629e-3
+ ute = -1.150766511e+00 lute = -3.397186617e-8
+ ua1 = 1.995991029e-09 lua1 = -4.077669889e-16
+ ub1 = -1.800173492e-18 lub1 = 5.063027425e-25
+ uc1 = -4.799819162e-11 luc1 = 3.940403026e-17 puc1 = -1.292469707e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.70 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {6.117125086e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.270061173e-8
+ k1 = 0.90707349
+ k2 = -1.692825012e-01 lk2 = 7.421933131e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586393070e-01 ldsub = -1.878912639e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {-1.237493850e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.104907129e-8
+ nfactor = 4.136313423e+00 lnfactor = -2.742984245e-7
+ eta0 = 6.941422985e-04 leta0 = -4.640229594e-16
+ etab = -0.043998
+ u0 = 3.312879428e-02 lu0 = -8.700050142e-10
+ ua = -1.204257462e-09 lua = 4.428756835e-18
+ ub = 2.231410867e-18 lub = 3.760868051e-27
+ uc = 5.934482814e-11 luc = 6.705512110e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.210096203e+05 lvsat = 3.507557157e-3
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.663234627e-01 lketa = 1.679154558e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.437579959e-01 lpclm = -4.142355779e-8
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.16e-8
+ alpha1 = 0.85
+ beta0 = 1.477216343e+01 lbeta0 = -9.128320512e-8
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.24096074
+ kt2 = -0.028878939
+ at = -3.156797014e+04 lat = 1.217109402e-2
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.71 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {2.095027150e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.034321807e-08 wvth0 = 4.305267901e-07 pvth0 = -5.677830361e-14
+ k1 = 0.90707349
+ k2 = -1.967637336e-01 lk2 = 1.104618554e-08 wk2 = 8.594874859e-09 pk2 = -1.133500691e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.587152994e-01 ldsub = -1.190086783e-11 wdsub = -9.210126205e-11 pdsub = 1.214640654e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = -1.969379114e+01 lnfactor = 2.868439596e-06 wnfactor = 1.717110574e-05 pnfactor = -2.264542596e-12
+ eta0 = -1.198575802e-02 leta0 = 1.672237627e-09 weta0 = 1.294150965e-08 peta0 = -1.706739234e-15
+ etab = -0.043998
+ u0 = 2.886857169e-02 lu0 = -3.081625991e-10 wu0 = 6.269970532e-09 pu0 = -8.268899837e-16
+ ua = -1.393114108e-09 lua = 2.933536017e-17 wua = 1.457959249e-16 pua = -1.922771238e-23
+ ub = 5.821356358e-18 lub = -4.696847332e-25 wub = -2.790295360e-24 pub = 3.679869424e-31
+ uc = 1.358483186e-10 luc = -3.383844714e-18 wuc = 7.491151233e-17 puc = -9.879405157e-24
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.807212357e+05 lvsat = -4.367270400e-03 wvsat = -2.962528449e-02 pvsat = 3.907012144e-9
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.042393423e-05 lb0 = -1.374718871e-12 wb0 = -1.063900085e-11 pb0 = 1.403082070e-18
+ b1 = -1.489699742e-08 lb1 = 1.964630917e-15 wb1 = 1.520435227e-14 pb1 = -2.005165182e-21
+ keta = -6.646568245e-01 lketa = 8.251224767e-08 wketa = 5.033874646e-07 pketa = -6.638724222e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.007979923e-01 lpclm = 3.806350441e-09 wpclm = 2.945748867e-08 ppclm = -3.884883063e-15
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.926680000e-09 lalpha0 = 3.762127085e-15
+ alpha1 = 0.85
+ beta0 = 1.851450637e+01 lbeta0 = -5.848271341e-07 wbeta0 = -3.728796034e-06 pbeta0 = 4.917573498e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -6.742232766e-01 lkt1 = 5.713909659e-08 wkt1 = 3.728796034e-07 pkt1 = -4.917573498e-14
+ kt2 = -0.028878939
+ at = 3.661133691e+05 lat = -4.027551869e-02 wat = -2.423717422e-01 pat = 3.196422774e-8
+ ute = -4.056885251e-01 lute = -1.204541279e-07 wute = -9.321990086e-07 pute = 1.229393374e-13
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.72 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {0.4913699+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56800772
+ k2 = -0.040590746
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 2.78042
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.025731
+ ua = -1.0529435e-9
+ ub = 1.832e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 9.1484e-8
+ b1 = 1.6098e-9
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.73 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.686658882e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.529877423e-7
+ k1 = 6.306233093e-01 lk1 = -1.249298787e-6
+ k2 = -6.740196593e-02 lk2 = 5.349342695e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.061974093e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -4.150850668e-8
+ nfactor = 2.879387786e+00 lnfactor = -1.974593481e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.354343754e-02 lu0 = 4.364598594e-8
+ ua = -1.313449938e-09 lua = 5.197593448e-15
+ ub = 2.047230912e-18 lub = -4.294261552e-24
+ uc = 6.360448918e-11 luc = -3.006247511e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.351684055e+00 la0 = 2.177936285e-7
+ ags = 3.551173841e-01 lags = -2.042550699e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.521064901e-07 lb0 = -1.209532709e-12
+ b1 = 2.676544836e-09 lb1 = -2.128356603e-14
+ keta = -6.543345349e-03 lketa = 3.983882560e-08 pketa = 5.551115123e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.729504833e-02 lpclm = 8.812755480e-07 ppclm = 2.220446049e-28
+ pdiblc1 = 0.39
+ pdiblc2 = -4.909208011e-04 lpdiblc2 = 2.895513261e-8
+ pdiblcb = 1.428571509e+00 lpdiblcb = -2.900148578e-05 wpdiblcb = -2.775557562e-22 ppdiblcb = -3.552713679e-27
+ drout = 0.56
+ pscbe1 = -1.305244910e+08 lpscbe1 = 7.093382338e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.823377938e-01 lkt1 = -8.064961658e-8
+ kt2 = -3.540316915e-02 lkt2 = 1.174215713e-7
+ at = 1.981929862e+05 lat = -4.627437017e-1
+ ute = -1.001224242e+00 lute = -2.278021137e-6
+ ua1 = 9.668660399e-10 lua1 = 3.075262429e-15
+ ub1 = -3.225707215e-19 lub1 = -4.926105023e-24
+ uc1 = 7.240266785e-11 luc1 = -7.698294787e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.74 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.261329009e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.983104483e-9
+ k1 = 4.569800848e-01 lk1 = 1.314914708e-7
+ k2 = 7.632929869e-03 lk2 = -6.173429272e-08 wk2 = -2.602085214e-24 pk2 = 6.071532166e-30
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.167594931e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 4.247992715e-8
+ nfactor = 2.386320130e+00 lnfactor = 1.946221841e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.997561279e-02 lu0 = -7.501906254e-9
+ ua = -6.233902280e-10 lua = -2.896792476e-16
+ ub = 1.507555669e-18 lub = -2.828239869e-27
+ uc = 2.621592345e-11 luc = -3.315325625e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.495909374e+00 la0 = -9.290689409e-7
+ ags = 3.392148694e-01 lags = -7.780016508e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.269093046e-02 lketa = 8.872369085e-08 wketa = 3.469446952e-24
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.606890755e-01 lpclm = 3.532385178e-06 wpclm = -2.220446049e-22 ppclm = -8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 2.958440708e-03 lpdiblc2 = 1.526220364e-9
+ pdiblcb = -4.385714527e+00 lpdiblcb = 1.723302489e-5
+ drout = 0.56
+ pscbe1 = 7.776031919e+08 lpscbe1 = -1.279409298e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.912647966e-01 lkt1 = -9.663152887e-9
+ kt2 = -2.057567252e-02 lkt2 = -4.849174381e-10
+ at = 140000.0
+ ute = -1.487467585e+00 lute = 1.588528060e-6
+ ua1 = 1.252925832e-09 lua1 = 8.005490075e-16
+ ub1 = -9.359247047e-19 lub1 = -4.878713775e-26
+ uc1 = -3.045817068e-11 luc1 = 4.810766883e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.75 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.074546213e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.983123382e-8
+ k1 = 4.422672016e-01 lk1 = 1.896350346e-7
+ k2 = 1.464013110e-02 lk2 = -8.942591814e-08 pk2 = 2.775557562e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-8.664948260e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.651125123e-8
+ nfactor = 3.260621691e+00 lnfactor = -1.508913887e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.897131030e-02 lu0 = -3.533022299e-9
+ ua = -2.470893049e-10 lua = -1.776775716e-15
+ ub = 9.417411723e-19 lub = 2.233203320e-24
+ uc = -2.649083339e-12 luc = 1.107557462e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.372621647e+00 la0 = -4.418505176e-7
+ ags = 2.060309996e-01 lags = 4.485266396e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.791565865e-02 lketa = -7.174871712e-08 pketa = 2.775557562e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.098057438e-01 lpclm = 9.229324121e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 1.439337851e-03 lpdiblc2 = 7.529534081e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.917747749e+08 lpscbe1 = 2.112427606e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.956911592e-01 lkt1 = 7.829305460e-9
+ kt2 = -2.362580522e-02 lkt2 = 1.156884401e-8
+ at = 1.681070864e+05 lat = -1.110758607e-1
+ ute = -1.732577830e+00 lute = 2.557174581e-6
+ ua1 = -6.478469656e-10 lua1 = 8.312176910e-15
+ ub1 = 7.966432982e-19 lub1 = -6.895689710e-24
+ uc1 = -6.637324182e-12 luc1 = -4.602948185e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.76 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.179855929e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.927603051e-8
+ k1 = 5.966824121e-01 lk1 = -1.117650811e-7
+ k2 = -4.957004899e-02 lk2 = 3.590471238e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.455643000e-01 ldsub = -5.573875314e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.015830594e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -4.736268633e-8
+ nfactor = 2.885647174e+00 lnfactor = -7.770082518e-07 wnfactor = 3.552713679e-21
+ eta0 = 1.537409836e-01 leta0 = -1.439336249e-7
+ etab = -5.631671062e-02 letab = -2.670815255e-8
+ u0 = 2.873101599e-02 lu0 = -3.063996420e-9
+ ua = -9.365879010e-10 lua = -4.309565068e-16
+ ub = 1.973747937e-18 lub = 2.188489244e-25
+ uc = 3.881630995e-11 luc = 2.982023293e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.048119000e+04 lvsat = 1.857958438e-2
+ a0 = 1.458514562e+00 la0 = -6.095032656e-7
+ ags = 3.405996804e-01 lags = 1.858645883e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.634123739e-02 lketa = 3.415428738e-08 wketa = 1.387778781e-23 pketa = -1.387778781e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.321841752e-01 lpclm = 2.438013063e-7
+ pdiblc1 = 4.388270976e-01 lpdiblc1 = -9.530468411e-8
+ pdiblc2 = 4.811682871e-03 lpdiblc2 = 9.471179099e-10
+ pdiblcb = -1.800242252e-03 lpdiblcb = -4.528316635e-8
+ drout = 7.148712196e-01 ldrout = -3.022901909e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.114225720e-08 lalpha0 = -2.229550126e-15
+ alpha1 = 9.956377930e-01 lalpha1 = -2.842676410e-7
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.250339102e-01 lkt1 = 6.510286367e-8
+ kt2 = -6.229275676e-05 lkt2 = -3.442432826e-8
+ at = 1.354586873e+05 lat = -4.735007080e-2
+ ute = 1.718178647e-01 lute = -1.159979192e-6
+ ua1 = 5.861327436e-09 lua1 = -4.392956931e-15
+ ub1 = -4.609958711e-18 lub1 = 3.657354026e-24
+ uc1 = -7.616316627e-11 luc1 = 8.967668832e-17 wuc1 = -5.169878828e-32 puc1 = 5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.77 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {3.129211304e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.444729961e-07 wvth0 = 2.241573576e-07 pvth0 = -2.133711297e-13
+ k1 = -2.052536689e-01 lk1 = 6.515826377e-07 wk1 = 5.236131922e-07 pk1 = -4.984174490e-13
+ k2 = 1.527060328e-01 lk2 = -1.566380466e-07 wk2 = -1.240193594e-07 pk2 = 1.180516718e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.908198630e-01 ldsub = 6.585125799e-08 wdsub = 1.803798063e-08 pdsub = -1.717001104e-14
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.442750761e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -6.724966788e-09 wvoff = -1.066947456e-08 pvoff = 1.015607011e-14
+ nfactor = -7.890653184e-01 lnfactor = 2.720880751e-06 wnfactor = 1.524175609e-06 pnfactor = -1.450833803e-12
+ eta0 = -4.380243871e-01 leta0 = 4.193565880e-07 weta0 = -1.187387758e-16 peta0 = 1.130255282e-22
+ etab = -1.624957128e-01 letab = 7.436162220e-08 wetab = 1.848826576e-09 petab = -1.759862890e-15
+ u0 = 4.493327137e-02 lu0 = -1.848661547e-08 wu0 = -1.403333341e-08 pu0 = 1.335806344e-14
+ ua = -1.085034838e-09 lua = -2.896526880e-16 wua = -1.905433225e-16 pua = 1.813745684e-22
+ ub = 2.884713468e-18 lub = -6.482818559e-25 wub = -4.796725881e-25 pub = 4.565912228e-31
+ uc = -1.084184211e-10 luc = 1.699701759e-16 wuc = 1.479238767e-16 puc = -1.408059277e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.738319570e+05 lvsat = -1.749861470e-01 wvsat = -1.721390679e-01 pvsat = 1.638559081e-7
+ a0 = -5.912794935e-01 la0 = 1.341656750e-06 wa0 = 6.827346854e-07 pa0 = -6.498821751e-13
+ ags = -6.424277010e+00 lags = 6.625222177e-06 wags = 5.555058348e-06 pags = -5.287754496e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 5.007755222e-16 lb0 = -4.766787048e-22 wb0 = -4.309834392e-22 pb0 = 4.102449471e-28
+ b1 = -2.465330662e-17 lb1 = 2.346701416e-23 wb1 = 2.121742458e-23 pb1 = -2.019646333e-29
+ keta = 2.153930525e-01 lketa = -1.959479902e-07 wketa = -1.451310063e-07 pketa = 1.381474474e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.272247601e-01 lpclm = 1.533339793e-07 wpclm = 2.851038538e-07 ppclm = -2.713849414e-13
+ pdiblc1 = -2.335276672e-01 lpdiblc1 = 5.446970418e-07 wpdiblc1 = 6.453869515e-07 ppdiblc1 = -6.143315767e-13
+ pdiblc2 = -1.116380561e-03 lpdiblc2 = 6.589928858e-09 wpdiblc2 = 9.225665055e-09 ppdiblc2 = -8.781735278e-15
+ pdiblcb = -5.498868177e-01 lpdiblcb = 4.764300311e-07 wpdiblcb = 4.118014838e-07 ppdiblcb = -3.919860082e-13
+ drout = -1.473984068e-01 ldrout = 5.184878833e-07 wdrout = 5.918148496e-13 pdrout = -5.633373101e-19
+ pscbe1 = -1.695736247e+09 lpscbe1 = 2.375643915e+03 wpscbe1 = 2.147910478e+03 ppscbe1 = -2.044555173e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.663126801e-05 lalpha0 = -2.532238385e-11 walpha0 = -2.289586861e-11 palpha0 = 2.179414231e-17
+ alpha1 = 5.587244140e-01 lalpha1 = 1.316219031e-7
+ beta0 = 4.244335176e+01 lbeta0 = -2.720794946e-05 wbeta0 = -2.459974719e-05 pbeta0 = 2.341603196e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.001571673e-01 lkt1 = 4.142316475e-08 wkt1 = 4.843683123e-08 pkt1 = -4.610609935e-14
+ kt2 = -3.864760086e-02 lkt2 = 2.304293399e-09 wkt2 = 2.179384960e-09 pkt2 = -2.074515135e-15
+ at = -1.534889695e+05 lat = 2.276937137e-01 wat = 2.335445331e-01 pat = -2.223066037e-7
+ ute = -1.464630003e+00 lute = 3.977244414e-07 wute = 4.989382498e-07 pute = -4.749298402e-13
+ ua1 = -4.163943466e-10 lua1 = 1.582687157e-15 wua1 = 1.549728046e-15 pua1 = -1.475156682e-21
+ ub1 = -5.182242992e-19 lub1 = -2.374902172e-25 wub1 = -2.831556330e-25 pub1 = 2.695304671e-31
+ uc1 = -2.310960574e-10 luc1 = 2.371543637e-16 wuc1 = 1.979658202e-16 puc1 = -1.884399029e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.78 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {9.570423974e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.659316617e-08 wvth0 = -2.905677931e-07 pvth0 = 1.922338611e-14
+ k1 = 1.502846004e+00 lk1 = -1.202751507e-07 wk1 = -1.047226384e-06 pk1 = 2.114151094e-13
+ k2 = -2.601192697e-01 lk2 = 2.990986392e-08 wk2 = 2.623242223e-07 pk2 = -5.652965222e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.379617820e-01 ldsub = 4.454872048e-08 wdsub = -3.607596137e-08 pdsub = 7.283051185e-15
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.103590344e-03 lcdscd = -1.221701108e-09 wcdscd = 6.488559690e-18 pcdscd = -2.932053905e-24
+ cit = 0.0
+ voff = {-1.435536461e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.050967303e-09 wvoff = 2.133894892e-08 pvoff = -4.307928297e-15
+ nfactor = 7.214289841e+00 lnfactor = -8.956833822e-07 wnfactor = -3.048351219e-06 pnfactor = 6.154041929e-13
+ eta0 = 8.851262253e-01 leta0 = -1.785500339e-07 weta0 = -4.801314901e-17 peta0 = 8.106582072e-23
+ etab = 3.926102897e-02 letab = -1.680841602e-08 wetab = -3.697653121e-09 petab = 7.464859019e-16
+ u0 = -1.113485300e-02 lu0 = 6.849504638e-09 wu0 = 2.387890131e-08 pu0 = -3.773755098e-15
+ ua = -2.165085484e-09 lua = 1.984016778e-16 wua = 3.810866424e-16 pua = -7.693415179e-23
+ ub = 8.041001028e-19 lub = 2.919077920e-25 wub = 9.593451749e-25 pub = -1.936735630e-31
+ uc = 4.091673843e-10 luc = -6.391701538e-17 wuc = -2.958477536e-16 puc = 5.972604036e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -3.040513344e+05 lvsat = 8.614833258e-02 wvsat = 3.333620339e-01 pvsat = -6.457043527e-8
+ a0 = 3.086589121e+00 la0 = -3.203021978e-07 wa0 = -1.365469369e-06 pa0 = 2.756623211e-13
+ ags = 1.387944883e+01 lags = -2.549645759e-06 wags = -1.111011670e-05 pags = 2.242921469e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.001551044e-15 lb0 = 2.021941264e-22 wb0 = 8.619668784e-22 pb0 = -1.740147354e-28
+ b1 = 4.930661323e-17 lb1 = -9.954068386e-24 wb1 = -4.243484916e-23 pb1 = 8.566789784e-30
+ keta = -3.273198435e-01 lketa = 4.929365591e-08 wketa = 2.902620126e-07 pketa = -5.859838534e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.373656324e+00 lpclm = -2.291523623e-07 wpclm = -5.702077079e-07 ppclm = 1.151141023e-13
+ pdiblc1 = 1.468417726e+00 lpdiblc1 = -2.243797444e-07 wpdiblc1 = -1.290773903e-06 ppdiblc1 = 2.605827265e-13
+ pdiblc2 = 1.755369350e-02 lpdiblc2 = -1.846722877e-09 wpdiblc2 = -1.845133010e-08 ppdiblc2 = 3.724972969e-15
+ pdiblcb = 9.952003177e-01 lpdiblcb = -2.217654887e-07 wpdiblcb = -8.236029677e-07 ppdiblcb = 1.662697907e-13
+ drout = 1.401077015e+00 ldrout = -1.812387389e-07 wdrout = -1.181649807e-12 pdrout = 2.380576722e-19
+ pscbe1 = 5.798401147e+09 lpscbe1 = -1.010814385e+03 wpscbe1 = -4.295820955e+03 ppscbe1 = 8.672446302e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.317032184e-05 lalpha0 = 1.073843837e-11 walpha0 = 4.579173722e-11 palpha0 = -9.244481702e-18
+ alpha1 = 0.85
+ beta0 = -4.367816456e+01 lbeta0 = 1.170872746e-05 wbeta0 = 4.919949439e-05 pbeta0 = -9.932443126e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.822670442e-01 lkt1 = -1.184914199e-08 wkt1 = -9.687366240e-08 pkt1 = 1.955695182e-14
+ kt2 = -3.731885617e-02 lkt2 = 1.703858922e-09 wkt2 = -4.358769908e-09 pkt2 = 8.799528249e-16
+ at = 6.101473761e+05 lat = -1.173790418e-01 wat = -4.670890662e-01 pat = 9.429640778e-8
+ ute = 8.702924697e-03 lute = -2.680467154e-07 wute = -9.978764997e-07 pute = 2.014523057e-13
+ ua1 = 5.597363148e-09 lua1 = -1.134815593e-15 wua1 = -3.099456090e-15 pua1 = 6.257212943e-22
+ ub1 = -2.458191401e-18 lub1 = 6.391440569e-25 wub1 = 5.663112691e-25 pub1 = -1.143274861e-31
+ uc1 = 4.120493553e-10 luc1 = -5.347082858e-17 wuc1 = -3.959316404e-16 puc1 = 7.993107551e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.79 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {6.013083237e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.522278438e-08 wvth0 = 8.954174513e-09 pvth0 = -4.124440824e-14
+ k1 = 9.070734930e-01 lk1 = -3.911853064e-16 wk1 = -2.552805967e-15 pk1 = 3.366666945e-22
+ k2 = -2.311582554e-01 lk2 = 2.406318540e-08 wk2 = 5.325225416e-08 pk2 = -1.432199422e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.587100988e-01 ldsub = -1.617046413e-11 wdsub = -6.092569117e-11 pdsub = 1.229976654e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000030e-03 lcdscd = -4.139417108e-18 wcdscd = -2.568172758e-17 pcdscd = 3.562514866e-24
+ cit = 0.0
+ voff = {-1.237493862e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.104907110e-08 wvoff = 1.034837105e-15 pvoff = -1.594769317e-22
+ nfactor = 1.670233163e+01 lnfactor = -2.811138747e-06 wnfactor = -1.081471738e-05 pnfactor = 2.183285961e-12
+ eta0 = -9.253153176e-03 leta0 = 2.008169411e-09 weta0 = 8.560960799e-09 peta0 = -1.728295256e-15
+ etab = -4.399799987e-02 letab = -1.689043350e-17 wetab = -1.102238301e-16 petab = 1.453642762e-23
+ u0 = 6.307564147e-02 lu0 = -8.132184197e-09 wu0 = -2.577321500e-08 pu0 = 6.250063795e-15
+ ua = -1.053281450e-09 lua = -2.605043222e-17 wua = -1.299347872e-16 pua = 2.623136543e-23
+ ub = 3.204175574e-18 lub = -1.926218441e-25 wub = -8.371924353e-25 pub = 1.690132463e-31
+ uc = -4.162243428e-10 luc = 1.027138919e-16 wuc = 4.092900467e-16 puc = -8.262788390e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.332879165e+04 lvsat = 1.803769534e-02 wvsat = 7.546092689e-02 pvsat = -1.250510189e-8
+ a0 = 1.500000009e+00 la0 = -1.194998767e-15 wa0 = -7.798348634e-15 pa0 = 1.028454211e-21
+ ags = 1.250000002e+00 lags = -2.558593337e-16 wags = -1.669697269e-15 pags = 2.202016347e-22
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 5.247153303e-07 lb0 = -1.059300556e-13 wb0 = -4.515868041e-13 pb0 = 9.116679560e-20
+ b1 = -7.498791184e-10 lb1 = 1.513863463e-16 wb1 = 6.453699654e-16 pb1 = -1.302879340e-22
+ keta = 5.641523391e-03 lketa = -1.792491779e-08 wketa = -1.479985699e-07 pketa = 2.987809930e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.157239903e+00 lpclm = -1.854619987e-07 wpclm = -6.140453605e-07 ppclm = 1.239640915e-13
+ pdiblc1 = 3.569721484e-01 lpdiblc1 = 2.045812408e-16 wpdiblc1 = 1.335060063e-15 ppdiblc1 = -1.760690482e-22
+ pdiblc2 = 8.406112142e-03 lpdiblc2 = -5.485285837e-18 wpdiblc2 = -3.579600505e-17 ppdiblc2 = 4.720814017e-24
+ pdiblcb = -1.032957699e-01 lpdiblcb = -1.624156365e-17 wpdiblcb = -1.059894394e-16 ppdiblcb = 1.397798544e-23
+ drout = 5.033266682e-01 ldrout = -1.083547252e-15 wdrout = -7.071037089e-15 pdrout = 9.325353822e-22
+ pscbe1 = 7.914198808e+08 lpscbe1 = -1.070451736e-07 wpscbe1 = -6.985588074e-07 ppscbe1 = 9.212660789e-14
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.419754858e-07 lalpha0 = -2.430152379e-14 walpha0 = -1.035989951e-13 palpha0 = 2.091466902e-20
+ alpha1 = 0.85
+ beta0 = 1.166438150e+01 lbeta0 = 5.361189194e-07 wbeta0 = 2.674656580e-06 pbeta0 = -5.399623452e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.070672635e-01 lkt1 = -2.703054890e-08 wkt1 = -1.152330104e-07 pkt1 = 2.326335536e-14
+ kt2 = -2.887893895e-02 lkt2 = -6.492847926e-18 wkt2 = -4.237121765e-17 pkt2 = 5.587946772e-24
+ at = -1.318808792e+05 lat = 3.242236440e-02 wat = 8.633249952e-02 pat = -1.742889134e-8
+ ute = -1.271989799e+00 lute = -9.499187629e-09 wute = -4.049566240e-08 pute = 8.175304847e-15
+ ua1 = -2.384732671e-11 lua1 = -1.225091633e-24 wua1 = -7.994730554e-24 pua1 = 1.054353063e-30
+ ub1 = 7.077531832e-19 lub1 = -1.740301883e-33 wub1 = -1.135690073e-32 pub1 = 1.497759125e-39
+ uc1 = 1.471862498e-10 luc1 = 2.519829960e-26 wuc1 = 1.644401971e-25 puc1 = -2.168650431e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.80 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {2.245797326e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.916540697e-07 wvth0 = -1.321973514e-06 pvth0 = 1.342796662e-13
+ k1 = 0.90707349
+ k2 = 5.578684387e-02 lk2 = -1.377942124e-08 wk2 = -2.087582337e-07 pk2 = 2.023221093e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.584431017e-01 ldsub = 1.904138854e-11 wdsub = 1.421608489e-10 pdsub = -1.448348944e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999994e-03 lcdscd = 6.485593312e-19 wcdscd = 5.563750849e-18 pcdscd = -5.581706972e-25
+ cit = 0.0
+ voff = {-2.075299991e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -9.076372987e-17 wvoff = -7.667200208e-16 pvoff = 7.811418179e-23
+ nfactor = -2.489978150e+01 lnfactor = 2.675389535e-06 wnfactor = 2.165154763e-05 pnfactor = -2.098397536e-12
+ eta0 = 2.626181318e-02 leta0 = -2.675579521e-09 weta0 = -1.997557282e-08 peta0 = 2.035131334e-15
+ etab = -0.043998
+ u0 = -4.640795805e-02 lu0 = 6.306622391e-09 wu0 = 7.105536087e-08 pu0 = -6.519785619e-15
+ ua = -1.636886090e-09 lua = 5.091593125e-17 wua = 3.555938929e-16 pua = -3.780064243e-23
+ ub = 2.250052681e-18 lub = -6.679116293e-26 wub = 2.832828653e-25 pub = 2.124384321e-32
+ uc = 1.332552160e-09 luc = -1.279165021e-16 wuc = -9.550101082e-16 puc = 9.729738484e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.270108485e+04 lvsat = 1.152642794e-02 wvsat = 5.473399398e-02 pvsat = -9.771613249e-9
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -9.563480884e-06 lb0 = 1.224511349e-12 wb0 = 6.562808203e-12 pb0 = -8.338986323e-19
+ b1 = 1.366732608e-08 lb1 = -1.749969092e-15 wb1 = -9.379018591e-15 pb1 = 1.191738453e-21
+ keta = -4.810040347e-01 lketa = 4.625438506e-08 wketa = 3.453299969e-07 pketa = -3.518256541e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.140289521e-01 lpclm = 8.769900912e-08 wpclm = 9.028500314e-07 ppclm = -7.608558969e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -2.878028247e-07 lalpha0 = 3.237806959e-14 walpha0 = 2.417309982e-13 palpha0 = -2.462779583e-20
+ alpha1 = 0.85
+ beta0 = 1.922122984e+01 lbeta0 = -4.604857975e-07 wbeta0 = -4.337024874e-06 pbeta0 = 3.847452166e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.412024352e-01 lkt1 = 1.703553167e-08 wkt1 = 1.723344106e-07 pkt1 = -1.466132369e-14
+ kt2 = -0.028878939
+ at = 3.185561747e+05 lat = -2.698172470e-02 wat = -2.014424989e-01 pat = 2.052316323e-8
+ ute = -2.151671721e+00 lute = 1.065141439e-07 wute = 5.704500013e-07 pute = -7.239682022e-14
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.81 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {0.4913699+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56800772
+ k2 = -0.040590746
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 2.78042
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.025731
+ ua = -1.0529435e-9
+ ub = 1.832e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 9.1484e-8
+ b1 = 1.6098e-9
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.82 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.187120042e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.449661691e-06 wvth0 = 3.799652268e-08 pvth0 = -7.581020989e-13
+ k1 = 7.679245717e-01 lk1 = -3.988717236e-06 wk1 = -1.044357338e-07 pk1 = 2.083689333e-12
+ k2 = -1.424839858e-01 lk2 = 2.032961794e-06 wk2 = 5.710978691e-08 pk2 = -1.139447672e-12
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.396630106e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 6.261931899e-07 wvoff = 2.545500732e-08 pvoff = -5.078752768e-13
+ nfactor = 1.984171048e+00 lnfactor = 1.588666433e-05 wnfactor = 6.809304973e-07 pnfactor = -1.358584425e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.015859985e-02 lu0 = 1.111798648e-07 wu0 = 2.574615863e-09 pu0 = -5.136842931e-14
+ ua = -1.855799642e-09 lua = 1.601849020e-14 wua = 4.125285401e-16 pua = -8.230720340e-21
+ ub = 2.759700979e-18 lub = -1.850937953e-23 wub = -5.419275314e-25 pub = 1.081247362e-29
+ uc = 6.616718905e-11 luc = -3.517554340e-16 wuc = -1.949271528e-18 puc = 3.889163357e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.059995482e+00 la0 = 6.037529330e-06 wa0 = 2.218676628e-07 pa0 = -4.426677206e-12
+ ags = 6.098023488e-01 lags = -5.285699177e-06 wags = -1.937215340e-07 pags = 3.865108994e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 6.204682837e-07 lb0 = -1.055423148e-11 wb0 = -3.562509678e-13 pb0 = 7.107876915e-18
+ b1 = 6.469143135e-09 lb1 = -9.695303596e-14 wb1 = -2.884771629e-15 pb1 = 5.755662025e-20
+ keta = -3.543441538e-02 lketa = 6.162700169e-07 wketa = 2.197547238e-08 pketa = -4.384520099e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.589161037e-01 lpclm = 3.507363183e-06 wpclm = 1.001151866e-07 ppclm = -1.997486290e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -8.268913408e-03 lpdiblc2 = 1.841407155e-07 wpdiblc2 = 5.916190072e-09 ppdiblc2 = -1.180391203e-13
+ pdiblcb = 1.225981116e+01 lpdiblcb = -2.451050903e-04 wpdiblcb = -8.238587476e-06 ppdiblcb = 1.643753169e-10
+ drout = 0.56
+ pscbe1 = -5.577131782e+08 lpscbe1 = 1.561660019e+04 wpscbe1 = 3.249333855e+02 ppscbe1 = -6.483032240e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.757211891e-01 lkt1 = -2.126633257e-07 wkt1 = -5.032801248e-09 pkt1 = 1.004138516e-13
+ kt2 = -3.508056030e-02 lkt2 = 1.109849178e-07 wkt2 = -2.453866191e-10 pkt2 = 4.895924623e-15
+ at = 1.981929863e+05 lat = -4.627437017e-1
+ ute = -8.896307601e-01 lute = -4.504521008e-06 wute = -8.488157329e-08 pute = 1.693547049e-12
+ ua1 = 4.953095126e-10 lua1 = 1.248370215e-14 wua1 = 3.586809845e-16 pua1 = -7.156360320e-21
+ ub1 = 1.294816353e-19 lub1 = -1.394539985e-23 wub1 = -3.438454883e-25 pub1 = 6.860364264e-30
+ uc1 = 9.625058006e-11 luc1 = -1.245640185e-15 wuc1 = -1.813948517e-17 puc1 = 3.619168495e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.83 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.909507229e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.003989620e-08 wvth0 = -4.930250957e-08 pvth0 = -6.391058306e-14
+ k1 = 6.033211652e-01 lk1 = -2.679810535e-06 wk1 = -1.113117087e-07 pk1 = 2.138366267e-12
+ k2 = -2.066163692e-03 lk2 = 9.163759830e-07 wk2 = 7.377440934e-09 pk2 = -7.439819753e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.075199276e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 3.705952184e-07 wvoff = -7.027909199e-09 pvoff = -2.495749902e-13
+ nfactor = 7.911571456e+00 lnfactor = -3.124731835e-05 wnfactor = -4.202682967e-06 pnfactor = 2.524806886e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 5.077532826e-02 lu0 = -1.322807162e-07 wu0 = -1.582092918e-08 pu0 = 9.491075579e-14
+ ua = 2.017236972e-09 lua = -1.477943606e-14 wua = -2.008545548e-15 pua = 1.102137270e-20
+ ub = -9.704715590e-19 lub = 1.115250860e-23 wub = 1.884866807e-24 pub = -8.485106170e-30
+ uc = 1.492738782e-10 luc = -1.012609936e-15 wuc = -9.360181824e-17 puc = 7.677017784e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 2.144127744e+00 la0 = -2.583361407e-06 wa0 = -4.930556356e-07 pa0 = 1.258307787e-12
+ ags = 1.761942869e-01 lags = -1.837699468e-06 wags = 1.239986717e-07 pags = 1.338635727e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -3.733988909e-07 lb0 = -2.651117977e-12 wb0 = 2.840191452e-13 pb0 = 2.016525169e-18
+ b1 = 1.235600041e-08 lb1 = -1.437646245e-13 wb1 = -9.398369306e-15 pb1 = 1.093519739e-19
+ keta = 2.241656438e-02 lketa = 1.562459101e-07 wketa = -2.670388401e-08 pketa = -5.135956067e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.092982737e+00 lpclm = -1.439946843e-05 wpclm = -1.866341298e-06 ppclm = 1.363954167e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 3.710228660e-02 lpdiblc2 = -1.766456678e-07 wpdiblc2 = -2.597090179e-08 ppdiblc2 = 1.355232396e-13
+ pdiblcb = -3.687943347e+01 lpdiblcb = 1.456443354e-04 wpdiblcb = 2.471576243e-05 ppdiblcb = -9.767375194e-11
+ drout = 0.56
+ pscbe1 = 1.808679028e+09 lpscbe1 = -3.200669031e+03 wpscbe1 = -7.842692750e+02 ppscbe1 = 2.337215321e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.282676684e-01 lkt1 = 2.051800245e-07 wkt1 = 2.814556841e-08 pkt1 = -1.634165957e-13
+ kt2 = -1.004165202e-01 lkt2 = 6.305286958e-07 wkt2 = 6.072950364e-08 pkt2 = -4.799691467e-13
+ at = 140000.0
+ ute = -3.396942908e+00 lute = 1.543332682e-05 wute = 1.452408034e-06 pute = -1.053079697e-11
+ ua1 = -6.949192448e-10 lua1 = 2.194825959e-14 wua1 = 1.481593296e-15 pua1 = -1.608562540e-20
+ ub1 = -2.619106371e-19 lub1 = -1.083309508e-23 wub1 = -5.126766683e-25 pub1 = 8.202889717e-30
+ uc1 = 2.708030707e-10 luc1 = -2.633660819e-15 wuc1 = -2.291489405e-16 puc1 = 2.039838929e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.84 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {3.704232332e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.515382927e-07 wvth0 = 1.042304588e-07 pvth0 = -6.706546036e-13
+ k1 = -4.293198183e-01 lk1 = 1.401063748e-06 wk1 = 6.629569781e-07 pk1 = -9.214514450e-13
+ k2 = 3.729117309e-01 lk2 = -5.654920341e-07 wk2 = -2.725128435e-07 pk2 = 3.621111219e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -1.621656431e+00 ldsub = 8.621646599e-06 wdsub = 1.659437695e-06 pdsub = -6.557900296e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {2.885946907e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.194802615e-06 wvoff = -2.854227260e-07 pvoff = 8.506081969e-13
+ nfactor = 3.725942809e+00 lnfactor = -1.470621203e-05 wnfactor = -3.539381328e-07 pnfactor = 1.003828728e-11
+ eta0 = -4.981389543e-01 leta0 = 2.284736349e-06 weta0 = 4.397509891e-07 peta0 = -1.737843579e-12
+ etab = 4.354170733e-01 letab = -1.997348129e-06 wetab = -3.844363993e-07 petab = 1.519246902e-12
+ u0 = 2.416659232e-02 lu0 = -2.712615822e-08 wu0 = 3.654622243e-09 pu0 = 1.794569416e-14
+ ua = 3.135504344e-09 lua = -1.919869564e-14 wua = -2.572908972e-15 pua = 1.325166979e-20
+ ub = -5.111143675e-18 lub = 2.751595206e-23 wub = 4.604017907e-24 pub = -1.923086774e-29
+ uc = -2.881685016e-10 luc = 7.161102928e-16 wuc = 2.171752061e-16 puc = -4.604520395e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = -3.658847585e-01 la0 = 7.335909313e-06 wa0 = 1.322363605e-06 pa0 = -5.916013015e-12
+ ags = -7.005904371e-01 lags = 1.627249424e-06 wags = 6.896052766e-07 pags = -8.965742688e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.939546512e-07 lb0 = -1.779507858e-12 wb0 = 4.517809143e-13 pb0 = 1.353550621e-18
+ b1 = -5.986302450e-09 lb1 = -7.127802632e-14 wb1 = 4.553373205e-15 pb1 = 5.421634772e-20
+ keta = 2.318643214e-01 lketa = -6.714667013e-07 wketa = -1.551298792e-07 pketa = 4.561646897e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.981965627e+00 lpclm = 9.608004593e-06 wpclm = 3.416585042e-06 ppclm = -7.237954557e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -6.485716908e-03 lpdiblc2 = -4.391064887e-09 wpdiblc2 = 6.028050252e-09 ppdiblc2 = 9.067189034e-15
+ pdiblcb = 6.590235130e-02 lpdiblcb = -3.592352750e-07 wpdiblcb = -6.914323728e-08 ppdiblcb = 2.732458457e-13
+ drout = 0.56
+ pscbe1 = 1.192755226e+09 lpscbe1 = -7.666114643e+02 wpscbe1 = -3.810617629e+02 ppscbe1 = 7.437872147e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.678350503e-01 lkt1 = 1.151921809e-06 wkt1 = 2.070013522e-07 pkt1 = -8.702333693e-13
+ kt2 = -8.816029381e-02 lkt2 = 5.820935477e-07 wkt2 = 4.908699713e-08 pkt2 = -4.339593464e-13
+ at = 1.547989822e+05 lat = -5.848381645e-02 wat = 1.012256994e-02 pat = -4.000319181e-8
+ ute = -8.094701062e+00 lute = 3.399830801e-05 wute = 4.839234518e-06 pute = -2.391513220e-11
+ ua1 = -2.131947734e-08 lua1 = 1.034540589e-13 wua1 = 1.572350355e-14 pua1 = -7.236795995e-20
+ ub1 = 1.773205346e-17 lub1 = -8.194309992e-23 wub1 = -1.288161491e-23 pub1 = 5.708346173e-29
+ uc1 = -1.210052667e-10 luc1 = -1.085280895e-15 wuc1 = 8.699191685e-17 puc1 = 7.904878808e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.85 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {8.126625796e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.833971508e-08 wvth0 = -2.241407457e-07 pvth0 = -2.971308852e-14
+ k1 = 6.382875525e-01 lk1 = -6.827787948e-07 wk1 = -3.164620115e-08 pk1 = 4.343313031e-13
+ k2 = 1.377507430e-02 lk2 = 1.354999824e-07 wk2 = -4.818232781e-08 pk2 = -7.575534940e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 5.208877163e+00 ldsub = -4.710742142e-06 wdsub = -3.318875389e-06 pdsub = 3.159174424e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-3.691774056e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 8.909024160e-08 wvoff = 2.035408227e-07 pvoff = -1.037904635e-13
+ nfactor = 2.902132580e-01 lnfactor = -8.000076798e-06 wnfactor = 1.974170091e-06 pnfactor = 5.494097074e-12
+ eta0 = 1.310018538e+00 leta0 = -1.244571905e-06 weta0 = -8.795017084e-07 peta0 = 8.371806960e-13
+ etab = -1.067150857e+00 letab = 9.354856657e-07 wetab = 7.688727985e-07 petab = -7.318754083e-13
+ u0 = 7.228735220e-03 lu0 = 5.934523236e-09 wu0 = 1.635532283e-08 pu0 = -6.844562002e-15
+ ua = -9.966303185e-09 lua = 6.374473543e-15 wua = 6.868290396e-15 pua = -5.176427870e-21
+ ub = 1.416526203e-17 lub = -1.010929799e-23 wub = -9.273255750e-24 pub = 7.855919041e-30
+ uc = -1.301082669e-10 luc = 4.075955238e-16 wuc = 1.284894387e-16 puc = -2.873479751e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.378147357e+04 lvsat = 1.097318736e-01 wvsat = 3.552129870e-02 pvsat = -6.933334804e-8
+ a0 = 8.550989633e+00 la0 = -1.006876839e-05 wa0 = -5.394763498e-06 pa0 = 7.195019752e-12
+ ags = 4.815035729e+00 lags = -9.138596492e-06 wags = -3.403399240e-06 pags = 7.092483481e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -8.338029628e-07 lb0 = -1.311352496e-12 wb0 = 6.342172152e-13 pb0 = 9.974566716e-19
+ b1 = -3.149500611e-08 lb1 = -2.148807231e-14 wb1 = 2.395610949e-14 pb1 = 1.634451541e-20
+ keta = -7.402086627e-01 lketa = 1.225904087e-06 wketa = 5.429904074e-07 pketa = -9.064830335e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.471614655e+00 lpclm = -2.988616142e-06 wpclm = -1.551256085e-06 ppclm = 2.458680149e-12
+ pdiblc1 = 5.499285885e-01 lpdiblc1 = -3.121615733e-07 wpdiblc1 = -8.450734923e-08 ppdiblc1 = 1.649482893e-13
+ pdiblc2 = -3.046528683e-02 lpdiblc2 = 4.241420204e-08 wpdiblc2 = 2.683279202e-08 ppdiblc2 = -3.154119114e-14
+ pdiblcb = 1.652317102e-01 lpdiblcb = -5.531143634e-07 wpdiblcb = -1.270498481e-07 ppdiblcb = 3.862726590e-13
+ drout = 4.420233479e+00 ldrout = -7.534716383e-06 wdrout = -2.818417106e-06 pdrout = 5.501214800e-12
+ pscbe1 = 3.311384645e+08 lpscbe1 = 9.151619228e+02 wpscbe1 = 3.566310875e+02 ppscbe1 = -6.961014437e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.897972713e-05 lalpha0 = -7.602523235e-11 walpha0 = -2.962554001e-11 palpha0 = 5.782552867e-17
+ alpha1 = 2.080852953e+00 lalpha1 = -2.402478493e-06 walpha1 = -8.254493775e-07 palpha1 = 1.611178956e-12
+ beta0 = 3.942284599e+01 lbeta0 = -4.989563339e-05 wbeta0 = -1.944391867e-05 pbeta0 = 3.795221542e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 1.600730101e-01 lkt1 = -2.688681037e-07 wkt1 = -3.689878470e-07 pkt1 = 2.540290049e-13
+ kt2 = 5.090511116e-01 lkt2 = -5.835920475e-07 wkt2 = -3.872479470e-07 pkt2 = 4.177145406e-13
+ at = -1.253319492e+03 lat = 2.461117062e-01 wat = 1.039875271e-01 pat = -2.232164183e-7
+ ute = 1.899759215e+01 lute = -1.888262436e-05 wute = -1.431948635e-05 pute = 1.348041104e-11
+ ua1 = 6.090476834e-08 lua1 = -5.703788403e-14 wua1 = -4.186780254e-14 pua1 = 4.004341619e-20
+ ub1 = -4.591090728e-17 lub1 = 4.228038594e-23 wub1 = 3.141482312e-23 pub1 = -2.937791401e-29
+ uc1 = -1.175732069e-09 luc1 = 9.734203110e-16 wuc1 = 8.363672937e-16 puc1 = -6.722036792e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.86 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {1.246742175e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.248524047e-07 wvth0 = -4.861368115e-07 pvth0 = 2.196759885e-13
+ k1 = -5.796825371e-01 lk1 = 4.765837920e-07 wk1 = 8.084157711e-07 pk1 = -3.653077270e-13
+ k2 = 3.094428308e-01 lk2 = -1.459405374e-07 wk2 = -2.432383836e-07 pk2 = 1.099148040e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.145343276e-01 ldsub = 4.327790972e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-3.948322855e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.135106343e-07 wvoff = 1.799123567e-07 pvoff = -8.129897565e-14
+ nfactor = -1.817246299e+01 lnfactor = 9.574193934e-06 wnfactor = 1.474654415e-05 pnfactor = -6.663683117e-12
+ eta0 = -4.380236780e-01 leta0 = 4.193562676e-07 weta0 = -5.395093970e-13 peta0 = 2.437940460e-19
+ etab = -1.600650675e-01 letab = 7.204793715e-8
+ u0 = 3.545515521e-03 lu0 = 9.440510085e-09 wu0 = 1.744751810e-08 pu0 = -7.884201926e-15
+ ua = -4.915110148e-09 lua = 1.566338864e-15 wua = 2.722734521e-15 pua = -1.230351998e-21
+ ub = 4.807537174e-18 lub = -1.201857491e-24 wub = -1.942233830e-24 pub = 8.776585651e-31
+ uc = 5.200149291e-10 luc = -2.112443941e-16 wuc = -3.300826393e-16 puc = 1.491580731e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.409208113e+05 lvsat = -1.770836388e-03 wvsat = -7.104259741e-02 pvsat = 3.210279996e-8
+ a0 = -5.109836523e+00 la0 = 2.934712471e-06 wa0 = 4.119693756e-06 pa0 = -1.861611334e-12
+ ags = -9.251723749e+00 lags = 4.251284586e-06 wags = 7.705704817e-06 pags = -3.482061598e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -4.210067388e-06 lb0 = 1.902449461e-12 wb0 = 3.202311977e-12 pb0 = -1.447063939e-18
+ b1 = -1.029351404e-07 lb1 = 4.651443419e-14 wb1 = 7.829576174e-14 pb1 = -3.538036711e-20
+ keta = 1.049055792e+00 lketa = -4.772627513e-07 wketa = -7.792415630e-07 pketa = 3.521244567e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.680194935e+00 lpclm = 9.634125218e-07 wpclm = 1.964137911e-06 ppclm = -8.875566034e-13
+ pdiblc1 = 3.927571236e-01 lpdiblc1 = -1.625530421e-07 wpdiblc1 = 1.690146985e-07 ppdiblc1 = -7.637453096e-14
+ pdiblc2 = 2.678778009e-02 lpdiblc2 = -1.208390456e-08 wpdiblc2 = -1.199913247e-08 ppdiblc2 = 5.422179979e-15
+ pdiblcb = -7.061662818e-01 lpdiblcb = 2.763528287e-07 wpdiblcb = 5.306726452e-07 ppdiblcb = -2.398008856e-13
+ drout = -7.558122148e+00 ldrout = 3.867252749e-06 wdrout = 5.636834212e-06 pdrout = -2.547178281e-12
+ pscbe1 = 2.065836567e+09 lpscbe1 = -7.360642418e+02 wpscbe1 = -7.132621750e+02 ppscbe1 = 3.223096249e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -8.136701321e-05 lalpha0 = 3.853054320e-11 walpha0 = 5.925108003e-11 palpha0 = -2.677443729e-17
+ alpha1 = -1.611705906e+00 lalpha1 = 1.112398126e-06 walpha1 = 1.650898755e-06 palpha1 = -7.460097803e-13
+ beta0 = -4.102353437e+01 lbeta0 = 2.667974759e-05 wbeta0 = 3.888783734e-05 pbeta0 = -1.757267483e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 1.910873679e-02 lkt1 = -1.346868903e-07 wkt1 = -1.944070319e-07 pkt1 = 8.784884400e-14
+ kt2 = -1.648870573e-01 lkt2 = 5.791689064e-08 wkt2 = 9.820115517e-08 pkt2 = -4.437523620e-14
+ at = 4.802075712e+05 lat = -2.121817679e-01 wat = -2.484653340e-01 pat = 1.122767636e-7
+ ute = -4.141744093e-01 lute = -4.049325934e-07 wute = -3.000718896e-07 pute = 1.355967855e-13
+ ua1 = 1.120784177e-09 lua1 = -1.306453975e-16 wua1 = 3.805008715e-16 pua1 = -1.719411143e-22
+ ub1 = -2.271600555e-18 lub1 = 7.409590158e-25 wub1 = 1.050518455e-24 pub1 = -4.747093299e-31
+ uc1 = -2.966613942e-10 luc1 = 1.366496379e-16 wuc1 = 2.478369135e-16 puc1 = -1.119927923e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.87 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.750340240e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.132025349e-8
+ k1 = 1.260614571e-01 lk1 = 1.576714902e-7
+ k2 = 8.475738853e-02 lk2 = -4.440945505e-08 wk2 = -2.775557562e-23 pk2 = -2.081668171e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.905328527e-01 ldsub = 5.412372020e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.103590353e-03 lcdscd = -1.221701112e-9
+ cit = 0.0
+ voff = {-1.154994111e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.271458427e-8
+ nfactor = 3.206634077e+00 lnfactor = -8.661382834e-8
+ eta0 = 8.851262253e-01 leta0 = -1.785500338e-7
+ etab = 3.439973846e-02 letab = -1.582701384e-08 wetab = 5.204170428e-24 petab = -1.301042607e-30
+ u0 = 2.025864782e-02 lu0 = 1.888163151e-9
+ ua = -1.664072323e-09 lua = 9.725664082e-17
+ ub = 2.065347559e-18 lub = 3.728589477e-26
+ uc = 2.021746693e-11 luc = 1.460458292e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.342184647e+05 lvsat = 1.257826697e-3
+ a0 = 1.291411731e+00 la0 = 4.211000822e-8
+ ags = -7.269793732e-01 lags = 3.991145728e-07 wags = -2.220446049e-22 pags = -2.220446049e-28
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.316735352e-16 lb0 = -2.658238496e-23
+ b1 = -6.482321705e-18 lb1 = 1.308657588e-24
+ keta = 5.428652146e-02 lketa = -2.774541862e-08 wketa = -2.775557562e-23 pketa = 8.673617380e-30
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.240064173e-01 lpclm = -7.781228934e-8
+ pdiblc1 = -2.285578198e-01 lpdiblc1 = 1.182073759e-07 wpdiblc1 = -5.551115123e-23 ppdiblc1 = 1.387778781e-29
+ pdiblc2 = -6.704200072e-03 lpdiblc2 = 3.050484931e-09 wpdiblc2 = -2.168404345e-25 ppdiblc2 = -4.878909776e-31
+ pdiblcb = -8.758737421e-02 lpdiblcb = -3.171226653e-9
+ drout = 1.401075462e+00 ldrout = -1.812384259e-7
+ pscbe1 = 1.507016608e+08 lpscbe1 = 1.293488348e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.031901082e-06 lalpha0 = -1.415246593e-12
+ alpha1 = 0.85
+ beta0 = 2.100422375e+01 lbeta0 = -1.349417775e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.096264800e-01 lkt1 = 1.386230826e-8
+ kt2 = -4.304931441e-02 lkt2 = 2.860729557e-9
+ at = -3.932844299e+03 lat = 6.592087176e-03 pat = -3.637978807e-24
+ ute = -1.303201518e+00 lute = -3.198134688e-9
+ ua1 = 1.522520005e-09 lua1 = -3.121821852e-16
+ ub1 = -1.713664128e-18 lub1 = 4.888381454e-25 pub1 = 1.925929944e-46
+ uc1 = -1.084804678e-10 luc1 = 5.161425266e-17 wuc1 = -1.292469707e-32 puc1 = -1.292469707e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.88 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {6.130803429e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.900108240e-8
+ k1 = 9.070734896e-01 lk1 = 5.142863913e-17
+ k2 = -1.611477193e-01 lk2 = 5.234114019e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -7.794653811e-18
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999996e-03 lcdscd = 5.442087753e-19
+ cit = 0.0
+ voff = {-1.237493848e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.104907131e-8
+ nfactor = 2.484263783e+00 lnfactor = 5.921900879e-8
+ eta0 = 2.001909455e-03 leta0 = -2.640137943e-10
+ etab = -4.399800002e-02 letab = 2.220584827e-18
+ u0 = 2.919169366e-02 lu0 = 8.475092343e-11
+ ua = -1.224106221e-09 lua = 8.435844238e-18
+ ub = 2.103521860e-18 lub = 2.957922859e-26
+ uc = 1.218677263e-10 luc = -5.916673095e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.325369855e+05 lvsat = 1.597285411e-3
+ a0 = 1.499999999e+00 la0 = 1.571054398e-16
+ ags = 1.250000000e+00 lags = 3.363798129e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -6.898412508e-08 lb0 = 1.392658415e-14
+ b1 = 9.858632274e-11 lb1 = -1.990270542e-17
+ keta = -1.889316341e-01 lketa = 2.135570583e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.499568007e-01 lpclm = -2.248687870e-8
+ pdiblc1 = 3.569721502e-01 lpdiblc1 = -2.689604095e-17
+ pdiblc2 = 8.406112095e-03 lpdiblc2 = 7.211488351e-19
+ pdiblcb = -1.032957700e-01 lpdiblcb = 2.135236432e-18
+ drout = 5.033266589e-01 ldrout = 1.424533824e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 1.407241821e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 5.774280622e-09 lalpha0 = 3.194912098e-15
+ alpha1 = 0.85
+ beta0 = 1.518074234e+01 lbeta0 = -1.737675240e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.585636645e-01 lkt1 = 3.553695993e-9
+ kt2 = -2.887893901e-02 lkt2 = 8.536227281e-19
+ at = -1.837987011e+04 lat = 9.508667194e-3
+ ute = -1.325229293e+00 lute = 1.248854588e-9
+ ua1 = -2.384733722e-11 lua1 = 1.610623404e-25
+ ub1 = 7.077531683e-19 lub1 = 2.287970107e-34
+ uc1 = 1.471862500e-10 luc1 = -3.312754956e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.89 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {-7.830981281e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.551283305e-07 wvth0 = 9.819012935e-07 pvth0 = -1.294941245e-13
+ k1 = 0.90707349
+ k2 = -4.031459864e-01 lk2 = 3.714908748e-08 wk2 = 1.403207628e-07 pk2 = -1.850564252e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.45863
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999998e-03 lcdscd = 2.552394060e-19 wcdscd = 1.963887386e-18 pcdscd = -2.589994191e-25
+ cit = 0.0
+ voff = {-2.075300001e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.193267707e-17
+ nfactor = 8.275709919e+00 lnfactor = -7.045626990e-07 wnfactor = -3.582792759e-06 pnfactor = 4.725022919e-13
+ eta0 = 8.801219272e-10 leta0 = -8.964436628e-17 weta0 = 5.138788330e-19 peta0 = -6.777085437e-26
+ etab = -0.043998
+ u0 = 1.793886886e-01 lu0 = -1.972337897e-08 wu0 = -1.006927941e-07 pu0 = 1.327946637e-14
+ ua = -1.238295631e-09 lua = 1.030715774e-17 wua = 5.241323476e-17 pua = -6.912309813e-24
+ ub = 4.818240523e-18 lub = -3.284405833e-25 wub = -1.670162989e-24 pub = 2.202627652e-31
+ uc = 7.700399988e-11 luc = 1.171365296e-26 wuc = -1.348304398e-28 puc = 1.778438317e-35
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.159709097e+04 lvsat = 1.359052964e-02 wvsat = 8.599900705e-02 pvsat = -1.134163505e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -8.178187945e-06 lb0 = 1.083376493e-12 wb0 = 5.509110064e-12 pb0 = -7.265469443e-19
+ b1 = 1.168755196e-08 lb1 = -1.548267082e-15 wb1 = -7.873139042e-15 pb1 = 1.038317450e-21
+ keta = -2.700000006e-02 lketa = 6.295935995e-18 wketa = 7.693845561e-20 pketa = -1.014466289e-26
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 9.696314362e-01 lpclm = -1.042101893e-07 wpclm = -5.299223370e-07 ppclm = 6.988668773e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.000000001e-08 lalpha0 = -1.407093779e-24 walpha0 = -1.540541173e-25 palpha0 = 2.031555584e-32
+ alpha1 = 0.85
+ beta0 = 1.095773815e+01 lbeta0 = 3.831664914e-07 wbeta0 = 1.948451340e-06 pbeta0 = -2.569637112e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -8.809131195e-02 lkt1 = -1.892836833e-08 wkt1 = -9.625320927e-08 pkt1 = 1.269396949e-14
+ kt2 = -0.028878939
+ at = 5.372048693e+04 lat = 6.909540389e-12 wat = -3.282912076e-14 pat = 4.307366908e-21
+ ute = -2.042108666e+00 lute = 9.579162324e-08 wute = 4.871128358e-07 pute = -6.424092790e-14
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.90 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {0.4913699+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56800772
+ k2 = -0.040590746
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 2.78042
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.025731
+ ua = -1.0529435e-9
+ ub = 1.832e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 9.1484e-8
+ b1 = 1.6098e-9
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.91 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.753697877e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.192323364e-7
+ k1 = 6.121972372e-01 lk1 = -8.816639883e-7
+ k2 = -5.732582613e-02 lk2 = 3.338963274e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.017062664e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.311152548e-7
+ nfactor = 2.999527454e+00 lnfactor = -4.371605856e-06 wnfactor = -2.842170943e-20
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.399768874e-02 lu0 = 3.458282001e-08 wu0 = -2.220446049e-22
+ ua = -1.240665649e-09 lua = 3.745409973e-15
+ ub = 1.951616170e-18 lub = -2.386567588e-24
+ uc = 6.326057033e-11 luc = -2.937629231e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.390829178e+00 la0 = -5.632251912e-7
+ ags = 3.209382116e-01 lags = 4.776837126e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 8.925150941e-08 lb0 = 4.454238660e-14
+ b1 = 2.167571440e-09 lb1 = -1.112858939e-14
+ keta = -2.666112675e-03 lketa = -3.751925933e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.631270000e-03 lpclm = 5.288499448e-07 ppclm = 1.776356839e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 5.528995573e-04 lpdiblc2 = 8.128953030e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -7.319501400e+07 lpscbe1 = 5.949551434e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.832257539e-01 lkt1 = -6.293314343e-8
+ kt2 = -3.544646383e-02 lkt2 = 1.182853816e-7
+ at = 1.981929862e+05 lat = -4.627437017e-1
+ ute = -1.016200285e+00 lute = -1.979220918e-6
+ ua1 = 1.030149760e-09 lua1 = 1.812633186e-15
+ ub1 = -3.832369470e-19 lub1 = -3.715699712e-24
+ uc1 = 6.920223587e-11 luc1 = -7.059748407e-16 puc1 = -3.308722450e-36
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.92 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.174342346e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.525913972e-8
+ k1 = 4.373408531e-01 lk1 = 5.087731700e-7
+ k2 = 8.934565372e-03 lk2 = -1.929984209e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.179994591e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.553724997e-9
+ nfactor = 1.644821634e+00 lnfactor = 6.400853618e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.718425420e-02 lu0 = 9.243630640e-9
+ ua = -9.777670666e-10 lua = 1.654871732e-15
+ ub = 1.840111304e-18 lub = -1.499894165e-24
+ uc = 9.701328365e-12 luc = 1.321337955e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.408917323e+00 la0 = -7.070599674e-7
+ ags = 3.610925198e-01 lags = 1.583814327e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 5.011079129e-08 lb0 = 3.557847194e-13
+ b1 = -1.658197099e-09 lb1 = 1.929346677e-14
+ keta = -1.740241834e-02 lketa = 7.966208966e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -6.899761706e-01 lpclm = 5.938871634e-06 ppclm = 3.552713679e-27
+ pdiblc1 = 0.39
+ pdiblc2 = -1.623723774e-03 lpdiblc2 = 2.543720274e-08 ppdiblc2 = 1.110223025e-28
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.392309919e+08 lpscbe1 = 2.844246136e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.862989458e-01 lkt1 = -3.849548711e-8
+ kt2 = -9.860889619e-03 lkt2 = -8.516805990e-8
+ at = 140000.0
+ ute = -1.231212620e+00 lute = -2.694684098e-7
+ ua1 = 1.514330084e-09 lua1 = -2.037511139e-15 wua1 = -1.323488980e-29
+ ub1 = -1.026378584e-18 lub1 = 1.398486053e-24
+ uc1 = -7.088796187e-11 luc1 = 4.080057410e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.93 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.258444758e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.849541224e-8
+ k1 = 5.592357205e-01 lk1 = 2.705915957e-8
+ k2 = -3.344055097e-02 lk2 = -2.553700375e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.527821500e-01 ldsub = -1.157040216e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.370079140e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 7.356542684e-8
+ nfactor = 3.198174774e+00 lnfactor = 2.621868556e-7
+ eta0 = 1.575872698e-01 leta0 = -3.066156572e-7
+ etab = -1.378278648e-01 letab = 2.680476500e-7
+ u0 = 2.961611194e-02 lu0 = -3.667817484e-10
+ ua = -7.010393526e-10 lua = 5.612767375e-16
+ ub = 1.754049020e-18 lub = -1.159786258e-24
+ uc = 3.566812735e-11 luc = 2.951609590e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.605932281e+00 la0 = -1.485639637e-6
+ ags = 3.277011992e-01 lags = 2.903399581e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 7.970976424e-08 lb0 = 2.388131005e-13
+ b1 = 8.033723719e-10 lb1 = 9.565637143e-15
+ keta = 5.453875497e-04 lketa = 8.734496589e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.112609403e+00 lpclm = -1.184732045e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.502894210e-03 lpdiblc2 = 9.129299537e-9
+ pdiblcb = -3.719925625e-02 lpdiblcb = 4.821000899e-8
+ drout = 0.56
+ pscbe1 = 6.245423126e+08 lpscbe1 = 3.424725263e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.591689679e-01 lkt1 = -1.457099312e-7
+ kt2 = -1.496516276e-02 lkt2 = -6.499657985e-8
+ at = 1.698930575e+05 lat = -1.181338060e-1
+ ute = -8.787696445e-01 lute = -1.662281110e-6
+ ua1 = 2.126322375e-09 lua1 = -4.456031847e-15
+ ub1 = -1.476118686e-18 lub1 = 3.175805416e-24
+ uc1 = 8.711055893e-12 luc1 = 9.343989506e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.94 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.784394203e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.403361498e-8
+ k1 = 5.910989287e-01 lk1 = -3.513403122e-8
+ k2 = -5.807107652e-02 lk2 = 2.253885108e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.26
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-6.567142512e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -6.567491050e-8
+ nfactor = 3.233958994e+00 lnfactor = 1.923403166e-7
+ eta0 = -1.433508281e-03 leta0 = 3.773978078e-09 weta0 = 6.938893904e-24
+ etab = 7.933901888e-02 letab = -1.558362640e-07 wetab = 1.179611964e-22 petab = 3.053113318e-28
+ u0 = 3.161666009e-02 lu0 = -4.271613666e-9
+ ua = 2.752158536e-10 lua = -1.344257251e-15
+ ub = 3.376251922e-19 lub = 1.604904499e-24
+ uc = 6.148628680e-11 luc = -2.087787897e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.674837450e+04 lvsat = 6.346786025e-3
+ a0 = 5.066918688e-01 la0 = 6.599468372e-7
+ ags = -2.598775476e-01 lags = 1.437223750e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.118978317e-07 lb0 = 1.759858233e-13
+ b1 = 4.226685500e-09 lb1 = 2.883737292e-15
+ keta = 6.946103312e-02 lketa = -1.257806426e-07 wketa = -1.665334537e-22 pketa = 4.440892099e-28
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.584889993e-01 lpclm = 6.775974424e-7
+ pdiblc1 = 4.239170811e-01 lpdiblc1 = -6.620210620e-8
+ pdiblc2 = 9.545914571e-03 lpdiblc2 = -4.617838089e-9
+ pdiblcb = -2.421622557e-02 lpdiblcb = 2.286867807e-8
+ drout = 2.176050537e-01 ldrout = 6.683141902e-7
+ pscbe1 = 8.629220470e+08 lpscbe1 = -1.228163479e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.195826690e-06 lalpha0 = 1.020019183e-11 walpha0 = 1.101142831e-26 palpha0 = 1.694065895e-32
+ alpha1 = 0.85
+ beta0 = 1.042942088e+01 lbeta0 = 6.696082211e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.901361166e-01 lkt1 = 1.099223579e-7
+ kt2 = -6.838621167e-02 lkt2 = 3.927495052e-8
+ at = 1.538056803e+05 lat = -8.673316007e-2
+ ute = -2.354634327e+00 lute = 1.218431122e-6
+ ua1 = -1.525599643e-09 lua1 = 2.672085355e-15 wua1 = -1.654361225e-30 pua1 = -6.617444900e-36
+ ub1 = 9.327016030e-19 lub1 = -1.525925138e-24 wub1 = -3.081487911e-39 pub1 = 1.540743956e-45
+ uc1 = 7.140092441e-11 luc1 = -2.892326820e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.95 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.218486251e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.713217742e-9
+ k1 = 6.257710814e-01 lk1 = -6.813779454e-8
+ k2 = -5.325740349e-02 lk2 = 1.795680719e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.145343276e-01 ldsub = 4.327790972e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.265594373e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.716768537e-9
+ nfactor = 3.816562507e+00 lnfactor = -3.622288973e-7
+ eta0 = -4.380244825e-01 leta0 = 4.193566312e-07 weta0 = 7.771561172e-22 peta0 = 1.332267630e-27
+ etab = -1.600650675e-01 letab = 7.204793715e-8
+ u0 = 2.956204634e-02 lu0 = -2.315865879e-9
+ ua = -8.551569683e-10 lua = -2.682768386e-16
+ ub = 1.911412579e-18 lub = 1.068461874e-25
+ uc = 2.781855420e-11 luc = 1.116979601e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.498700947e+04 lvsat = 4.609863593e-2
+ a0 = 1.033165535e+00 la0 = 1.588065578e-7
+ ags = 2.238489687e+00 lags = -9.409245514e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 5.649984863e-07 lb0 = -2.553120810e-13
+ b1 = 1.381407783e-08 lb1 = -6.242319304e-15
+ keta = -1.128952678e-01 lketa = 4.780085550e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.248591510e+00 lpclm = -3.600504257e-7
+ pdiblc1 = 6.447801384e-01 lpdiblc1 = -2.764374541e-07 wpdiblc1 = 3.552713679e-21
+ pdiblc2 = 8.895504641e-03 lpdiblc2 = -3.998725234e-9
+ pdiblcb = 8.513601992e-02 lpdiblcb = -8.122164671e-08 wpdiblcb = 1.353084311e-22 ppdiblcb = -1.908195824e-29
+ drout = 8.471347030e-01 ldrout = 6.907687805e-8
+ pscbe1 = 1.002269402e+09 lpscbe1 = -2.554584477e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 6.984094440e-06 lalpha0 = -1.393643679e-12
+ alpha1 = 0.85
+ beta0 = 1.696331585e+01 lbeta0 = 4.765917258e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.707775674e-01 lkt1 = -3.692777228e-9
+ kt2 = -1.845629469e-02 lkt2 = -8.252388786e-9
+ at = 1.097132702e+05 lat = -4.476243271e-2
+ ute = -8.616208324e-01 lute = -2.027400563e-7
+ ua1 = 1.688160728e-09 lua1 = -3.870320810e-16
+ ub1 = -7.051401785e-19 lub1 = 3.310533463e-26
+ uc1 = 7.289584949e-11 luc1 = -3.034625898e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.96 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.750340240e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.132025349e-8
+ k1 = 1.260614571e-01 lk1 = 1.576714902e-7
+ k2 = 8.475738853e-02 lk2 = -4.440945505e-08 wk2 = -2.220446049e-22 pk2 = 2.775557562e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.905328527e-01 ldsub = 5.412372020e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.103590353e-03 lcdscd = -1.221701112e-9
+ cit = 0.0
+ voff = {-1.154994111e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.271458427e-8
+ nfactor = 3.206634077e+00 lnfactor = -8.661382834e-8
+ eta0 = 8.851262253e-01 leta0 = -1.785500338e-7
+ etab = 3.439973846e-02 letab = -1.582701384e-08 wetab = 9.714451465e-23 petab = 5.204170428e-30
+ u0 = 2.025864782e-02 lu0 = 1.888163151e-9
+ ua = -1.664072323e-09 lua = 9.725664082e-17
+ ub = 2.065347559e-18 lub = 3.728589477e-26
+ uc = 2.021746693e-11 luc = 1.460458292e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.342184647e+05 lvsat = 1.257826697e-3
+ a0 = 1.291411731e+00 la0 = 4.211000822e-8
+ ags = -7.269793732e-01 lags = 3.991145728e-07 wags = 1.776356839e-21 pags = 8.881784197e-28
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.316735352e-16 lb0 = -2.658238496e-23
+ b1 = -6.482321705e-18 lb1 = 1.308657588e-24
+ keta = 5.428652146e-02 lketa = -2.774541862e-08 wketa = -1.110223025e-22 pketa = 9.714451465e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.240064173e-01 lpclm = -7.781228934e-8
+ pdiblc1 = -2.285578198e-01 lpdiblc1 = 1.182073759e-07 wpdiblc1 = -4.440892099e-22 ppdiblc1 = 1.110223025e-28
+ pdiblc2 = -6.704200072e-03 lpdiblc2 = 3.050484931e-09 wpdiblc2 = 1.734723476e-23 ppdiblc2 = 5.204170428e-30
+ pdiblcb = -8.758737421e-02 lpdiblcb = -3.171226653e-9
+ drout = 1.401075462e+00 ldrout = -1.812384259e-7
+ pscbe1 = 1.507016608e+08 lpscbe1 = 1.293488348e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.031901082e-06 lalpha0 = -1.415246593e-12
+ alpha1 = 0.85
+ beta0 = 2.100422375e+01 lbeta0 = -1.349417775e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.096264800e-01 lkt1 = 1.386230826e-8
+ kt2 = -4.304931441e-02 lkt2 = 2.860729557e-9
+ at = -3.932844299e+03 lat = 6.592087176e-03 pat = -2.910383046e-23
+ ute = -1.303201518e+00 lute = -3.198134688e-9
+ ua1 = 1.522520005e-09 lua1 = -3.121821852e-16
+ ub1 = -1.713664128e-18 lub1 = 4.888381454e-25 wub1 = 6.162975822e-39 pub1 = -1.540743956e-45
+ uc1 = -1.084804678e-10 luc1 = 5.161425266e-17 wuc1 = -2.584939414e-31 puc1 = -1.292469707e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.97 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {6.130803429e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.900108240e-8
+ k1 = 9.070734896e-01 lk1 = 5.142908321e-17
+ k2 = -1.611477193e-01 lk2 = 5.234114019e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -7.792877454e-18
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999996e-03 lcdscd = 5.442105100e-19
+ cit = 0.0
+ voff = {-1.237493848e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.104907131e-8
+ nfactor = 2.484263783e+00 lnfactor = 5.921900879e-8
+ eta0 = 2.001909455e-03 leta0 = -2.640137943e-10
+ etab = -4.399800002e-02 letab = 2.220668094e-18
+ u0 = 2.919169366e-02 lu0 = 8.475092343e-11
+ ua = -1.224106221e-09 lua = 8.435844238e-18
+ ub = 2.103521860e-18 lub = 2.957922859e-26
+ uc = 1.218677263e-10 luc = -5.916673095e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.325369855e+05 lvsat = 1.597285411e-3
+ a0 = 1.499999999e+00 la0 = 1.571152097e-16
+ ags = 1.250000000e+00 lags = 3.363354040e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -6.898412508e-08 lb0 = 1.392658415e-14
+ b1 = 9.858632274e-11 lb1 = -1.990270542e-17
+ keta = -1.889316341e-01 lketa = 2.135570583e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.499568007e-01 lpclm = -2.248687870e-8
+ pdiblc1 = 3.569721502e-01 lpdiblc1 = -2.689404255e-17
+ pdiblc2 = 8.406112095e-03 lpdiblc2 = 7.211176101e-19
+ pdiblcb = -1.032957700e-01 lpdiblcb = 2.135180921e-18
+ drout = 5.033266589e-01 ldrout = 1.424531604e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 1.407623291e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 5.774280622e-09 lalpha0 = 3.194912098e-15
+ alpha1 = 0.85
+ beta0 = 1.518074234e+01 lbeta0 = -1.737675240e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.585636645e-01 lkt1 = 3.553695993e-9
+ kt2 = -2.887893901e-02 lkt2 = 8.536504836e-19
+ at = -1.837987011e+04 lat = 9.508667194e-3
+ ute = -1.325229293e+00 lute = 1.248854588e-9
+ ua1 = -2.384733722e-11 lua1 = 1.610621982e-25
+ ub1 = 7.077531683e-19 lub1 = 2.287943144e-34
+ uc1 = 1.471862500e-10 luc1 = -3.313685534e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.98 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {1.194873363e+01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.523958373e-06 wvth0 = -7.556472499e-06 pvth0 = 9.965551497e-13
+ k1 = 0.90707349
+ k2 = 9.875103659e-01 lk2 = -1.462520629e-07 wk2 = -7.922978880e-07 pk2 = 1.044890378e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.45863
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000021e-03 lcdscd = -2.765170037e-18 wcdscd = -1.339528488e-17 pcdscd = 1.766586877e-24
+ cit = 0.0
+ voff = {-2.075300001e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.193356525e-17
+ nfactor = 8.275710773e+00 lnfactor = -7.045628116e-07 wnfactor = -3.582793332e-06 pnfactor = 4.725023674e-13
+ eta0 = 8.801220094e-10 leta0 = -8.964436551e-17 weta0 = 5.138827172e-19 peta0 = -6.777136663e-26
+ etab = -0.043998
+ u0 = -8.291482853e-01 lu0 = 1.132834857e-07 wu0 = 5.756643738e-07 pu0 = -7.591919328e-14
+ ua = -1.238295196e-09 lua = 1.030710037e-17 wua = 5.241294305e-17 pua = -6.912271342e-24
+ ub = 4.818322194e-18 lub = -3.284513543e-25 wub = -1.670217761e-24 pub = 2.202699885e-31
+ uc = 7.700399988e-11 luc = 1.192049981e-26 wuc = 9.165161187e-28 puc = -1.209751646e-34
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -6.662743445e+05 lvsat = 1.069453224e-01 wvsat = 5.607202436e-01 pvsat = -7.394834644e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -8.178175521e-06 lb0 = 1.083374855e-12 wb0 = 5.509101732e-12 pb0 = -7.265458456e-19
+ b1 = 1.168756218e-08 lb1 = -1.548268431e-15 wb1 = -7.873145898e-15 pb1 = 1.038318354e-21
+ keta = -2.700000006e-02 lketa = 6.177169887e-18 wketa = -5.266898029e-19 pketa = 6.949996134e-26
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 9.696314183e-01 lpclm = -1.042101869e-07 wpclm = -5.299223250e-07 ppclm = 6.988668614e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.000000001e-08 lalpha0 = -1.169646621e-24 walpha0 = 1.053708986e-24 palpha0 = -1.389134033e-31
+ alpha1 = 0.85
+ beta0 = 1.091651628e+01 lbeta0 = 3.886028724e-07 wbeta0 = 1.976096043e-06 pbeta0 = -2.606095223e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -8.428655518e-02 lkt1 = -1.943014346e-08 wkt1 = -9.880480092e-08 pkt1 = 1.303047595e-14
+ kt2 = -0.028878939
+ at = 5.372048693e+04 lat = 6.960239261e-12 wat = 2.253800631e-13 pat = -2.980232239e-20
+ ute = -2.052414123e+00 lute = 9.715071713e-08 wute = 4.940240046e-07 pute = -6.515237975e-14
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.99 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {0.4913699+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56800772
+ k2 = -0.040590746
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 2.78042
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.025731
+ ua = -1.0529435e-9
+ ub = 1.832e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 9.1484e-8
+ b1 = 1.6098e-9
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.100 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.753697877e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.192323364e-7
+ k1 = 6.121972372e-01 lk1 = -8.816639883e-7
+ k2 = -5.732582613e-02 lk2 = 3.338963274e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.017062664e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.311152548e-7
+ nfactor = 2.999527454e+00 lnfactor = -4.371605856e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.399768874e-02 lu0 = 3.458282001e-8
+ ua = -1.240665649e-09 lua = 3.745409973e-15
+ ub = 1.951616170e-18 lub = -2.386567588e-24
+ uc = 6.326057033e-11 luc = -2.937629231e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.390829178e+00 la0 = -5.632251912e-7
+ ags = 3.209382116e-01 lags = 4.776837126e-07 wags = -8.881784197e-22
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 8.925150941e-08 lb0 = 4.454238660e-14
+ b1 = 2.167571440e-09 lb1 = -1.112858939e-14
+ keta = -2.666112675e-03 lketa = -3.751925933e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.631270000e-03 lpclm = 5.288499448e-07 ppclm = -4.440892099e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 5.528995573e-04 lpdiblc2 = 8.128953030e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -7.319501400e+07 lpscbe1 = 5.949551434e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.832257539e-01 lkt1 = -6.293314343e-8
+ kt2 = -3.544646383e-02 lkt2 = 1.182853816e-7
+ at = 1.981929862e+05 lat = -4.627437017e-1
+ ute = -1.016200285e+00 lute = -1.979220918e-6
+ ua1 = 1.030149760e-09 lua1 = 1.812633186e-15
+ ub1 = -3.832369470e-19 lub1 = -3.715699712e-24
+ uc1 = 6.920223587e-11 luc1 = -7.059748407e-16 wuc1 = -1.033975766e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.101 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.174342346e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.525913972e-8
+ k1 = 4.373408531e-01 lk1 = 5.087731700e-7
+ k2 = 8.934565372e-03 lk2 = -1.929984209e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.179994591e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.553724997e-9
+ nfactor = 1.644821634e+00 lnfactor = 6.400853618e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.718425420e-02 lu0 = 9.243630640e-9
+ ua = -9.777670666e-10 lua = 1.654871732e-15
+ ub = 1.840111304e-18 lub = -1.499894165e-24
+ uc = 9.701328365e-12 luc = 1.321337955e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.408917323e+00 la0 = -7.070599674e-7
+ ags = 3.610925198e-01 lags = 1.583814327e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 5.011079129e-08 lb0 = 3.557847194e-13
+ b1 = -1.658197099e-09 lb1 = 1.929346677e-14 pb1 = -1.323488980e-35
+ keta = -1.740241834e-02 lketa = 7.966208966e-08 wketa = 2.775557562e-23
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -6.899761706e-01 lpclm = 5.938871634e-06 wpclm = 4.440892099e-22 ppclm = 7.105427358e-27
+ pdiblc1 = 0.39
+ pdiblc2 = -1.623723774e-03 lpdiblc2 = 2.543720274e-08 ppdiblc2 = 2.775557562e-29
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.392309919e+08 lpscbe1 = 2.844246136e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.862989458e-01 lkt1 = -3.849548711e-8
+ kt2 = -9.860889619e-03 lkt2 = -8.516805990e-8
+ at = 140000.0
+ ute = -1.231212620e+00 lute = -2.694684098e-7
+ ua1 = 1.514330084e-09 lua1 = -2.037511139e-15
+ ub1 = -1.026378584e-18 lub1 = 1.398486053e-24
+ uc1 = -7.088796187e-11 luc1 = 4.080057410e-16 wuc1 = -1.033975766e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.102 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.258444758e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.849541224e-8
+ k1 = 5.592357205e-01 lk1 = 2.705915957e-8
+ k2 = -3.344055097e-02 lk2 = -2.553700375e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.527821500e-01 ldsub = -1.157040216e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.370079140e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 7.356542684e-8
+ nfactor = 3.198174774e+00 lnfactor = 2.621868556e-7
+ eta0 = 1.575872697e-01 leta0 = -3.066156572e-7
+ etab = -1.378278648e-01 letab = 2.680476500e-7
+ u0 = 2.961611194e-02 lu0 = -3.667817484e-10
+ ua = -7.010393526e-10 lua = 5.612767375e-16
+ ub = 1.754049020e-18 lub = -1.159786258e-24
+ uc = 3.566812735e-11 luc = 2.951609590e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.605932281e+00 la0 = -1.485639637e-6
+ ags = 3.277011992e-01 lags = 2.903399581e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 7.970976424e-08 lb0 = 2.388131005e-13
+ b1 = 8.033723719e-10 lb1 = 9.565637143e-15
+ keta = 5.453875497e-04 lketa = 8.734496589e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.112609403e+00 lpclm = -1.184732045e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.502894210e-03 lpdiblc2 = 9.129299537e-9
+ pdiblcb = -3.719925625e-02 lpdiblcb = 4.821000899e-8
+ drout = 0.56
+ pscbe1 = 6.245423126e+08 lpscbe1 = 3.424725263e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.591689679e-01 lkt1 = -1.457099312e-7
+ kt2 = -1.496516276e-02 lkt2 = -6.499657985e-8
+ at = 1.698930575e+05 lat = -1.181338060e-1
+ ute = -8.787696445e-01 lute = -1.662281110e-6
+ ua1 = 2.126322375e-09 lua1 = -4.456031847e-15
+ ub1 = -1.476118686e-18 lub1 = 3.175805416e-24
+ uc1 = 8.711055893e-12 luc1 = 9.343989506e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.103 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.784394203e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.403361498e-8
+ k1 = 5.910989287e-01 lk1 = -3.513403122e-8
+ k2 = -5.807107652e-02 lk2 = 2.253885108e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.26
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-6.567142512e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -6.567491050e-8
+ nfactor = 3.233958994e+00 lnfactor = 1.923403166e-7
+ eta0 = -1.433508281e-03 leta0 = 3.773978078e-09 weta0 = 1.734723476e-24
+ etab = 7.933901887e-02 letab = -1.558362640e-07 wetab = 1.214306433e-23 petab = 8.326672685e-29
+ u0 = 3.161666009e-02 lu0 = -4.271613666e-9
+ ua = 2.752158536e-10 lua = -1.344257251e-15
+ ub = 3.376251922e-19 lub = 1.604904499e-24
+ uc = 6.148628680e-11 luc = -2.087787897e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.674837450e+04 lvsat = 6.346786025e-3
+ a0 = 5.066918688e-01 la0 = 6.599468372e-7
+ ags = -2.598775475e-01 lags = 1.437223750e-06 pags = 1.776356839e-27
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.118978317e-07 lb0 = 1.759858233e-13
+ b1 = 4.226685500e-09 lb1 = 2.883737292e-15
+ keta = 6.946103312e-02 lketa = -1.257806426e-07 wketa = -5.551115123e-23 pketa = 2.775557562e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.584889993e-01 lpclm = 6.775974424e-7
+ pdiblc1 = 4.239170811e-01 lpdiblc1 = -6.620210620e-8
+ pdiblc2 = 9.545914571e-03 lpdiblc2 = -4.617838089e-09 wpdiblc2 = 2.775557562e-23
+ pdiblcb = -2.421622557e-02 lpdiblcb = 2.286867807e-8
+ drout = 2.176050537e-01 ldrout = 6.683141902e-7
+ pscbe1 = 8.629220470e+08 lpscbe1 = -1.228163479e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.195826690e-06 lalpha0 = 1.020019183e-11 walpha0 = 3.917527381e-27 palpha0 = -1.090554920e-32
+ alpha1 = 0.85
+ beta0 = 1.042942088e+01 lbeta0 = 6.696082211e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.901361166e-01 lkt1 = 1.099223579e-7
+ kt2 = -6.838621167e-02 lkt2 = 3.927495052e-8
+ at = 1.538056803e+05 lat = -8.673316007e-2
+ ute = -2.354634327e+00 lute = 1.218431122e-6
+ ua1 = -1.525599643e-09 lua1 = 2.672085355e-15 wua1 = -8.271806126e-31 pua1 = -8.271806126e-37
+ ub1 = 9.327016030e-19 lub1 = -1.525925138e-24 pub1 = -7.703719778e-46
+ uc1 = 7.140092441e-11 luc1 = -2.892326820e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.104 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.218486251e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.713217742e-9
+ k1 = 6.257710814e-01 lk1 = -6.813779454e-8
+ k2 = -5.325740349e-02 lk2 = 1.795680719e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.145343276e-01 ldsub = 4.327790972e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.265594373e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.716768537e-9
+ nfactor = 3.816562507e+00 lnfactor = -3.622288973e-7
+ eta0 = -4.380244825e-01 leta0 = 4.193566312e-07 weta0 = 2.775557562e-22 peta0 = 3.053113318e-28
+ etab = -1.600650675e-01 letab = 7.204793715e-8
+ u0 = 2.956204634e-02 lu0 = -2.315865879e-9
+ ua = -8.551569683e-10 lua = -2.682768386e-16
+ ub = 1.911412579e-18 lub = 1.068461874e-25
+ uc = 2.781855420e-11 luc = 1.116979601e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.498700947e+04 lvsat = 4.609863593e-2
+ a0 = 1.033165535e+00 la0 = 1.588065578e-7
+ ags = 2.238489687e+00 lags = -9.409245514e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 5.649984863e-07 lb0 = -2.553120810e-13
+ b1 = 1.381407783e-08 lb1 = -6.242319304e-15
+ keta = -1.128952678e-01 lketa = 4.780085550e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.248591510e+00 lpclm = -3.600504257e-7
+ pdiblc1 = 6.447801384e-01 lpdiblc1 = -2.764374541e-7
+ pdiblc2 = 8.895504641e-03 lpdiblc2 = -3.998725234e-9
+ pdiblcb = 8.513601992e-02 lpdiblcb = -8.122164671e-08 wpdiblcb = -7.806255642e-23 ppdiblcb = 7.719519468e-29
+ drout = 8.471347030e-01 ldrout = 6.907687805e-8
+ pscbe1 = 1.002269402e+09 lpscbe1 = -2.554584477e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 6.984094440e-06 lalpha0 = -1.393643679e-12
+ alpha1 = 0.85
+ beta0 = 1.696331585e+01 lbeta0 = 4.765917258e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.707775674e-01 lkt1 = -3.692777228e-9
+ kt2 = -1.845629469e-02 lkt2 = -8.252388786e-9
+ at = 1.097132702e+05 lat = -4.476243271e-2
+ ute = -8.616208324e-01 lute = -2.027400563e-7
+ ua1 = 1.688160728e-09 lua1 = -3.870320810e-16
+ ub1 = -7.051401785e-19 lub1 = 3.310533463e-26
+ uc1 = 7.289584949e-11 luc1 = -3.034625898e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.105 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.750340240e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.132025349e-8
+ k1 = 1.260614571e-01 lk1 = 1.576714902e-7
+ k2 = 8.475738853e-02 lk2 = -4.440945505e-08 pk2 = 4.163336342e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.905328527e-01 ldsub = 5.412372020e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.103590353e-03 lcdscd = -1.221701112e-9
+ cit = 0.0
+ voff = {-1.154994111e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.271458427e-8
+ nfactor = 3.206634077e+00 lnfactor = -8.661382834e-8
+ eta0 = 8.851262253e-01 leta0 = -1.785500338e-7
+ etab = 3.439973846e-02 letab = -1.582701384e-08 wetab = -1.040834086e-23 petab = -2.602085214e-30
+ u0 = 2.025864782e-02 lu0 = 1.888163151e-9
+ ua = -1.664072323e-09 lua = 9.725664082e-17
+ ub = 2.065347559e-18 lub = 3.728589477e-26
+ uc = 2.021746693e-11 luc = 1.460458292e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.342184647e+05 lvsat = 1.257826697e-3
+ a0 = 1.291411731e+00 la0 = 4.211000822e-8
+ ags = -7.269793732e-01 lags = 3.991145728e-07 pags = 3.330669074e-28
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.316735352e-16 lb0 = -2.658238496e-23
+ b1 = -6.482321705e-18 lb1 = 1.308657588e-24
+ keta = 5.428652146e-02 lketa = -2.774541862e-08 pketa = 6.938893904e-30
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.240064173e-01 lpclm = -7.781228934e-8
+ pdiblc1 = -2.285578198e-01 lpdiblc1 = 1.182073759e-07 wpdiblc1 = -1.110223025e-22 ppdiblc1 = -8.326672685e-29
+ pdiblc2 = -6.704200072e-03 lpdiblc2 = 3.050484931e-09 wpdiblc2 = -1.084202172e-24 ppdiblc2 = -1.870248748e-30
+ pdiblcb = -8.758737421e-02 lpdiblcb = -3.171226653e-9
+ drout = 1.401075462e+00 ldrout = -1.812384259e-7
+ pscbe1 = 1.507016608e+08 lpscbe1 = 1.293488348e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.031901082e-06 lalpha0 = -1.415246593e-12
+ alpha1 = 0.85
+ beta0 = 2.100422375e+01 lbeta0 = -1.349417775e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.096264800e-01 lkt1 = 1.386230826e-8
+ kt2 = -4.304931441e-02 lkt2 = 2.860729557e-9
+ at = -3.932844299e+03 lat = 6.592087176e-3
+ ute = -1.303201518e+00 lute = -3.198134688e-9
+ ua1 = 1.522520005e-09 lua1 = -3.121821852e-16
+ ub1 = -1.713664128e-18 lub1 = 4.888381454e-25 pub1 = -3.851859889e-46
+ uc1 = -1.084804678e-10 luc1 = 5.161425266e-17 wuc1 = -5.169878828e-32 puc1 = 2.261821987e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.106 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {6.130803429e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.900108240e-8
+ k1 = 9.070734896e-01 lk1 = 5.142908321e-17
+ k2 = -1.611477193e-01 lk2 = 5.234114019e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -7.795097900e-18
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999996e-03 lcdscd = 5.442070405e-19
+ cit = 0.0
+ voff = {-1.237493848e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.104907131e-8
+ nfactor = 2.484263783e+00 lnfactor = 5.921900879e-8
+ eta0 = 2.001909455e-03 leta0 = -2.640137943e-10
+ etab = -4.399800002e-02 letab = 2.220557072e-18
+ u0 = 2.919169366e-02 lu0 = 8.475092343e-11
+ ua = -1.224106221e-09 lua = 8.435844238e-18
+ ub = 2.103521860e-18 lub = 2.957922859e-26
+ uc = 1.218677263e-10 luc = -5.916673095e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.325369855e+05 lvsat = 1.597285411e-3
+ a0 = 1.499999999e+00 la0 = 1.571063279e-16
+ ags = 1.250000000e+00 lags = 3.363709311e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -6.898412508e-08 lb0 = 1.392658415e-14
+ b1 = 9.858632274e-11 lb1 = -1.990270542e-17
+ keta = -1.889316341e-01 lketa = 2.135570583e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.499568007e-01 lpclm = -2.248687870e-8
+ pdiblc1 = 3.569721502e-01 lpdiblc1 = -2.689581891e-17
+ pdiblc2 = 8.406112095e-03 lpdiblc2 = 7.211453656e-19
+ pdiblcb = -1.032957700e-01 lpdiblcb = 2.135291943e-18
+ drout = 5.033266589e-01 ldrout = 1.424531604e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 1.407337189e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 5.774280622e-09 lalpha0 = 3.194912098e-15
+ alpha1 = 0.85
+ beta0 = 1.518074234e+01 lbeta0 = -1.737675240e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.585636645e-01 lkt1 = 3.553695993e-9
+ kt2 = -2.887893901e-02 lkt2 = 8.535949725e-19
+ at = -1.837987011e+04 lat = 9.508667194e-3
+ ute = -1.325229293e+00 lute = 1.248854588e-9
+ ua1 = -2.384733722e-11 lua1 = 1.610623275e-25
+ ub1 = 7.077531683e-19 lub1 = 2.287966255e-34
+ uc1 = 1.471862500e-10 luc1 = -3.312858353e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.107 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {-3.880355590e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.635977419e-07 wvth0 = 2.900730368e-06 pvth0 = -3.825512216e-13
+ k1 = 0.90707349
+ k2 = -6.061728085e-01 lk2 = 6.392446782e-08 wk2 = 2.605402149e-07 pk2 = -3.436030408e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.585249057e-01 ldsub = 1.385994477e-11 wdsub = 6.942867459e-11 pdsub = -9.156323034e-18
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000001e-03 lcdscd = -9.109032972e-20
+ cit = 0.0
+ voff = {-2.075300001e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.193223298e-17
+ nfactor = 6.715065360e+00 lnfactor = -4.987433340e-07 wnfactor = -2.551781032e-06 pnfactor = 3.365314343e-13
+ eta0 = 1.494627088e-02 leta0 = -1.971128926e-09 weta0 = -9.873983253e-09 peta0 = 1.302190785e-15
+ etab = -0.043998
+ u0 = 1.684154364e-01 lu0 = -1.827621550e-08 wu0 = -8.335814279e-08 pu0 = 1.099335523e-14
+ ua = 1.137846112e-09 lua = -3.030607914e-16 wua = -1.517342041e-15 pua = 2.001085858e-22
+ ub = -2.380164850e-18 lub = 6.208923157e-25 wub = 3.085333133e-24 pub = -4.068968189e-31
+ uc = 3.003892365e-10 luc = -2.946026837e-17 wuc = -1.475754356e-16 puc = 1.946239602e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.928588791e+05 lvsat = -1.954612624e-02 wvsat = -7.291385621e-02 pvsat = 9.615952271e-9
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.002439095e-05 lb0 = -1.317197815e-12 wb0 = -6.516096164e-12 pb0 = 8.593492782e-19
+ b1 = 3.616590999e-07 lb1 = -4.770286479e-14 wb1 = -2.390755428e-13 pb1 = 3.152952166e-20
+ keta = -2.700000006e-02 lketa = 6.282308007e-18
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.545414356e-01 lpclm = 5.723495320e-08 wpclm = 2.788054358e-07 ppclm = -3.676913968e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.000000001e-08 lalpha0 = -1.379975490e-24
+ alpha1 = 0.85
+ beta0 = 1.390773688e+01 lbeta0 = -5.882290701e-9
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.491681706e-01 lkt1 = 2.869080887e-08 wkt1 = 1.422476705e-07 pkt1 = -1.875976503e-14
+ kt2 = -0.028878939
+ at = 5.372048693e+04 lat = 6.915419362e-12
+ ute = 5.697718714e-02 lute = -1.810379182e-07 wute = -8.995073951e-07 pute = 1.186279348e-13
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.108 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {0.4913699+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56800772
+ k2 = -0.040590746
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 2.78042
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.025731
+ ua = -1.0529435e-9
+ ub = 1.832e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 9.1484e-8
+ b1 = 1.6098e-9
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.109 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.753697877e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.192323364e-7
+ k1 = 6.121972372e-01 lk1 = -8.816639883e-7
+ k2 = -5.732582613e-02 lk2 = 3.338963274e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.017062664e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.311152548e-7
+ nfactor = 2.999527454e+00 lnfactor = -4.371605856e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.399768874e-02 lu0 = 3.458282001e-8
+ ua = -1.240665649e-09 lua = 3.745409973e-15
+ ub = 1.951616170e-18 lub = -2.386567588e-24
+ uc = 6.326057033e-11 luc = -2.937629231e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.390829178e+00 la0 = -5.632251912e-7
+ ags = 3.209382116e-01 lags = 4.776837126e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 8.925150941e-08 lb0 = 4.454238660e-14
+ b1 = 2.167571440e-09 lb1 = -1.112858939e-14
+ keta = -2.666112675e-03 lketa = -3.751925933e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.631270000e-03 lpclm = 5.288499448e-07 ppclm = 1.776356839e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 5.528995573e-04 lpdiblc2 = 8.128953030e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -7.319501400e+07 lpscbe1 = 5.949551434e+03 ppscbe1 = -1.525878906e-17
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.832257539e-01 lkt1 = -6.293314343e-8
+ kt2 = -3.544646383e-02 lkt2 = 1.182853816e-07 wkt2 = 2.220446049e-22
+ at = 1.981929862e+05 lat = -4.627437017e-1
+ ute = -1.016200285e+00 lute = -1.979220918e-6
+ ua1 = 1.030149760e-09 lua1 = 1.812633186e-15
+ ub1 = -3.832369470e-19 lub1 = -3.715699712e-24
+ uc1 = 6.920223587e-11 luc1 = -7.059748407e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.110 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.174342346e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.525913972e-8
+ k1 = 4.373408531e-01 lk1 = 5.087731700e-7
+ k2 = 8.934565372e-03 lk2 = -1.929984209e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.179994591e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.553724997e-9
+ nfactor = 1.644821634e+00 lnfactor = 6.400853618e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.718425420e-02 lu0 = 9.243630640e-9
+ ua = -9.777670666e-10 lua = 1.654871732e-15
+ ub = 1.840111304e-18 lub = -1.499894165e-24
+ uc = 9.701328365e-12 luc = 1.321337955e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.408917322e+00 la0 = -7.070599674e-7
+ ags = 3.610925198e-01 lags = 1.583814327e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 5.011079129e-08 lb0 = 3.557847194e-13
+ b1 = -1.658197099e-09 lb1 = 1.929346677e-14 pb1 = 2.646977960e-35
+ keta = -1.740241834e-02 lketa = 7.966208966e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -6.899761706e-01 lpclm = 5.938871634e-06 ppclm = 1.065814104e-26
+ pdiblc1 = 0.39
+ pdiblc2 = -1.623723774e-03 lpdiblc2 = 2.543720274e-08 ppdiblc2 = -5.551115123e-29
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.392309919e+08 lpscbe1 = 2.844246136e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.862989458e-01 lkt1 = -3.849548711e-8
+ kt2 = -9.860889619e-03 lkt2 = -8.516805990e-8
+ at = 140000.0
+ ute = -1.231212620e+00 lute = -2.694684098e-7
+ ua1 = 1.514330084e-09 lua1 = -2.037511139e-15
+ ub1 = -1.026378584e-18 lub1 = 1.398486053e-24
+ uc1 = -7.088796187e-11 luc1 = 4.080057410e-16 puc1 = 8.271806126e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.111 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.258444758e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.849541224e-8
+ k1 = 5.592357205e-01 lk1 = 2.705915957e-8
+ k2 = -3.344055097e-02 lk2 = -2.553700375e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.527821500e-01 ldsub = -1.157040216e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.370079140e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 7.356542684e-8
+ nfactor = 3.198174774e+00 lnfactor = 2.621868556e-7
+ eta0 = 1.575872697e-01 leta0 = -3.066156572e-7
+ etab = -1.378278648e-01 letab = 2.680476500e-7
+ u0 = 2.961611194e-02 lu0 = -3.667817484e-10
+ ua = -7.010393526e-10 lua = 5.612767375e-16
+ ub = 1.754049020e-18 lub = -1.159786258e-24
+ uc = 3.566812735e-11 luc = 2.951609590e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.605932281e+00 la0 = -1.485639637e-6
+ ags = 3.277011992e-01 lags = 2.903399581e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 7.970976424e-08 lb0 = 2.388131005e-13
+ b1 = 8.033723719e-10 lb1 = 9.565637143e-15
+ keta = 5.453875496e-04 lketa = 8.734496589e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.112609403e+00 lpclm = -1.184732045e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.502894210e-03 lpdiblc2 = 9.129299537e-9
+ pdiblcb = -3.719925625e-02 lpdiblcb = 4.821000899e-8
+ drout = 0.56
+ pscbe1 = 6.245423126e+08 lpscbe1 = 3.424725263e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.591689679e-01 lkt1 = -1.457099312e-7
+ kt2 = -1.496516276e-02 lkt2 = -6.499657985e-8
+ at = 1.698930575e+05 lat = -1.181338060e-1
+ ute = -8.787696445e-01 lute = -1.662281110e-6
+ ua1 = 2.126322375e-09 lua1 = -4.456031847e-15
+ ub1 = -1.476118686e-18 lub1 = 3.175805416e-24 wub1 = -6.162975822e-39
+ uc1 = 8.711055893e-12 luc1 = 9.343989506e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.112 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.784394203e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.403361498e-8
+ k1 = 5.910989287e-01 lk1 = -3.513403122e-8
+ k2 = -5.807107652e-02 lk2 = 2.253885108e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.26
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-6.567142512e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -6.567491050e-8
+ nfactor = 3.233958994e+00 lnfactor = 1.923403166e-7
+ eta0 = -1.433508281e-03 leta0 = 3.773978078e-09 peta0 = -6.938893904e-30
+ etab = 7.933901888e-02 letab = -1.558362640e-07 wetab = -5.551115123e-23 petab = 1.179611964e-28
+ u0 = 3.161666009e-02 lu0 = -4.271613666e-9
+ ua = 2.752158536e-10 lua = -1.344257251e-15
+ ub = 3.376251922e-19 lub = 1.604904499e-24
+ uc = 6.148628680e-11 luc = -2.087787897e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.674837450e+04 lvsat = 6.346786025e-3
+ a0 = 5.066918688e-01 la0 = 6.599468372e-7
+ ags = -2.598775476e-01 lags = 1.437223750e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.118978317e-07 lb0 = 1.759858233e-13
+ b1 = 4.226685500e-09 lb1 = 2.883737292e-15
+ keta = 6.946103312e-02 lketa = -1.257806426e-07 wketa = 5.551115123e-23 pketa = -1.665334537e-28
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.584889993e-01 lpclm = 6.775974424e-7
+ pdiblc1 = 4.239170811e-01 lpdiblc1 = -6.620210620e-8
+ pdiblc2 = 9.545914571e-03 lpdiblc2 = -4.617838089e-9
+ pdiblcb = -2.421622557e-02 lpdiblcb = 2.286867807e-8
+ drout = 2.176050537e-01 ldrout = 6.683141902e-7
+ pscbe1 = 8.629220470e+08 lpscbe1 = -1.228163479e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.195826690e-06 lalpha0 = 1.020019183e-11 walpha0 = 1.101142831e-26 palpha0 = 2.117582368e-33
+ alpha1 = 0.85
+ beta0 = 1.042942088e+01 lbeta0 = 6.696082211e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.901361166e-01 lkt1 = 1.099223579e-7
+ kt2 = -6.838621167e-02 lkt2 = 3.927495052e-8
+ at = 1.538056803e+05 lat = -8.673316007e-2
+ ute = -2.354634327e+00 lute = 1.218431122e-6
+ ua1 = -1.525599643e-09 lua1 = 2.672085355e-15 wua1 = 1.654361225e-30 pua1 = 4.963083675e-36
+ ub1 = 9.327016030e-19 lub1 = -1.525925138e-24 wub1 = 1.540743956e-39 pub1 = 4.622231867e-45
+ uc1 = 7.140092441e-11 luc1 = -2.892326820e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.113 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.218486251e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.713217742e-9
+ k1 = 6.257710814e-01 lk1 = -6.813779454e-8
+ k2 = -5.325740349e-02 lk2 = 1.795680719e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.145343276e-01 ldsub = 4.327790972e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.265594373e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.716768537e-9
+ nfactor = 3.816562507e+00 lnfactor = -3.622288973e-7
+ eta0 = -4.380244825e-01 leta0 = 4.193566312e-07 weta0 = -9.992007222e-22 peta0 = -1.720845688e-27
+ etab = -1.600650675e-01 letab = 7.204793715e-8
+ u0 = 2.956204634e-02 lu0 = -2.315865879e-9
+ ua = -8.551569683e-10 lua = -2.682768386e-16
+ ub = 1.911412579e-18 lub = 1.068461874e-25
+ uc = 2.781855420e-11 luc = 1.116979601e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.498700947e+04 lvsat = 4.609863593e-2
+ a0 = 1.033165535e+00 la0 = 1.588065578e-7
+ ags = 2.238489687e+00 lags = -9.409245514e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 5.649984863e-07 lb0 = -2.553120810e-13
+ b1 = 1.381407783e-08 lb1 = -6.242319304e-15
+ keta = -1.128952678e-01 lketa = 4.780085550e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.248591510e+00 lpclm = -3.600504257e-7
+ pdiblc1 = 6.447801384e-01 lpdiblc1 = -2.764374541e-7
+ pdiblc2 = 8.895504641e-03 lpdiblc2 = -3.998725234e-9
+ pdiblcb = 8.513601992e-02 lpdiblcb = -8.122164671e-08 wpdiblcb = 3.469446952e-24 ppdiblcb = 1.023486851e-28
+ drout = 8.471347030e-01 ldrout = 6.907687805e-8
+ pscbe1 = 1.002269402e+09 lpscbe1 = -2.554584477e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 6.984094440e-06 lalpha0 = -1.393643679e-12
+ alpha1 = 0.85
+ beta0 = 1.696331585e+01 lbeta0 = 4.765917258e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.707775674e-01 lkt1 = -3.692777228e-9
+ kt2 = -1.845629469e-02 lkt2 = -8.252388786e-9
+ at = 1.097132702e+05 lat = -4.476243271e-2
+ ute = -8.616208324e-01 lute = -2.027400563e-7
+ ua1 = 1.688160728e-09 lua1 = -3.870320810e-16
+ ub1 = -7.051401785e-19 lub1 = 3.310533463e-26
+ uc1 = 7.289584949e-11 luc1 = -3.034625898e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.114 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.750340240e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.132025349e-8
+ k1 = 1.260614571e-01 lk1 = 1.576714902e-7
+ k2 = 8.475738853e-02 lk2 = -4.440945505e-08 wk2 = -1.110223025e-22 pk2 = -8.326672685e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.905328527e-01 ldsub = 5.412372020e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.103590353e-03 lcdscd = -1.221701112e-9
+ cit = 0.0
+ voff = {-1.154994111e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.271458427e-8
+ nfactor = 3.206634077e+00 lnfactor = -8.661382834e-8
+ eta0 = 8.851262253e-01 leta0 = -1.785500338e-7
+ etab = 3.439973846e-02 letab = -1.582701384e-08 wetab = -5.551115123e-23 petab = 5.377642776e-29
+ u0 = 2.025864782e-02 lu0 = 1.888163151e-9
+ ua = -1.664072323e-09 lua = 9.725664082e-17
+ ub = 2.065347559e-18 lub = 3.728589477e-26
+ uc = 2.021746693e-11 luc = 1.460458292e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.342184647e+05 lvsat = 1.257826697e-3
+ a0 = 1.291411731e+00 la0 = 4.211000822e-8
+ ags = -7.269793732e-01 lags = 3.991145728e-07 wags = -1.776356839e-21
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.316735352e-16 lb0 = -2.658238496e-23
+ b1 = -6.482321705e-18 lb1 = 1.308657588e-24
+ keta = 5.428652146e-02 lketa = -2.774541862e-08 wketa = -2.220446049e-22 pketa = 6.938893904e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.240064173e-01 lpclm = -7.781228934e-8
+ pdiblc1 = -2.285578198e-01 lpdiblc1 = 1.182073759e-07 wpdiblc1 = -4.440892099e-22 ppdiblc1 = -1.665334537e-28
+ pdiblc2 = -6.704200072e-03 lpdiblc2 = 3.050484931e-09 wpdiblc2 = 2.515349040e-23 ppdiblc2 = -1.192622390e-30
+ pdiblcb = -8.758737421e-02 lpdiblcb = -3.171226653e-9
+ drout = 1.401075462e+00 ldrout = -1.812384259e-7
+ pscbe1 = 1.507016608e+08 lpscbe1 = 1.293488348e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.031901082e-06 lalpha0 = -1.415246593e-12
+ alpha1 = 0.85
+ beta0 = 2.100422375e+01 lbeta0 = -1.349417775e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.096264800e-01 lkt1 = 1.386230826e-8
+ kt2 = -4.304931441e-02 lkt2 = 2.860729557e-9
+ at = -3.932844299e+03 lat = 6.592087176e-3
+ ute = -1.303201518e+00 lute = -3.198134688e-9
+ ua1 = 1.522520005e-09 lua1 = -3.121821852e-16
+ ub1 = -1.713664128e-18 lub1 = 4.888381454e-25
+ uc1 = -1.084804678e-10 luc1 = 5.161425266e-17 wuc1 = -4.135903063e-31 puc1 = 1.421716678e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.115 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {6.130803429e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.900108240e-8
+ k1 = 9.070734896e-01 lk1 = 5.142908321e-17
+ k2 = -1.611477193e-01 lk2 = 5.234114019e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -7.794653811e-18
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999996e-03 lcdscd = 5.442105100e-19
+ cit = 0.0
+ voff = {-1.237493848e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.104907131e-8
+ nfactor = 2.484263783e+00 lnfactor = 5.921900879e-8
+ eta0 = 2.001909455e-03 leta0 = -2.640137943e-10
+ etab = -4.399800002e-02 letab = 2.220668094e-18
+ u0 = 2.919169366e-02 lu0 = 8.475092343e-11
+ ua = -1.224106221e-09 lua = 8.435844238e-18
+ ub = 2.103521860e-18 lub = 2.957922859e-26
+ uc = 1.218677263e-10 luc = -5.916673095e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.325369855e+05 lvsat = 1.597285411e-3
+ a0 = 1.499999999e+00 la0 = 1.571081043e-16
+ ags = 1.250000000e+00 lags = 3.363354040e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -6.898412508e-08 lb0 = 1.392658415e-14
+ b1 = 9.858632274e-11 lb1 = -1.990270542e-17
+ keta = -1.889316341e-01 lketa = 2.135570583e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.499568007e-01 lpclm = -2.248687870e-8
+ pdiblc1 = 3.569721502e-01 lpdiblc1 = -2.689759526e-17
+ pdiblc2 = 8.406112095e-03 lpdiblc2 = 7.211453656e-19
+ pdiblcb = -1.032957700e-01 lpdiblcb = 2.135180921e-18
+ drout = 5.033266589e-01 ldrout = 1.424531604e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 1.407241821e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 5.774280622e-09 lalpha0 = 3.194912098e-15
+ alpha1 = 0.85
+ beta0 = 1.518074234e+01 lbeta0 = -1.737675240e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.585636645e-01 lkt1 = 3.553695993e-9
+ kt2 = -2.887893901e-02 lkt2 = 8.536504836e-19
+ at = -1.837987011e+04 lat = 9.508667194e-3
+ ute = -1.325229293e+00 lute = 1.248854588e-9
+ ua1 = -2.384733722e-11 lua1 = 1.610621982e-25
+ ub1 = 7.077531683e-19 lub1 = 2.287973959e-34
+ uc1 = 1.471862500e-10 luc1 = -3.312858353e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.116 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {7.086112022e-02+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.250733090e-08 wvth0 = 4.089666711e-07 pvth0 = -5.393493355e-14
+ k1 = 0.90707349
+ k2 = -1.561746687e-01 lk2 = 4.578263143e-09 wk2 = -2.324301201e-08 pk2 = 3.065311667e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.585241313e-01 ldsub = 1.396207225e-11 wdsub = 6.991703044e-11 pdsub = -9.220727893e-18
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000001e-03 lcdscd = -9.108686028e-20
+ cit = 0.0
+ voff = {-2.075300001e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.193267707e-17
+ nfactor = 6.715065591e+00 lnfactor = -4.987433644e-07 wnfactor = -2.551781177e-06 pnfactor = 3.365314534e-13
+ eta0 = 1.494623607e-02 leta0 = -1.971124532e-09 weta0 = -9.873962242e-09 peta0 = 1.302188014e-15
+ etab = -0.043998
+ u0 = -1.320960968e-01 lu0 = 2.135554602e-08 wu0 = 1.061540464e-07 pu0 = -1.399970180e-14
+ ua = 1.137850984e-09 lua = -3.030614339e-16 wua = -1.517345114e-15 pua = 2.001089909e-22
+ ub = -2.380311201e-18 lub = 6.209116165e-25 wub = 3.085425426e-24 pub = -4.069089906e-31
+ uc = 3.020282860e-10 luc = -2.967642787e-17 wuc = -1.486090727e-16 puc = 1.959871312e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.689527288e+05 lvsat = -1.639335923e-02 wvsat = -5.783787281e-02 pvsat = 7.627716504e-9
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.002426040e-05 lb0 = -1.317180597e-12 wb0 = -6.516013832e-12 pb0 = 8.593384202e-19
+ b1 = 3.616598576e-07 lb1 = -4.770296472e-14 wb1 = -2.390760206e-13 pb1 = 3.152958468e-20
+ keta = -2.700000006e-02 lketa = 6.282308007e-18
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.545414263e-01 lpclm = 5.723495198e-08 wpclm = 2.788054300e-07 ppclm = -3.676913891e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.000000001e-08 lalpha0 = -1.379922550e-24
+ alpha1 = 0.85
+ beta0 = 1.390773688e+01 lbeta0 = -5.882290701e-9
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.491681634e-01 lkt1 = 2.869080791e-08 wkt1 = 1.422476659e-07 pkt1 = -1.875976443e-14
+ kt2 = -0.028878939
+ at = 5.372048693e+04 lat = 6.915302947e-12
+ ute = 6.696761924e-02 lute = -1.823554664e-07 wute = -9.058076813e-07 pute = 1.194588228e-13
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.117 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {0.4913699+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56800772
+ k2 = -0.040590746
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 2.78042
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.025731
+ ua = -1.0529435e-9
+ ub = 1.832e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 9.1484e-8
+ b1 = 1.6098e-9
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.118 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.753697877e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.192323364e-7
+ k1 = 6.121972372e-01 lk1 = -8.816639883e-7
+ k2 = -5.732582613e-02 lk2 = 3.338963274e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.017062664e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.311152548e-7
+ nfactor = 2.999527454e+00 lnfactor = -4.371605856e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.399768874e-02 lu0 = 3.458282001e-8
+ ua = -1.240665649e-09 lua = 3.745409973e-15
+ ub = 1.951616170e-18 lub = -2.386567588e-24
+ uc = 6.326057033e-11 luc = -2.937629231e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.390829178e+00 la0 = -5.632251912e-7
+ ags = 3.209382116e-01 lags = 4.776837126e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 8.925150941e-08 lb0 = 4.454238660e-14
+ b1 = 2.167571440e-09 lb1 = -1.112858939e-14
+ keta = -2.666112675e-03 lketa = -3.751925933e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.631270000e-03 lpclm = 5.288499448e-07 ppclm = 8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 5.528995573e-04 lpdiblc2 = 8.128953030e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -7.319501400e+07 lpscbe1 = 5.949551434e+03 ppscbe1 = 7.629394531e-18
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.832257539e-01 lkt1 = -6.293314343e-8
+ kt2 = -3.544646383e-02 lkt2 = 1.182853816e-7
+ at = 1.981929863e+05 lat = -4.627437017e-1
+ ute = -1.016200285e+00 lute = -1.979220918e-6
+ ua1 = 1.030149760e-09 lua1 = 1.812633186e-15
+ ub1 = -3.832369470e-19 lub1 = -3.715699712e-24
+ uc1 = 6.920223587e-11 luc1 = -7.059748407e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.119 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.174342346e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.525913972e-8
+ k1 = 4.373408531e-01 lk1 = 5.087731700e-7
+ k2 = 8.934565372e-03 lk2 = -1.929984209e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.179994591e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.553724997e-9
+ nfactor = 1.644821634e+00 lnfactor = 6.400853618e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.718425420e-02 lu0 = 9.243630640e-9
+ ua = -9.777670666e-10 lua = 1.654871732e-15
+ ub = 1.840111304e-18 lub = -1.499894165e-24
+ uc = 9.701328365e-12 luc = 1.321337955e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.408917323e+00 la0 = -7.070599674e-7
+ ags = 3.610925198e-01 lags = 1.583814327e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 5.011079129e-08 lb0 = 3.557847194e-13
+ b1 = -1.658197099e-09 lb1 = 1.929346677e-14
+ keta = -1.740241834e-02 lketa = 7.966208966e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -6.899761706e-01 lpclm = 5.938871634e-06 ppclm = -1.776356839e-27
+ pdiblc1 = 0.39
+ pdiblc2 = -1.623723774e-03 lpdiblc2 = 2.543720274e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.392309919e+08 lpscbe1 = 2.844246136e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.862989458e-01 lkt1 = -3.849548711e-8
+ kt2 = -9.860889619e-03 lkt2 = -8.516805990e-8
+ at = 140000.0
+ ute = -1.231212620e+00 lute = -2.694684098e-7
+ ua1 = 1.514330084e-09 lua1 = -2.037511139e-15
+ ub1 = -1.026378584e-18 lub1 = 1.398486053e-24
+ uc1 = -7.088796187e-11 luc1 = 4.080057410e-16 wuc1 = -1.033975766e-31 puc1 = 4.135903063e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.120 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.258444758e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.849541224e-8
+ k1 = 5.592357205e-01 lk1 = 2.705915957e-8
+ k2 = -3.344055097e-02 lk2 = -2.553700375e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.527821500e-01 ldsub = -1.157040216e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.370079140e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 7.356542684e-8
+ nfactor = 3.198174774e+00 lnfactor = 2.621868556e-7
+ eta0 = 1.575872698e-01 leta0 = -3.066156572e-7
+ etab = -1.378278648e-01 letab = 2.680476500e-7
+ u0 = 2.961611194e-02 lu0 = -3.667817484e-10
+ ua = -7.010393526e-10 lua = 5.612767375e-16
+ ub = 1.754049020e-18 lub = -1.159786258e-24
+ uc = 3.566812735e-11 luc = 2.951609590e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.605932281e+00 la0 = -1.485639637e-6
+ ags = 3.277011992e-01 lags = 2.903399581e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 7.970976424e-08 lb0 = 2.388131005e-13
+ b1 = 8.033723719e-10 lb1 = 9.565637143e-15
+ keta = 5.453875497e-04 lketa = 8.734496589e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.112609403e+00 lpclm = -1.184732045e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.502894210e-03 lpdiblc2 = 9.129299537e-9
+ pdiblcb = -3.719925625e-02 lpdiblcb = 4.821000899e-8
+ drout = 0.56
+ pscbe1 = 6.245423126e+08 lpscbe1 = 3.424725263e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.591689679e-01 lkt1 = -1.457099312e-7
+ kt2 = -1.496516276e-02 lkt2 = -6.499657985e-8
+ at = 1.698930575e+05 lat = -1.181338060e-1
+ ute = -8.787696445e-01 lute = -1.662281110e-6
+ ua1 = 2.126322375e-09 lua1 = -4.456031847e-15
+ ub1 = -1.476118686e-18 lub1 = 3.175805416e-24
+ uc1 = 8.711055893e-12 luc1 = 9.343989506e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.121 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.784394203e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.403361498e-8
+ k1 = 5.910989287e-01 lk1 = -3.513403122e-8
+ k2 = -5.807107652e-02 lk2 = 2.253885108e-08 wk2 = 2.220446049e-22
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.26
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-6.567142512e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -6.567491050e-8
+ nfactor = 3.233958994e+00 lnfactor = 1.923403166e-7
+ eta0 = -1.433508281e-03 leta0 = 3.773978078e-09 peta0 = 3.469446952e-30
+ etab = 7.933901887e-02 letab = -1.558362640e-07 wetab = 3.469446952e-23 petab = -1.838806885e-28
+ u0 = 3.161666009e-02 lu0 = -4.271613666e-9
+ ua = 2.752158536e-10 lua = -1.344257251e-15 pua = -1.654361225e-36
+ ub = 3.376251922e-19 lub = 1.604904499e-24
+ uc = 6.148628680e-11 luc = -2.087787897e-17 wuc = -2.067951531e-31
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.674837450e+04 lvsat = 6.346786025e-3
+ a0 = 5.066918688e-01 la0 = 6.599468372e-7
+ ags = -2.598775475e-01 lags = 1.437223750e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.118978317e-07 lb0 = 1.759858233e-13
+ b1 = 4.226685500e-09 lb1 = 2.883737292e-15
+ keta = 6.946103312e-02 lketa = -1.257806426e-07 wketa = -2.775557562e-23 pketa = 1.387778781e-28
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.584889993e-01 lpclm = 6.775974424e-7
+ pdiblc1 = 4.239170811e-01 lpdiblc1 = -6.620210620e-8
+ pdiblc2 = 9.545914571e-03 lpdiblc2 = -4.617838089e-9
+ pdiblcb = -2.421622557e-02 lpdiblcb = 2.286867807e-8
+ drout = 2.176050537e-01 ldrout = 6.683141902e-7
+ pscbe1 = 8.629220470e+08 lpscbe1 = -1.228163479e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.195826690e-06 lalpha0 = 1.020019183e-11 walpha0 = -4.446922973e-27 palpha0 = 5.505714157e-33
+ alpha1 = 0.85
+ beta0 = 1.042942088e+01 lbeta0 = 6.696082211e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.901361166e-01 lkt1 = 1.099223579e-7
+ kt2 = -6.838621167e-02 lkt2 = 3.927495052e-8
+ at = 1.538056803e+05 lat = -8.673316007e-2
+ ute = -2.354634327e+00 lute = 1.218431122e-6
+ ua1 = -1.525599643e-09 lua1 = 2.672085355e-15 wua1 = -8.271806126e-31 pua1 = -1.654361225e-36
+ ub1 = 9.327016030e-19 lub1 = -1.525925138e-24 pub1 = -2.311115933e-45
+ uc1 = 7.140092441e-11 luc1 = -2.892326820e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.122 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {7.657712718e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.294721152e-07 wvth0 = -1.513862001e-07 pvth0 = 1.441016475e-13
+ k1 = 6.257710822e-01 lk1 = -6.813779531e-08 wk1 = -5.009823667e-16 pk1 = 4.768754280e-22
+ k2 = 4.737212088e-02 lk2 = -7.783052510e-08 wk2 = -6.245390297e-08 pk2 = 5.944868361e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.145343278e-01 ldsub = 4.327790950e-08 wdsub = -1.477626910e-16 pdsub = 1.406528227e-22
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.265594364e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.716769472e-09 wvoff = -6.095808303e-16 pvoff = 5.802482939e-22
+ nfactor = 3.816562516e+00 lnfactor = -3.622289064e-07 wnfactor = -5.922814239e-15 pnfactor = 5.637822653e-21
+ eta0 = -4.380244830e-01 leta0 = 4.193566317e-07 weta0 = 3.380755953e-16 peta0 = -3.218079622e-22
+ etab = -1.600650676e-01 letab = 7.204793725e-08 wetab = 6.792655327e-17 petab = -6.465783464e-23
+ u0 = -1.362103671e-02 lu0 = 3.878929040e-08 wu0 = 2.680080320e-08 pu0 = -2.551117535e-14
+ ua = -8.551569649e-10 lua = -2.682768418e-16 wua = -2.129189366e-24 pua = 2.026731467e-30
+ ub = 1.911407154e-18 lub = 1.068513516e-25 wub = 3.367101732e-30 pub = -3.205080160e-36
+ uc = 2.781855432e-11 luc = 1.116979589e-17 wuc = -7.614879963e-26 puc = 7.248449291e-32
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.284586148e+05 lvsat = 2.016794202e-01 wvsat = 1.014395847e-01 pvsat = -9.655841331e-8
+ a0 = 1.033165529e+00 la0 = 1.588065634e-07 wa0 = 3.682956162e-15 pa0 = -3.505736146e-21
+ ags = 2.238489660e+00 lags = -9.409245264e-07 wags = 1.627397239e-14 pags = -1.549089035e-20
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 5.649984843e-07 lb0 = -2.553120791e-13 wb0 = 1.227103407e-21 pb0 = -1.168056740e-27
+ b1 = 1.381407792e-08 lb1 = -6.242319397e-15 wb1 = -6.041060156e-23 pb1 = 5.750371683e-29
+ keta = -1.128952687e-01 lketa = 4.780085636e-08 wketa = 5.615223841e-16 pketa = -5.345026644e-22
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.248591517e+00 lpclm = -3.600504323e-07 wpclm = -4.301984546e-15 ppclm = 4.094976802e-21
+ pdiblc1 = 6.447801371e-01 lpdiblc1 = -2.764374528e-07 wpdiblc1 = 8.063683055e-16 ppdiblc1 = -7.675673430e-22
+ pdiblc2 = 8.895504672e-03 lpdiblc2 = -3.998725264e-09 wpdiblc2 = -1.943281647e-17 ppdiblc2 = 1.849771725e-23
+ pdiblcb = 8.513601967e-02 lpdiblcb = -8.122164648e-08 wpdiblcb = 1.561279621e-16 ppdiblcb = -1.486152911e-22
+ drout = 8.471347039e-01 ldrout = 6.907687722e-08 wdrout = -5.419309446e-16 pdrout = 5.158540262e-22
+ pscbe1 = 1.002269392e+09 lpscbe1 = -2.554584381e+02 wpscbe1 = 6.240154266e-06 ppscbe1 = -5.939882278e-12
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 6.984094428e-06 lalpha0 = -1.393643668e-12 walpha0 = 7.324625932e-21 palpha0 = -6.972178911e-27
+ alpha1 = 0.85
+ beta0 = 1.696331591e+01 lbeta0 = 4.765916758e-07 wbeta0 = -3.261334314e-14 pbeta0 = 3.104401003e-20
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.707775675e-01 lkt1 = -3.692777148e-09 wkt1 = 5.233502520e-17 pkt1 = -4.981792756e-23
+ kt2 = -1.845629470e-02 lkt2 = -8.252388772e-09 wkt2 = 8.530176565e-18 pkt2 = -8.119727113e-24
+ at = 1.097132692e+05 lat = -4.476243172e-02 wat = 6.481269374e-10 pat = -6.169396220e-16
+ ute = -8.616208302e-01 lute = -2.027400583e-07 wute = -1.339671485e-15 pute = 1.275207495e-21
+ ua1 = 1.688160724e-09 lua1 = -3.870320767e-16 wua1 = 2.775349774e-24 pua1 = -2.641806427e-30
+ ub1 = -7.051401795e-19 lub1 = 3.310533556e-26 wub1 = 6.089081742e-34 pub1 = -5.796078464e-40
+ uc1 = 7.289584960e-11 luc1 = -3.034625908e-17 wuc1 = -6.743962175e-26 puc1 = 6.419459221e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.123 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {8.718873043e-02+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 7.716644221e-08 wvth0 = 3.027724002e-07 pvth0 = -6.112399493e-14
+ k1 = 1.260614555e-01 lk1 = 1.576714905e-07 wk1 = 1.001961181e-15 pk1 = -2.022777501e-22
+ k2 = -1.165016602e-01 lk2 = -3.779077027e-09 wk2 = 1.249078059e-07 pk2 = -2.521651277e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.905328522e-01 ldsub = 5.412372030e-08 wdsub = 2.955236056e-16 pdsub = -5.966116490e-23
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.103590353e-03 lcdscd = -1.221701112e-9
+ cit = 0.0
+ voff = {-1.154994130e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.271458387e-08 wvoff = 1.219161661e-15 pvoff = -2.461255644e-22
+ nfactor = 3.206634057e+00 lnfactor = -8.661382449e-08 wnfactor = 1.184564269e-14 pnfactor = -2.391409737e-21
+ eta0 = 8.851262264e-01 leta0 = -1.785500340e-07 weta0 = -6.761524673e-16 peta0 = 1.365019209e-22
+ etab = 3.439973868e-02 letab = -1.582701388e-08 wetab = -1.358529678e-16 petab = 2.742613341e-23
+ u0 = 1.066248139e-01 lu0 = -1.554752483e-08 wu0 = -5.360160640e-08 pu0 = 1.082114590e-14
+ ua = -1.664072330e-09 lua = 9.725664221e-17 wua = 4.258378733e-24 pua = -8.596855019e-31
+ ub = 2.065358409e-18 lub = 3.728370425e-26 wub = -6.734203463e-30 pub = 1.359507726e-36
+ uc = 2.021746668e-11 luc = 1.460458297e-17 wuc = 1.522973925e-25 puc = -3.074594148e-32
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.611097133e+05 lvsat = -6.473530545e-02 wvsat = -2.028791694e-01 pvsat = 4.095744959e-8
+ a0 = 1.291411743e+00 la0 = 4.211000583e-08 wa0 = -7.365905219e-15 pa0 = 1.487036272e-21
+ ags = -7.269793207e-01 lags = 3.991145622e-07 wags = -3.254795722e-14 pags = 6.570814559e-21
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.086040475e-15 lb0 = -8.248939372e-22 wb0 = -2.454206663e-21 pb0 = 4.954576953e-28
+ b1 = -2.011568142e-16 lb1 = 4.060973881e-23 wb1 = 1.208212196e-22 pb1 = -2.439150864e-29
+ keta = 5.428652327e-02 lketa = -2.774541899e-08 wketa = -1.123044990e-15 pketa = 2.267214125e-22
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.240064034e-01 lpclm = -7.781228654e-08 wpclm = 8.603970869e-15 ppclm = -1.736978117e-21
+ pdiblc1 = -2.285578172e-01 lpdiblc1 = 1.182073753e-07 wpdiblc1 = -1.612737721e-15 ppdiblc1 = 3.255810899e-22
+ pdiblc2 = -6.704200135e-03 lpdiblc2 = 3.050484944e-09 wpdiblc2 = 3.886562014e-17 ppdiblc2 = -7.846230501e-24
+ pdiblcb = -8.758737370e-02 lpdiblcb = -3.171226754e-09 wpdiblcb = -3.122559988e-16 ppdiblcb = 6.303857436e-23
+ drout = 1.401075460e+00 ldrout = -1.812384256e-07 wdrout = 1.083861889e-15 pdrout = -2.188116355e-22
+ pscbe1 = 1.507016809e+08 lpscbe1 = 1.293488307e+02 wpscbe1 = -1.248030281e-05 ppscbe1 = 2.519536018e-12
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.031901106e-06 lalpha0 = -1.415246597e-12 walpha0 = -1.464927897e-20 palpha0 = 2.957412147e-27
+ alpha1 = 0.85
+ beta0 = 2.100422364e+01 lbeta0 = -1.349417753e-06 wbeta0 = 6.522657259e-14 pbeta0 = -1.316800535e-20
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.096264798e-01 lkt1 = 1.386230822e-08 wkt1 = -1.046736031e-16 pkt1 = 2.113131892e-23
+ kt2 = -4.304931438e-02 lkt2 = 2.860729551e-09 wkt2 = -1.706057517e-17 pkt2 = 3.444189378e-24
+ at = -3.932842210e+03 lat = 6.592086754e-03 wat = -1.296253758e-09 pat = 2.616889979e-16
+ ute = -1.303201522e+00 lute = -3.198133816e-09 wute = 2.679350075e-15 pute = -5.409095394e-22
+ ua1 = 1.522520014e-09 lua1 = -3.121821870e-16 wua1 = -5.550709474e-24 pua1 = 1.120583230e-30
+ ub1 = -1.713664126e-18 lub1 = 4.888381450e-25 wub1 = -1.217813267e-33 pub1 = 2.458549722e-40
+ uc1 = -1.084804680e-10 luc1 = 5.161425270e-17 wuc1 = 1.348793211e-25 puc1 = -2.722957731e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.124 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {6.130803429e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.900108240e-8
+ k1 = 9.070734896e-01 lk1 = 5.143085957e-17
+ k2 = -1.611477193e-01 lk2 = 5.234114019e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -7.794653811e-18
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999996e-03 lcdscd = 5.442070405e-19
+ cit = 0.0
+ voff = {-1.237493848e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.104907131e-8
+ nfactor = 2.484263783e+00 lnfactor = 5.921900879e-8
+ eta0 = 2.001909455e-03 leta0 = -2.640137943e-10
+ etab = -4.399800002e-02 letab = 2.220557072e-18
+ u0 = 2.919169366e-02 lu0 = 8.475092343e-11
+ ua = -1.224106221e-09 lua = 8.435844238e-18
+ ub = 2.103521860e-18 lub = 2.957922859e-26
+ uc = 1.218677263e-10 luc = -5.916673095e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.325369855e+05 lvsat = 1.597285411e-3
+ a0 = 1.499999999e+00 la0 = 1.571045516e-16
+ ags = 1.250000000e+00 lags = 3.363709311e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -6.898412508e-08 lb0 = 1.392658415e-14
+ b1 = 9.858632274e-11 lb1 = -1.990270542e-17
+ keta = -1.889316341e-01 lketa = 2.135570583e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.499568007e-01 lpclm = -2.248687870e-8
+ pdiblc1 = 3.569721502e-01 lpdiblc1 = -2.689670708e-17
+ pdiblc2 = 8.406112095e-03 lpdiblc2 = 7.211453656e-19
+ pdiblcb = -1.032957700e-01 lpdiblcb = 2.135402966e-18
+ drout = 5.033266589e-01 ldrout = 1.424531604e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 1.407623291e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 5.774280622e-09 lalpha0 = 3.194912098e-15
+ alpha1 = 0.85
+ beta0 = 1.518074234e+01 lbeta0 = -1.737675240e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.585636645e-01 lkt1 = 3.553695993e-9
+ kt2 = -2.887893901e-02 lkt2 = 8.536504836e-19
+ at = -1.837987011e+04 lat = 9.508667194e-3
+ ute = -1.325229293e+00 lute = 1.248854588e-9
+ ua1 = -2.384733722e-11 lua1 = 1.610623533e-25
+ ub1 = 7.077531683e-19 lub1 = 2.287958552e-34
+ uc1 = 1.471862500e-10 luc1 = -3.312858353e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.125 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {-6.442655289e-02+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.034920452e-08 wvth0 = 4.929305303e-07 pvth0 = -6.500817126e-14
+ k1 = 0.90707349
+ k2 = -4.372192880e-01 lk2 = 4.164270857e-08 wk2 = 1.511822721e-07 pk2 = -1.993806923e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.585234882e-01 ldsub = 1.404687923e-11 wdsub = 7.031613209e-11 pdsub = -9.273361816e-18
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000001e-03 lcdscd = -9.108686028e-20
+ cit = 0.0
+ voff = {-2.075300001e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.193267707e-17
+ nfactor = 6.715065073e+00 lnfactor = -4.987432961e-07 wnfactor = -2.551780856e-06 pnfactor = 3.365314110e-13
+ eta0 = 1.494623677e-02 leta0 = -1.971124625e-09 weta0 = -9.873962680e-09 peta0 = 1.302188072e-15
+ etab = -0.043998
+ u0 = 1.372433864e-01 lu0 = -1.416521437e-08 wu0 = -6.100665572e-08 pu0 = 8.045618763e-15
+ ua = 1.137845817e-09 lua = -3.030607526e-16 wua = -1.517341907e-15 pua = 2.001085681e-22
+ ub = -2.380181685e-18 lub = 6.208945359e-25 wub = 3.085345045e-24 pub = -4.068983898e-31
+ uc = 3.033951073e-10 luc = -2.985668563e-17 wuc = -1.494573658e-16 puc = 1.971058685e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.330544178e+05 lvsat = -2.484715409e-02 wvsat = -9.762143231e-02 pvsat = 1.287441211e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.002434794e-05 lb0 = -1.317192142e-12 wb0 = -6.516068161e-12 pb0 = 8.593455852e-19
+ b1 = 3.616569266e-07 lb1 = -4.770257818e-14 wb1 = -2.390742016e-13 pb1 = 3.152934478e-20
+ keta = -2.700000006e-02 lketa = 6.282308007e-18
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.545414303e-01 lpclm = 5.723495250e-08 wpclm = 2.788054324e-07 ppclm = -3.676913923e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.000000001e-08 lalpha0 = -1.379922550e-24
+ alpha1 = 0.85
+ beta0 = 1.390773688e+01 lbeta0 = -5.882290701e-9
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.491681677e-01 lkt1 = 2.869080848e-08 wkt1 = 1.422476686e-07 pkt1 = -1.875976478e-14
+ kt2 = -0.028878939
+ at = 5.372048693e+04 lat = 6.915419362e-12
+ ute = 7.529872056e-02 lute = -1.834541803e-07 wute = -9.109782294e-07 pute = 1.201407199e-13
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.126 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {0.4913699+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56800772
+ k2 = -0.040590746
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 2.78042
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.025731
+ ua = -1.0529435e-9
+ ub = 1.832e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 9.1484e-8
+ b1 = 1.6098e-9
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.127 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.753697877e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.192323364e-7
+ k1 = 6.121972372e-01 lk1 = -8.816639883e-7
+ k2 = -5.732582613e-02 lk2 = 3.338963274e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.017062664e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.311152548e-7
+ nfactor = 2.999527454e+00 lnfactor = -4.371605856e-06 wnfactor = 7.105427358e-21
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.399768874e-02 lu0 = 3.458282001e-8
+ ua = -1.240665649e-09 lua = 3.745409973e-15
+ ub = 1.951616170e-18 lub = -2.386567588e-24
+ uc = 6.326057033e-11 luc = -2.937629231e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.390829178e+00 la0 = -5.632251912e-7
+ ags = 3.209382116e-01 lags = 4.776837126e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 8.925150941e-08 lb0 = 4.454238660e-14 wb0 = -2.117582368e-28
+ b1 = 2.167571440e-09 lb1 = -1.112858939e-14
+ keta = -2.666112675e-03 lketa = -3.751925933e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.631270000e-03 lpclm = 5.288499448e-07 ppclm = -4.440892099e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 5.528995573e-04 lpdiblc2 = 8.128953030e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -7.319501400e+07 lpscbe1 = 5.949551434e+03 ppscbe1 = 3.814697266e-18
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.832257539e-01 lkt1 = -6.293314343e-8
+ kt2 = -3.544646383e-02 lkt2 = 1.182853816e-7
+ at = 1.981929863e+05 lat = -4.627437017e-01 wat = -4.656612873e-16
+ ute = -1.016200285e+00 lute = -1.979220918e-6
+ ua1 = 1.030149760e-09 lua1 = 1.812633186e-15
+ ub1 = -3.832369470e-19 lub1 = -3.715699712e-24
+ uc1 = 6.920223587e-11 luc1 = -7.059748407e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.128 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.174342346e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.525913972e-8
+ k1 = 4.373408531e-01 lk1 = 5.087731700e-7
+ k2 = 8.934565372e-03 lk2 = -1.929984209e-07 pk2 = -2.220446049e-28
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.179994591e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.553724997e-9
+ nfactor = 1.644821634e+00 lnfactor = 6.400853618e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.718425420e-02 lu0 = 9.243630640e-9
+ ua = -9.777670666e-10 lua = 1.654871732e-15
+ ub = 1.840111304e-18 lub = -1.499894165e-24
+ uc = 9.701328365e-12 luc = 1.321337955e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.408917323e+00 la0 = -7.070599674e-7
+ ags = 3.610925198e-01 lags = 1.583814327e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 5.011079129e-08 lb0 = 3.557847194e-13
+ b1 = -1.658197099e-09 lb1 = 1.929346677e-14
+ keta = -1.740241834e-02 lketa = 7.966208966e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -6.899761706e-01 lpclm = 5.938871634e-06 wpclm = 2.220446049e-22 ppclm = 3.552713679e-27
+ pdiblc1 = 0.39
+ pdiblc2 = -1.623723774e-03 lpdiblc2 = 2.543720274e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.392309919e+08 lpscbe1 = 2.844246136e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.862989458e-01 lkt1 = -3.849548711e-8
+ kt2 = -9.860889619e-03 lkt2 = -8.516805990e-8
+ at = 140000.0
+ ute = -1.231212620e+00 lute = -2.694684098e-7
+ ua1 = 1.514330084e-09 lua1 = -2.037511139e-15
+ ub1 = -1.026378584e-18 lub1 = 1.398486053e-24
+ uc1 = -7.088796187e-11 luc1 = 4.080057410e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.129 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.258444758e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.849541224e-8
+ k1 = 5.592357205e-01 lk1 = 2.705915957e-8
+ k2 = -3.344055097e-02 lk2 = -2.553700375e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.527821500e-01 ldsub = -1.157040216e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.370079140e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 7.356542684e-8
+ nfactor = 3.198174774e+00 lnfactor = 2.621868556e-7
+ eta0 = 1.575872698e-01 leta0 = -3.066156572e-7
+ etab = -1.378278648e-01 letab = 2.680476500e-7
+ u0 = 2.961611194e-02 lu0 = -3.667817484e-10
+ ua = -7.010393526e-10 lua = 5.612767375e-16
+ ub = 1.754049020e-18 lub = -1.159786258e-24
+ uc = 3.566812735e-11 luc = 2.951609590e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.605932281e+00 la0 = -1.485639637e-06 wa0 = -3.552713679e-21
+ ags = 3.277011992e-01 lags = 2.903399581e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 7.970976424e-08 lb0 = 2.388131005e-13
+ b1 = 8.033723719e-10 lb1 = 9.565637143e-15
+ keta = 5.453875497e-04 lketa = 8.734496589e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.112609403e+00 lpclm = -1.184732045e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.502894210e-03 lpdiblc2 = 9.129299537e-9
+ pdiblcb = -3.719925625e-02 lpdiblcb = 4.821000899e-8
+ drout = 0.56
+ pscbe1 = 6.245423126e+08 lpscbe1 = 3.424725263e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.591689679e-01 lkt1 = -1.457099312e-7
+ kt2 = -1.496516276e-02 lkt2 = -6.499657985e-8
+ at = 1.698930575e+05 lat = -1.181338060e-1
+ ute = -8.787696445e-01 lute = -1.662281110e-6
+ ua1 = 2.126322375e-09 lua1 = -4.456031847e-15
+ ub1 = -1.476118686e-18 lub1 = 3.175805416e-24
+ uc1 = 8.711055893e-12 luc1 = 9.343989506e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.130 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.784394203e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.403361498e-8
+ k1 = 5.910989287e-01 lk1 = -3.513403122e-8
+ k2 = -5.807107652e-02 lk2 = 2.253885108e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.26
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-6.567142512e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -6.567491050e-8
+ nfactor = 3.233958994e+00 lnfactor = 1.923403166e-7
+ eta0 = -1.433508281e-03 leta0 = 3.773978078e-09 weta0 = -1.734723476e-24 peta0 = -1.734723476e-30
+ etab = 7.933901888e-02 letab = -1.558362640e-07 wetab = -2.949029909e-23 petab = 3.642919300e-29
+ u0 = 3.161666009e-02 lu0 = -4.271613666e-9
+ ua = 2.752158536e-10 lua = -1.344257251e-15
+ ub = 3.376251922e-19 lub = 1.604904499e-24
+ uc = 6.148628680e-11 luc = -2.087787897e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.674837450e+04 lvsat = 6.346786025e-3
+ a0 = 5.066918688e-01 la0 = 6.599468372e-7
+ ags = -2.598775476e-01 lags = 1.437223750e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.118978317e-07 lb0 = 1.759858233e-13
+ b1 = 4.226685500e-09 lb1 = 2.883737292e-15
+ keta = 6.946103312e-02 lketa = -1.257806426e-07 wketa = -1.387778781e-23 pketa = -9.714451465e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.584889993e-01 lpclm = 6.775974424e-7
+ pdiblc1 = 4.239170811e-01 lpdiblc1 = -6.620210620e-8
+ pdiblc2 = 9.545914571e-03 lpdiblc2 = -4.617838089e-9
+ pdiblcb = -2.421622557e-02 lpdiblcb = 2.286867807e-8
+ drout = 2.176050537e-01 ldrout = 6.683141902e-7
+ pscbe1 = 8.629220470e+08 lpscbe1 = -1.228163479e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.195826690e-06 lalpha0 = 1.020019183e-11 walpha0 = -1.058791184e-27 palpha0 = 4.446922973e-33
+ alpha1 = 0.85
+ beta0 = 1.042942088e+01 lbeta0 = 6.696082211e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.901361166e-01 lkt1 = 1.099223579e-7
+ kt2 = -6.838621167e-02 lkt2 = 3.927495052e-8
+ at = 1.538056803e+05 lat = -8.673316007e-2
+ ute = -2.354634327e+00 lute = 1.218431122e-6
+ ua1 = -1.525599643e-09 lua1 = 2.672085355e-15 wua1 = 4.135903063e-31 pua1 = 1.654361225e-36
+ ub1 = 9.327016030e-19 lub1 = -1.525925138e-24 wub1 = -3.851859889e-40 pub1 = 3.851859889e-46
+ uc1 = 7.140092441e-11 luc1 = -2.892326820e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.131 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.137264256e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.044458513e-8
+ k1 = 6.257710813e-01 lk1 = -6.813779451e-8
+ k2 = -5.660819148e-02 lk2 = 2.114635860e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.145343276e-01 ldsub = 4.327790973e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.265594374e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.716768506e-9
+ nfactor = 3.816562506e+00 lnfactor = -3.622288970e-7
+ eta0 = -4.380244824e-01 leta0 = 4.193566311e-07 weta0 = 3.469446952e-23 peta0 = -2.775557562e-29
+ etab = -1.600650675e-01 letab = 7.204793714e-8
+ u0 = 3.099996783e-02 lu0 = -3.684596026e-9
+ ua = -8.551569684e-10 lua = -2.682768385e-16
+ ub = 1.911412760e-18 lub = 1.068460154e-25
+ uc = 2.781855419e-11 luc = 1.116979601e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.042946423e+04 lvsat = 4.091806665e-2
+ a0 = 1.033165535e+00 la0 = 1.588065576e-7
+ ags = 2.238489687e+00 lags = -9.409245522e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 5.649984864e-07 lb0 = -2.553120810e-13
+ b1 = 1.381407782e-08 lb1 = -6.242319301e-15
+ keta = -1.128952678e-01 lketa = 4.780085547e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.248591510e+00 lpclm = -3.600504255e-7
+ pdiblc1 = 6.447801385e-01 lpdiblc1 = -2.764374541e-7
+ pdiblc2 = 8.895504640e-03 lpdiblc2 = -3.998725233e-9
+ pdiblcb = 8.513601993e-02 lpdiblcb = -8.122164672e-08 wpdiblcb = -3.989863995e-23 ppdiblcb = -1.084202172e-29
+ drout = 8.471347030e-01 ldrout = 6.907687808e-8
+ pscbe1 = 1.002269402e+09 lpscbe1 = -2.554584480e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 6.984094440e-06 lalpha0 = -1.393643680e-12
+ alpha1 = 0.85
+ beta0 = 1.696331585e+01 lbeta0 = 4.765917275e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.707775674e-01 lkt1 = -3.692777231e-9
+ kt2 = -1.845629469e-02 lkt2 = -8.252388786e-9
+ at = 1.097132703e+05 lat = -4.476243274e-2
+ ute = -8.616208325e-01 lute = -2.027400562e-7
+ ua1 = 1.688160728e-09 lua1 = -3.870320811e-16
+ ub1 = -7.051401785e-19 lub1 = 3.310533460e-26
+ uc1 = 7.289584949e-11 luc1 = -3.034625897e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.132 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.912784230e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.459968901e-8
+ k1 = 1.260614572e-01 lk1 = 1.576714902e-7
+ k2 = 9.145896450e-02 lk2 = -4.576237591e-08 wk2 = -5.551115123e-23 pk2 = 4.163336342e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.905328527e-01 ldsub = 5.412372020e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.103590353e-03 lcdscd = -1.221701112e-9
+ cit = 0.0
+ voff = {-1.154994110e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.271458428e-8
+ nfactor = 3.206634077e+00 lnfactor = -8.661382847e-8
+ eta0 = 8.851262252e-01 leta0 = -1.785500338e-7
+ etab = 3.439973846e-02 letab = -1.582701384e-08 wetab = -1.040834086e-23 petab = -8.239936511e-30
+ u0 = 1.738280483e-02 lu0 = 2.468741208e-9
+ ua = -1.664072323e-09 lua = 9.725664078e-17
+ ub = 2.065347197e-18 lub = 3.728596771e-26
+ uc = 2.021746693e-11 luc = 1.460458292e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.233335552e+05 lvsat = 3.455283115e-3
+ a0 = 1.291411731e+00 la0 = 4.211000830e-8
+ ags = -7.269793749e-01 lags = 3.991145732e-07 wags = -4.440892099e-22 pags = 3.330669074e-28
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 5.428652140e-02 lketa = -2.774541861e-08 pketa = -2.081668171e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.240064177e-01 lpclm = -7.781228943e-8
+ pdiblc1 = -2.285578199e-01 lpdiblc1 = 1.182073759e-07 wpdiblc1 = -2.220446049e-22
+ pdiblc2 = -6.704200070e-03 lpdiblc2 = 3.050484931e-09 wpdiblc2 = 4.011548038e-24 ppdiblc2 = 2.493664997e-30
+ pdiblcb = -8.758737422e-02 lpdiblcb = -3.171226649e-9
+ drout = 1.401075462e+00 ldrout = -1.812384259e-7
+ pscbe1 = 1.507016602e+08 lpscbe1 = 1.293488349e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.031901081e-06 lalpha0 = -1.415246593e-12
+ alpha1 = 0.85
+ beta0 = 2.100422375e+01 lbeta0 = -1.349417775e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.096264800e-01 lkt1 = 1.386230826e-8
+ kt2 = -4.304931441e-02 lkt2 = 2.860729557e-9
+ at = -3.932844369e+03 lat = 6.592087190e-3
+ ute = -1.303201517e+00 lute = -3.198134717e-9
+ ua1 = 1.522520004e-09 lua1 = -3.121821851e-16
+ ub1 = -1.713664128e-18 lub1 = 4.888381454e-25 wub1 = -1.540743956e-39
+ uc1 = -1.084804678e-10 luc1 = 5.161425266e-17 wuc1 = 2.584939414e-32 puc1 = -2.261821987e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.133 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {6.130803429e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.900108240e-8
+ k1 = 9.070734896e-01 lk1 = 5.142908321e-17
+ k2 = -1.611477193e-01 lk2 = 5.234114019e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -7.794653811e-18
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999996e-03 lcdscd = 5.442105100e-19
+ cit = 0.0
+ voff = {-1.237493848e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.104907131e-8
+ nfactor = 2.484263783e+00 lnfactor = 5.921900879e-8
+ eta0 = 2.001909455e-03 leta0 = -2.640137943e-10
+ etab = -4.399800002e-02 letab = 2.220557072e-18
+ u0 = 2.919169366e-02 lu0 = 8.475092343e-11
+ ua = -1.224106221e-09 lua = 8.435844238e-18
+ ub = 2.103521860e-18 lub = 2.957922859e-26
+ uc = 1.218677263e-10 luc = -5.916673095e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.325369855e+05 lvsat = 1.597285411e-3
+ a0 = 1.499999999e+00 la0 = 1.571063279e-16
+ ags = 1.250000000e+00 lags = 3.363709311e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -6.898412508e-08 lb0 = 1.392658415e-14
+ b1 = 9.858632274e-11 lb1 = -1.990270542e-17
+ keta = -1.889316341e-01 lketa = 2.135570583e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.499568007e-01 lpclm = -2.248687870e-8
+ pdiblc1 = 3.569721502e-01 lpdiblc1 = -2.689626299e-17
+ pdiblc2 = 8.406112095e-03 lpdiblc2 = 7.211592434e-19
+ pdiblcb = -1.032957700e-01 lpdiblcb = 2.135291943e-18
+ drout = 5.033266589e-01 ldrout = 1.424531604e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 1.407337189e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 5.774280622e-09 lalpha0 = 3.194912098e-15
+ alpha1 = 0.85
+ beta0 = 1.518074234e+01 lbeta0 = -1.737675240e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.585636645e-01 lkt1 = 3.553695993e-9
+ kt2 = -2.887893901e-02 lkt2 = 8.535949725e-19
+ at = -1.837987011e+04 lat = 9.508667194e-3
+ ute = -1.325229293e+00 lute = 1.248854588e-9
+ ua1 = -2.384733722e-11 lua1 = 1.610623533e-25
+ ub1 = 7.077531683e-19 lub1 = 2.287966255e-34
+ uc1 = 1.471862500e-10 luc1 = -3.312858353e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.134 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {2.343188208e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.571694377e-07 wvth0 = -9.531599387e-07 pvth0 = 1.257036859e-13
+ k1 = 0.90707349
+ k2 = 1.002030108e-02 lk2 = -1.733969567e-08 wk2 = -1.174441367e-07 pk2 = 1.548865020e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.585222866e-01 ldsub = 1.420534621e-11 wdsub = 7.103784591e-11 pdsub = -9.368542157e-18
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000001e-03 lcdscd = -9.108339083e-20
+ cit = 0.0
+ voff = {-2.075300001e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.193267707e-17
+ nfactor = 6.715065176e+00 lnfactor = -4.987433096e-07 wnfactor = -2.551780918e-06 pnfactor = 3.365314192e-13
+ eta0 = 1.494620783e-02 leta0 = -1.971120808e-09 weta0 = -9.873945296e-09 peta0 = 1.302185780e-15
+ etab = -0.043998
+ u0 = -2.506096201e-01 lu0 = 3.698522798e-08 wu0 = 1.719502713e-07 pu0 = -2.267697372e-14
+ ua = 1.137843041e-09 lua = -3.030603864e-16 wua = -1.517340239e-15 pua = 2.001083481e-22
+ ub = -2.380190426e-18 lub = 6.208956887e-25 wub = 3.085350295e-24 pub = -4.068990822e-31
+ uc = 3.059431155e-10 luc = -3.019271950e-17 wuc = -1.509877810e-16 puc = 1.991241955e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.172609747e+05 lvsat = -9.576199013e-03 wvsat = -2.807218497e-02 pvsat = 3.702187826e-9
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.002439566e-05 lb0 = -1.317198436e-12 wb0 = -6.516096826e-12 pb0 = 8.593493655e-19
+ b1 = 3.616608296e-07 lb1 = -4.770309291e-14 wb1 = -2.390765458e-13 pb1 = 3.152965394e-20
+ keta = -2.700000006e-02 lketa = 6.282363518e-18
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.545414373e-01 lpclm = 5.723495342e-08 wpclm = 2.788054366e-07 ppclm = -3.676913979e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.000000001e-08 lalpha0 = -1.379922550e-24
+ alpha1 = 0.85
+ beta0 = 1.390773688e+01 lbeta0 = -5.882290701e-9
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.491681764e-01 lkt1 = 2.869080963e-08 wkt1 = 1.422476738e-07 pkt1 = -1.875976547e-14
+ kt2 = -0.028878939
+ at = 5.372048693e+04 lat = 6.915302947e-12
+ ute = 9.082946736e-02 lute = -1.855023908e-07 wute = -9.203064929e-07 pute = 1.213709406e-13
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.135 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {0.4913699+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56800772
+ k2 = -0.040590746
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 2.78042
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.025731
+ ua = -1.0529435e-9
+ ub = 1.832e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 9.1484e-8
+ b1 = 1.6098e-9
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.136 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.753697877e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.192323364e-7
+ k1 = 6.121972372e-01 lk1 = -8.816639883e-7
+ k2 = -5.732582613e-02 lk2 = 3.338963274e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.017062664e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.311152548e-7
+ nfactor = 2.999527454e+00 lnfactor = -4.371605856e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.399768874e-02 lu0 = 3.458282001e-8
+ ua = -1.240665649e-09 lua = 3.745409973e-15
+ ub = 1.951616170e-18 lub = -2.386567588e-24
+ uc = 6.326057033e-11 luc = -2.937629231e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.390829178e+00 la0 = -5.632251912e-7
+ ags = 3.209382116e-01 lags = 4.776837126e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 8.925150941e-08 lb0 = 4.454238660e-14
+ b1 = 2.167571440e-09 lb1 = -1.112858939e-14 wb1 = -1.323488980e-29
+ keta = -2.666112675e-03 lketa = -3.751925933e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.631270000e-03 lpclm = 5.288499448e-07 ppclm = 8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 5.528995573e-04 lpdiblc2 = 8.128953030e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -7.319501400e+07 lpscbe1 = 5.949551434e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.832257539e-01 lkt1 = -6.293314343e-08 wkt1 = -1.776356839e-21
+ kt2 = -3.544646383e-02 lkt2 = 1.182853816e-7
+ at = 1.981929863e+05 lat = -4.627437017e-1
+ ute = -1.016200285e+00 lute = -1.979220918e-06 wute = -7.105427358e-21
+ ua1 = 1.030149760e-09 lua1 = 1.812633186e-15
+ ub1 = -3.832369470e-19 lub1 = -3.715699712e-24
+ uc1 = 6.920223587e-11 luc1 = -7.059748407e-16 wuc1 = -2.067951531e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.137 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.174342346e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.525913972e-8
+ k1 = 4.373408531e-01 lk1 = 5.087731700e-7
+ k2 = 8.934565372e-03 lk2 = -1.929984209e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.179994591e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.553724997e-9
+ nfactor = 1.644821634e+00 lnfactor = 6.400853618e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.718425420e-02 lu0 = 9.243630640e-9
+ ua = -9.777670666e-10 lua = 1.654871732e-15
+ ub = 1.840111304e-18 lub = -1.499894165e-24
+ uc = 9.701328365e-12 luc = 1.321337955e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.408917323e+00 la0 = -7.070599674e-7
+ ags = 3.610925198e-01 lags = 1.583814327e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 5.011079129e-08 lb0 = 3.557847194e-13
+ b1 = -1.658197099e-09 lb1 = 1.929346677e-14 pb1 = 5.293955920e-35
+ keta = -1.740241834e-02 lketa = 7.966208966e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -6.899761706e-01 lpclm = 5.938871634e-06 wpclm = -4.440892099e-22 ppclm = -1.776356839e-27
+ pdiblc1 = 0.39
+ pdiblc2 = -1.623723774e-03 lpdiblc2 = 2.543720274e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.392309919e+08 lpscbe1 = 2.844246136e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.862989458e-01 lkt1 = -3.849548711e-8
+ kt2 = -9.860889619e-03 lkt2 = -8.516805990e-8
+ at = 140000.0
+ ute = -1.231212620e+00 lute = -2.694684098e-7
+ ua1 = 1.514330084e-09 lua1 = -2.037511139e-15
+ ub1 = -1.026378584e-18 lub1 = 1.398486053e-24
+ uc1 = -7.088796187e-11 luc1 = 4.080057410e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.138 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.258444758e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.849541224e-8
+ k1 = 5.592357205e-01 lk1 = 2.705915957e-8
+ k2 = -3.344055097e-02 lk2 = -2.553700375e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.527821500e-01 ldsub = -1.157040216e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.370079140e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 7.356542684e-8
+ nfactor = 3.198174774e+00 lnfactor = 2.621868556e-7
+ eta0 = 1.575872697e-01 leta0 = -3.066156572e-7
+ etab = -1.378278647e-01 letab = 2.680476500e-7
+ u0 = 2.961611194e-02 lu0 = -3.667817484e-10
+ ua = -7.010393526e-10 lua = 5.612767375e-16
+ ub = 1.754049020e-18 lub = -1.159786258e-24
+ uc = 3.566812735e-11 luc = 2.951609590e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.605932281e+00 la0 = -1.485639637e-6
+ ags = 3.277011992e-01 lags = 2.903399581e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 7.970976424e-08 lb0 = 2.388131005e-13
+ b1 = 8.033723719e-10 lb1 = 9.565637143e-15
+ keta = 5.453875497e-04 lketa = 8.734496589e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.112609403e+00 lpclm = -1.184732045e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.502894210e-03 lpdiblc2 = 9.129299537e-9
+ pdiblcb = -3.719925625e-02 lpdiblcb = 4.821000899e-8
+ drout = 0.56
+ pscbe1 = 6.245423126e+08 lpscbe1 = 3.424725263e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.591689679e-01 lkt1 = -1.457099312e-7
+ kt2 = -1.496516276e-02 lkt2 = -6.499657985e-8
+ at = 1.698930575e+05 lat = -1.181338060e-1
+ ute = -8.787696445e-01 lute = -1.662281110e-6
+ ua1 = 2.126322375e-09 lua1 = -4.456031847e-15
+ ub1 = -1.476118686e-18 lub1 = 3.175805416e-24
+ uc1 = 8.711055893e-12 luc1 = 9.343989506e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.139 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.784394203e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.403361498e-8
+ k1 = 5.910989287e-01 lk1 = -3.513403122e-8
+ k2 = -5.807107652e-02 lk2 = 2.253885108e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.26
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-6.567142512e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -6.567491050e-8
+ nfactor = 3.233958994e+00 lnfactor = 1.923403166e-7
+ eta0 = -1.433508281e-03 leta0 = 3.773978078e-09 weta0 = -3.469446952e-24
+ etab = 7.933901887e-02 letab = -1.558362640e-07 wetab = -2.428612866e-23 petab = -1.665334537e-28
+ u0 = 3.161666009e-02 lu0 = -4.271613666e-9
+ ua = 2.752158536e-10 lua = -1.344257251e-15
+ ub = 3.376251922e-19 lub = 1.604904499e-24
+ uc = 6.148628680e-11 luc = -2.087787897e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.674837450e+04 lvsat = 6.346786025e-3
+ a0 = 5.066918688e-01 la0 = 6.599468372e-7
+ ags = -2.598775476e-01 lags = 1.437223750e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.118978317e-07 lb0 = 1.759858233e-13
+ b1 = 4.226685500e-09 lb1 = 2.883737292e-15
+ keta = 6.946103312e-02 lketa = -1.257806426e-07 wketa = 1.110223025e-22
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.584889993e-01 lpclm = 6.775974424e-7
+ pdiblc1 = 4.239170811e-01 lpdiblc1 = -6.620210620e-8
+ pdiblc2 = 9.545914571e-03 lpdiblc2 = -4.617838089e-9
+ pdiblcb = -2.421622557e-02 lpdiblcb = 2.286867807e-8
+ drout = 2.176050537e-01 ldrout = 6.683141902e-7
+ pscbe1 = 8.629220470e+08 lpscbe1 = -1.228163479e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.195826690e-06 lalpha0 = 1.020019183e-11 walpha0 = -4.023406499e-27 palpha0 = 2.604626313e-32
+ alpha1 = 0.85
+ beta0 = 1.042942088e+01 lbeta0 = 6.696082211e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.901361166e-01 lkt1 = 1.099223579e-7
+ kt2 = -6.838621167e-02 lkt2 = 3.927495052e-8
+ at = 1.538056803e+05 lat = -8.673316007e-02 wat = 9.313225746e-16
+ ute = -2.354634327e+00 lute = 1.218431122e-6
+ ua1 = -1.525599643e-09 lua1 = 2.672085355e-15 pua1 = 6.617444900e-36
+ ub1 = 9.327016030e-19 lub1 = -1.525925138e-24
+ uc1 = 7.140092441e-11 luc1 = -2.892326820e-17 wuc1 = -4.135903063e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.140 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.137264256e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.044458513e-8
+ k1 = 6.257710813e-01 lk1 = -6.813779451e-8
+ k2 = -5.660819148e-02 lk2 = 2.114635860e-08 pk2 = 1.110223025e-28
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.145343276e-01 ldsub = 4.327790973e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.265594374e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.716768506e-9
+ nfactor = 3.816562506e+00 lnfactor = -3.622288970e-7
+ eta0 = -4.380244824e-01 leta0 = 4.193566311e-07 weta0 = -7.771561172e-22 peta0 = -4.857225733e-28
+ etab = -1.600650675e-01 letab = 7.204793714e-8
+ u0 = 3.099996783e-02 lu0 = -3.684596026e-9
+ ua = -8.551569684e-10 lua = -2.682768385e-16
+ ub = 1.911412760e-18 lub = 1.068460154e-25
+ uc = 2.781855419e-11 luc = 1.116979601e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.042946423e+04 lvsat = 4.091806665e-2
+ a0 = 1.033165535e+00 la0 = 1.588065576e-7
+ ags = 2.238489687e+00 lags = -9.409245522e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 5.649984864e-07 lb0 = -2.553120810e-13
+ b1 = 1.381407782e-08 lb1 = -6.242319301e-15
+ keta = -1.128952678e-01 lketa = 4.780085547e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.248591510e+00 lpclm = -3.600504255e-7
+ pdiblc1 = 6.447801385e-01 lpdiblc1 = -2.764374541e-7
+ pdiblc2 = 8.895504640e-03 lpdiblc2 = -3.998725233e-9
+ pdiblcb = 8.513601993e-02 lpdiblcb = -8.122164672e-08 wpdiblcb = -1.387778781e-22 ppdiblcb = -9.194034423e-29
+ drout = 8.471347030e-01 ldrout = 6.907687808e-8
+ pscbe1 = 1.002269402e+09 lpscbe1 = -2.554584480e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 6.984094440e-06 lalpha0 = -1.393643680e-12
+ alpha1 = 0.85
+ beta0 = 1.696331585e+01 lbeta0 = 4.765917275e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.707775674e-01 lkt1 = -3.692777231e-9
+ kt2 = -1.845629469e-02 lkt2 = -8.252388786e-9
+ at = 1.097132703e+05 lat = -4.476243274e-2
+ ute = -8.616208325e-01 lute = -2.027400562e-7
+ ua1 = 1.688160728e-09 lua1 = -3.870320811e-16
+ ub1 = -7.051401785e-19 lub1 = 3.310533460e-26
+ uc1 = 7.289584949e-11 luc1 = -3.034625897e-17 wuc1 = 4.135903063e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.141 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.912784230e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.459968901e-8
+ k1 = 1.260614572e-01 lk1 = 1.576714902e-7
+ k2 = 9.145896450e-02 lk2 = -4.576237591e-08 pk2 = -9.714451465e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.905328527e-01 ldsub = 5.412372020e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.103590353e-03 lcdscd = -1.221701112e-9
+ cit = 0.0
+ voff = {-1.154994110e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.271458428e-8
+ nfactor = 3.206634077e+00 lnfactor = -8.661382847e-8
+ eta0 = 8.851262252e-01 leta0 = -1.785500338e-7
+ etab = 3.439973846e-02 letab = -1.582701384e-08 wetab = -2.775557562e-23 petab = -1.387778781e-29
+ u0 = 1.738280483e-02 lu0 = 2.468741208e-9
+ ua = -1.664072323e-09 lua = 9.725664078e-17
+ ub = 2.065347197e-18 lub = 3.728596771e-26
+ uc = 2.021746693e-11 luc = 1.460458292e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.233335552e+05 lvsat = 3.455283115e-3
+ a0 = 1.291411731e+00 la0 = 4.211000830e-8
+ ags = -7.269793749e-01 lags = 3.991145732e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 5.428652140e-02 lketa = -2.774541861e-08 pketa = -1.387778781e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.240064177e-01 lpclm = -7.781228943e-8
+ pdiblc1 = -2.285578199e-01 lpdiblc1 = 1.182073759e-07 ppdiblc1 = 2.220446049e-28
+ pdiblc2 = -6.704200070e-03 lpdiblc2 = 3.050484931e-09 wpdiblc2 = 2.602085214e-24 ppdiblc2 = -6.505213035e-31
+ pdiblcb = -8.758737422e-02 lpdiblcb = -3.171226649e-9
+ drout = 1.401075462e+00 ldrout = -1.812384259e-7
+ pscbe1 = 1.507016602e+08 lpscbe1 = 1.293488349e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.031901081e-06 lalpha0 = -1.415246593e-12
+ alpha1 = 0.85
+ beta0 = 2.100422375e+01 lbeta0 = -1.349417775e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.096264800e-01 lkt1 = 1.386230826e-8
+ kt2 = -4.304931441e-02 lkt2 = 2.860729557e-9
+ at = -3.932844369e+03 lat = 6.592087190e-3
+ ute = -1.303201517e+00 lute = -3.198134717e-9
+ ua1 = 1.522520004e-09 lua1 = -3.121821851e-16
+ ub1 = -1.713664128e-18 lub1 = 4.888381454e-25 wub1 = 6.162975822e-39 pub1 = -1.540743956e-45
+ uc1 = -1.084804678e-10 luc1 = 5.161425266e-17 wuc1 = -5.169878828e-32 puc1 = -6.462348536e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.142 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {6.130803429e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.900108240e-8
+ k1 = 9.070734896e-01 lk1 = 5.142553050e-17
+ k2 = -1.611477193e-01 lk2 = 5.234114019e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -7.794653811e-18
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999996e-03 lcdscd = 5.442105100e-19
+ cit = 0.0
+ voff = {-1.237493848e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.104907131e-8
+ nfactor = 2.484263783e+00 lnfactor = 5.921900879e-8
+ eta0 = 2.001909455e-03 leta0 = -2.640137943e-10
+ etab = -4.399800002e-02 letab = 2.220446049e-18
+ u0 = 2.919169366e-02 lu0 = 8.475092343e-11
+ ua = -1.224106221e-09 lua = 8.435844238e-18
+ ub = 2.103521860e-18 lub = 2.957922859e-26
+ uc = 1.218677263e-10 luc = -5.916673095e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.325369855e+05 lvsat = 1.597285411e-3
+ a0 = 1.499999999e+00 la0 = 1.571081043e-16
+ ags = 1.250000000e+00 lags = 3.363354040e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -6.898412508e-08 lb0 = 1.392658415e-14
+ b1 = 9.858632274e-11 lb1 = -1.990270542e-17
+ keta = -1.889316341e-01 lketa = 2.135570583e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.499568007e-01 lpclm = -2.248687870e-8
+ pdiblc1 = 3.569721502e-01 lpdiblc1 = -2.689581891e-17
+ pdiblc2 = 8.406112095e-03 lpdiblc2 = 7.211453656e-19
+ pdiblcb = -1.032957700e-01 lpdiblcb = 2.135180921e-18
+ drout = 5.033266589e-01 ldrout = 1.424531604e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 1.407432556e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 5.774280622e-09 lalpha0 = 3.194912098e-15
+ alpha1 = 0.85
+ beta0 = 1.518074234e+01 lbeta0 = -1.737675240e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.585636645e-01 lkt1 = 3.553695993e-9
+ kt2 = -2.887893901e-02 lkt2 = 8.536504836e-19
+ at = -1.837987011e+04 lat = 9.508667194e-3
+ ute = -1.325229293e+00 lute = 1.248854588e-9
+ ua1 = -2.384733722e-11 lua1 = 1.610623016e-25
+ ub1 = 7.077531683e-19 lub1 = 2.287973959e-34
+ uc1 = 1.471862500e-10 luc1 = -3.312858353e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.143 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {-6.272620538e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.790920355e-07 wvth0 = 3.963296238e-06 pvth0 = -5.226834711e-13
+ k1 = 0.90707349
+ k2 = -8.057537200e-01 lk2 = 9.024539800e-08 wk2 = 3.480626245e-07 pk2 = -4.590284698e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.292022457e+00 ldsub = -2.417896307e-07 wdsub = -1.046182832e-06 pdsub = 1.379716380e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000001e-03 lcdscd = -9.109379917e-20
+ cit = 0.0
+ voff = {-2.075300001e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.193178889e-17
+ nfactor = -6.851256624e-01 lnfactor = 4.772012583e-07 wnfactor = 1.671004781e-06 pnfactor = -2.203737815e-13
+ eta0 = -1.034733598e-02 leta0 = 1.364617042e-09 weta0 = 4.559360192e-09 peta0 = -6.012929814e-16
+ etab = -0.043998
+ u0 = 8.925923967e-01 lu0 = -1.137813972e-07 wu0 = -4.803973820e-07 pu0 = 6.335528713e-14
+ ua = -2.896755218e-09 lua = 2.290264665e-16 wua = 7.849306339e-16 pua = -1.035174369e-22
+ ub = 1.246657437e-17 lub = -1.337110499e-24 wub = -5.386688792e-24 pub = 7.104019046e-31
+ uc = -1.724233205e-10 luc = 3.289472445e-17 wuc = 1.219834151e-16 puc = -1.608729477e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.531722760e+05 lvsat = -5.387651734e-02 wvsat = -2.197539227e-01 pvsat = 2.898136708e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -9.545585136e-06 lb0 = 1.263710202e-12 wb0 = 4.651160457e-12 pb0 = -6.133996923e-19
+ b1 = 1.210993705e-08 lb1 = -1.603971650e-15 wb1 = -3.961162091e-14 pb1 = 5.224020177e-21
+ keta = -7.798041805e-01 lketa = 9.928056812e-08 wketa = 4.295741551e-07 pketa = -5.665266915e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 8.437960589e-03 lpclm = 2.255296745e-08 wpclm = 1.287409769e-07 ppclm = -1.697848877e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.999997786e-08 lalpha0 = 2.920105005e-21 walpha0 = 1.264088677e-20 palpha0 = -1.667092819e-27
+ alpha1 = 0.85
+ beta0 = 1.390773666e+01 lbeta0 = -5.882262790e-09 wbeta0 = 1.207688456e-13 pbeta0 = -1.592709964e-20
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.998872423e-01 lkt1 = -4.184609246e-09 wkt1 = -4.218321692e-15 pkt1 = 5.563167704e-22
+ kt2 = -0.028878939
+ at = 5.372048932e+04 lat = -3.078503069e-10 wat = -1.361951232e-09 pat = 1.796154538e-16
+ ute = -1.122200093e+00 lute = -2.552683935e-08 wute = -2.281130090e-07 pute = 3.008377174e-14
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.144 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {0.4913699+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56800772
+ k2 = -0.040590746
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 2.78042
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.025731
+ ua = -1.0529435e-9
+ ub = 1.832e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 9.1484e-8
+ b1 = 1.6098e-9
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.145 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.753697877e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.192323364e-7
+ k1 = 6.121972372e-01 lk1 = -8.816639883e-7
+ k2 = -5.732582613e-02 lk2 = 3.338963274e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.017062664e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.311152548e-7
+ nfactor = 2.999527454e+00 lnfactor = -4.371605856e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.399768874e-02 lu0 = 3.458282001e-8
+ ua = -1.240665649e-09 lua = 3.745409973e-15
+ ub = 1.951616170e-18 lub = -2.386567588e-24
+ uc = 6.326057033e-11 luc = -2.937629231e-16 wuc = -2.067951531e-31
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.390829178e+00 la0 = -5.632251912e-7
+ ags = 3.209382116e-01 lags = 4.776837126e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 8.925150941e-08 lb0 = 4.454238660e-14
+ b1 = 2.167571440e-09 lb1 = -1.112858939e-14
+ keta = -2.666112675e-03 lketa = -3.751925933e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.631270000e-03 lpclm = 5.288499448e-07 ppclm = 8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 5.528995573e-04 lpdiblc2 = 8.128953030e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -7.319501400e+07 lpscbe1 = 5.949551434e+03 ppscbe1 = -7.629394531e-18
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.832257539e-01 lkt1 = -6.293314343e-8
+ kt2 = -3.544646383e-02 lkt2 = 1.182853816e-7
+ at = 1.981929863e+05 lat = -4.627437017e-1
+ ute = -1.016200285e+00 lute = -1.979220918e-6
+ ua1 = 1.030149760e-09 lua1 = 1.812633186e-15
+ ub1 = -3.832369470e-19 lub1 = -3.715699712e-24
+ uc1 = 6.920223587e-11 luc1 = -7.059748407e-16 puc1 = -8.271806126e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.146 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.174342346e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.525913972e-8
+ k1 = 4.373408531e-01 lk1 = 5.087731700e-7
+ k2 = 8.934565372e-03 lk2 = -1.929984209e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.179994591e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.553724997e-9
+ nfactor = 1.644821634e+00 lnfactor = 6.400853618e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.718425420e-02 lu0 = 9.243630640e-9
+ ua = -9.777670666e-10 lua = 1.654871732e-15
+ ub = 1.840111304e-18 lub = -1.499894165e-24
+ uc = 9.701328365e-12 luc = 1.321337955e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.408917323e+00 la0 = -7.070599674e-7
+ ags = 3.610925198e-01 lags = 1.583814327e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 5.011079129e-08 lb0 = 3.557847194e-13
+ b1 = -1.658197099e-09 lb1 = 1.929346677e-14
+ keta = -1.740241834e-02 lketa = 7.966208966e-08 wketa = 2.775557562e-23
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -6.899761706e-01 lpclm = 5.938871634e-06 wpclm = 2.220446049e-22 ppclm = 3.552713679e-27
+ pdiblc1 = 0.39
+ pdiblc2 = -1.623723774e-03 lpdiblc2 = 2.543720274e-08 ppdiblc2 = 2.775557562e-29
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.392309919e+08 lpscbe1 = 2.844246136e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.862989458e-01 lkt1 = -3.849548711e-8
+ kt2 = -9.860889619e-03 lkt2 = -8.516805990e-8
+ at = 140000.0
+ ute = -1.231212620e+00 lute = -2.694684098e-7
+ ua1 = 1.514330084e-09 lua1 = -2.037511139e-15
+ ub1 = -1.026378584e-18 lub1 = 1.398486053e-24
+ uc1 = -7.088796187e-11 luc1 = 4.080057410e-16 wuc1 = -1.033975766e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.147 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.258444758e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.849541224e-8
+ k1 = 5.592357205e-01 lk1 = 2.705915957e-8
+ k2 = -3.344055097e-02 lk2 = -2.553700375e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.527821500e-01 ldsub = -1.157040216e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.370079140e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 7.356542684e-08 wvoff = 4.440892099e-22
+ nfactor = 3.198174774e+00 lnfactor = 2.621868556e-7
+ eta0 = 1.575872698e-01 leta0 = -3.066156572e-7
+ etab = -1.378278647e-01 letab = 2.680476500e-7
+ u0 = 2.961611194e-02 lu0 = -3.667817484e-10
+ ua = -7.010393526e-10 lua = 5.612767375e-16
+ ub = 1.754049020e-18 lub = -1.159786258e-24
+ uc = 3.566812735e-11 luc = 2.951609590e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.605932281e+00 la0 = -1.485639637e-6
+ ags = 3.277011992e-01 lags = 2.903399581e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 7.970976424e-08 lb0 = 2.388131005e-13
+ b1 = 8.033723719e-10 lb1 = 9.565637143e-15
+ keta = 5.453875497e-04 lketa = 8.734496589e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.112609403e+00 lpclm = -1.184732045e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.502894210e-03 lpdiblc2 = 9.129299537e-9
+ pdiblcb = -3.719925625e-02 lpdiblcb = 4.821000899e-8
+ drout = 0.56
+ pscbe1 = 6.245423126e+08 lpscbe1 = 3.424725263e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.591689679e-01 lkt1 = -1.457099312e-7
+ kt2 = -1.496516276e-02 lkt2 = -6.499657985e-8
+ at = 1.698930575e+05 lat = -1.181338060e-1
+ ute = -8.787696445e-01 lute = -1.662281110e-6
+ ua1 = 2.126322375e-09 lua1 = -4.456031847e-15
+ ub1 = -1.476118686e-18 lub1 = 3.175805416e-24
+ uc1 = 8.711055893e-12 luc1 = 9.343989506e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.148 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.784394203e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.403361498e-8
+ k1 = 5.910989287e-01 lk1 = -3.513403122e-8
+ k2 = -5.807107652e-02 lk2 = 2.253885108e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.26
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-6.567142512e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -6.567491050e-8
+ nfactor = 3.233958994e+00 lnfactor = 1.923403166e-7
+ eta0 = -1.433508281e-03 leta0 = 3.773978078e-09 peta0 = 1.734723476e-30
+ etab = 7.933901888e-02 letab = -1.558362640e-07 wetab = -6.245004514e-23 petab = 2.133709875e-28
+ u0 = 3.161666009e-02 lu0 = -4.271613666e-9
+ ua = 2.752158536e-10 lua = -1.344257251e-15 pua = 1.654361225e-36
+ ub = 3.376251922e-19 lub = 1.604904499e-24
+ uc = 6.148628680e-11 luc = -2.087787897e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.674837450e+04 lvsat = 6.346786025e-3
+ a0 = 5.066918688e-01 la0 = 6.599468372e-7
+ ags = -2.598775475e-01 lags = 1.437223750e-06 pags = 1.776356839e-27
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.118978317e-07 lb0 = 1.759858233e-13
+ b1 = 4.226685500e-09 lb1 = 2.883737292e-15
+ keta = 6.946103312e-02 lketa = -1.257806426e-07 wketa = -8.326672685e-23 pketa = 5.551115123e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.584889993e-01 lpclm = 6.775974424e-7
+ pdiblc1 = 4.239170811e-01 lpdiblc1 = -6.620210620e-8
+ pdiblc2 = 9.545914571e-03 lpdiblc2 = -4.617838089e-9
+ pdiblcb = -2.421622557e-02 lpdiblcb = 2.286867807e-8
+ drout = 2.176050537e-01 ldrout = 6.683141902e-7
+ pscbe1 = 8.629220470e+08 lpscbe1 = -1.228163479e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.195826690e-06 lalpha0 = 1.020019183e-11 walpha0 = 1.058791184e-28 palpha0 = -1.005851625e-32
+ alpha1 = 0.85
+ beta0 = 1.042942088e+01 lbeta0 = 6.696082211e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.901361166e-01 lkt1 = 1.099223579e-7
+ kt2 = -6.838621167e-02 lkt2 = 3.927495052e-8
+ at = 1.538056803e+05 lat = -8.673316007e-2
+ ute = -2.354634327e+00 lute = 1.218431122e-6
+ ua1 = -1.525599643e-09 lua1 = 2.672085355e-15 pua1 = -3.308722450e-36
+ ub1 = 9.327016030e-19 lub1 = -1.525925138e-24 wub1 = -7.703719778e-40 pub1 = 7.703719778e-46
+ uc1 = 7.140092441e-11 luc1 = -2.892326820e-17 wuc1 = 2.067951531e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.149 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.137264256e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.044458513e-8
+ k1 = 6.257710813e-01 lk1 = -6.813779451e-8
+ k2 = -5.660819148e-02 lk2 = 2.114635860e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.145343276e-01 ldsub = 4.327790973e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.265594374e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.716768506e-9
+ nfactor = 3.816562506e+00 lnfactor = -3.622288970e-7
+ eta0 = -4.380244824e-01 leta0 = 4.193566311e-07 weta0 = -3.191891196e-22 peta0 = -1.387778781e-29
+ etab = -1.600650675e-01 letab = 7.204793714e-8
+ u0 = 3.099996783e-02 lu0 = -3.684596026e-9
+ ua = -8.551569684e-10 lua = -2.682768385e-16
+ ub = 1.911412760e-18 lub = 1.068460154e-25
+ uc = 2.781855419e-11 luc = 1.116979601e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.042946423e+04 lvsat = 4.091806665e-2
+ a0 = 1.033165535e+00 la0 = 1.588065576e-7
+ ags = 2.238489688e+00 lags = -9.409245522e-07 wags = 7.105427358e-21
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 5.649984864e-07 lb0 = -2.553120810e-13
+ b1 = 1.381407782e-08 lb1 = -6.242319301e-15
+ keta = -1.128952678e-01 lketa = 4.780085547e-08 wketa = -2.220446049e-22
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.248591510e+00 lpclm = -3.600504255e-7
+ pdiblc1 = 6.447801385e-01 lpdiblc1 = -2.764374541e-7
+ pdiblc2 = 8.895504640e-03 lpdiblc2 = -3.998725233e-9
+ pdiblcb = 8.513601993e-02 lpdiblcb = -8.122164672e-08 wpdiblcb = 6.678685383e-23 ppdiblcb = -5.724587471e-29
+ drout = 8.471347030e-01 ldrout = 6.907687808e-8
+ pscbe1 = 1.002269402e+09 lpscbe1 = -2.554584480e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 6.984094440e-06 lalpha0 = -1.393643680e-12
+ alpha1 = 0.85
+ beta0 = 1.696331585e+01 lbeta0 = 4.765917275e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.707775674e-01 lkt1 = -3.692777231e-9
+ kt2 = -1.845629469e-02 lkt2 = -8.252388786e-9
+ at = 1.097132703e+05 lat = -4.476243274e-2
+ ute = -8.616208325e-01 lute = -2.027400562e-7
+ ua1 = 1.688160728e-09 lua1 = -3.870320811e-16
+ ub1 = -7.051401785e-19 lub1 = 3.310533460e-26
+ uc1 = 7.289584949e-11 luc1 = -3.034625897e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.150 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.912784230e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.459968901e-8
+ k1 = 1.260614572e-01 lk1 = 1.576714902e-7
+ k2 = 9.145896450e-02 lk2 = -4.576237591e-08 pk2 = -3.469446952e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.905328527e-01 ldsub = 5.412372020e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.103590353e-03 lcdscd = -1.221701112e-09 pcdscd = 3.469446952e-30
+ cit = 0.0
+ voff = {-1.154994110e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.271458428e-8
+ nfactor = 3.206634077e+00 lnfactor = -8.661382847e-8
+ eta0 = 8.851262252e-01 leta0 = -1.785500338e-7
+ etab = 3.439973846e-02 letab = -1.582701384e-08 wetab = 2.428612866e-23 petab = -9.540979118e-30
+ u0 = 1.738280483e-02 lu0 = 2.468741208e-9
+ ua = -1.664072323e-09 lua = 9.725664078e-17
+ ub = 2.065347197e-18 lub = 3.728596771e-26
+ uc = 2.021746693e-11 luc = 1.460458292e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.233335552e+05 lvsat = 3.455283115e-3
+ a0 = 1.291411731e+00 la0 = 4.211000830e-8
+ ags = -7.269793749e-01 lags = 3.991145732e-07 pags = 3.330669074e-28
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 5.428652140e-02 lketa = -2.774541861e-08 wketa = 2.775557562e-23 pketa = 2.081668171e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.240064177e-01 lpclm = -7.781228943e-8
+ pdiblc1 = -2.285578199e-01 lpdiblc1 = 1.182073759e-07 wpdiblc1 = -2.220446049e-22 ppdiblc1 = 5.551115123e-29
+ pdiblc2 = -6.704200070e-03 lpdiblc2 = 3.050484931e-09 wpdiblc2 = 4.770489559e-24 ppdiblc2 = -3.415236843e-30
+ pdiblcb = -8.758737422e-02 lpdiblcb = -3.171226649e-9
+ drout = 1.401075462e+00 ldrout = -1.812384259e-7
+ pscbe1 = 1.507016602e+08 lpscbe1 = 1.293488349e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.031901081e-06 lalpha0 = -1.415246593e-12
+ alpha1 = 0.85
+ beta0 = 2.100422375e+01 lbeta0 = -1.349417775e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.096264800e-01 lkt1 = 1.386230826e-8
+ kt2 = -4.304931441e-02 lkt2 = 2.860729557e-9
+ at = -3.932844369e+03 lat = 6.592087190e-3
+ ute = -1.303201517e+00 lute = -3.198134717e-9
+ ua1 = 1.522520004e-09 lua1 = -3.121821851e-16
+ ub1 = -1.713664128e-18 lub1 = 4.888381454e-25 wub1 = -3.081487911e-39
+ uc1 = -1.084804678e-10 luc1 = 5.161425266e-17 wuc1 = -1.033975766e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.151 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {6.130803429e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.900108240e-8
+ k1 = 9.070734896e-01 lk1 = 5.143085957e-17
+ k2 = -1.611477193e-01 lk2 = 5.234114019e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -7.794653811e-18
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999996e-03 lcdscd = 5.442070405e-19
+ cit = 0.0
+ voff = {-1.237493848e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.104907131e-8
+ nfactor = 2.484263783e+00 lnfactor = 5.921900879e-8
+ eta0 = 2.001909455e-03 leta0 = -2.640137943e-10
+ etab = -4.399800002e-02 letab = 2.220501560e-18
+ u0 = 2.919169366e-02 lu0 = 8.475092343e-11
+ ua = -1.224106221e-09 lua = 8.435844238e-18
+ ub = 2.103521860e-18 lub = 2.957922859e-26
+ uc = 1.218677263e-10 luc = -5.916673095e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.325369855e+05 lvsat = 1.597285411e-3
+ a0 = 1.499999999e+00 la0 = 1.571063279e-16
+ ags = 1.250000000e+00 lags = 3.363886947e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -6.898412508e-08 lb0 = 1.392658415e-14
+ b1 = 9.858632274e-11 lb1 = -1.990270542e-17
+ keta = -1.889316341e-01 lketa = 2.135570583e-08 pketa = 5.551115123e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.499568007e-01 lpclm = -2.248687870e-8
+ pdiblc1 = 3.569721502e-01 lpdiblc1 = -2.689581891e-17
+ pdiblc2 = 8.406112095e-03 lpdiblc2 = 7.211592434e-19
+ pdiblcb = -1.032957700e-01 lpdiblcb = 2.135180921e-18
+ drout = 5.033266589e-01 ldrout = 1.424540486e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 1.407337189e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 5.774280622e-09 lalpha0 = 3.194912098e-15
+ alpha1 = 0.85
+ beta0 = 1.518074234e+01 lbeta0 = -1.737675240e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.585636645e-01 lkt1 = 3.553695993e-9
+ kt2 = -2.887893901e-02 lkt2 = 8.535394613e-19
+ at = -1.837987011e+04 lat = 9.508667194e-3
+ ute = -1.325229293e+00 lute = 1.248854588e-9
+ ua1 = -2.384733722e-11 lua1 = 1.610623533e-25
+ ub1 = 7.077531683e-19 lub1 = 2.287973959e-34
+ uc1 = 1.471862500e-10 luc1 = -3.312858353e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.152 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {-7.424725632e-02+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.164436871e-08 wvth0 = 4.882898279e-07 pvth0 = -6.439615079e-14
+ k1 = 0.90707349
+ k2 = -3.400228006e-01 lk2 = 2.882433862e-08 wk2 = 8.695896763e-08 pk2 = -1.146823561e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.305277426e+00 ldsub = -2.435377092e-07 wdsub = -1.053613991e-06 pdsub = 1.389516668e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000001e-03 lcdscd = -9.108686028e-20
+ cit = 0.0
+ voff = {-2.075300001e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.193267707e-17
+ nfactor = -6.851267237e-01 lnfactor = 4.772013983e-07 wnfactor = 1.671005376e-06 pnfactor = -2.203738600e-13
+ eta0 = -1.034739498e-02 leta0 = 1.364624824e-09 weta0 = 4.559393272e-09 peta0 = -6.012973441e-16
+ etab = -0.043998
+ u0 = 1.106030932e-01 lu0 = -1.065186585e-08 wu0 = -4.198915474e-08 pu0 = 5.537571716e-15
+ ua = -2.896658749e-09 lua = 2.290137441e-16 wua = 7.848765503e-16 pua = -1.035103043e-22
+ ub = 1.246658459e-17 lub = -1.337111847e-24 wub = -5.386694525e-24 pub = 7.104026606e-31
+ uc = -1.739688444e-10 luc = 3.309854969e-17 wuc = 1.228498853e-16 puc = -1.620156572e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.391586935e+05 lvsat = 7.240079398e-04 wvsat = 1.235534015e-02 pvsat = -1.629434615e-9
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -9.545565207e-06 lb0 = 1.263707574e-12 wb0 = 4.651149284e-12 pb0 = -6.133982187e-19
+ b1 = 1.211326448e-08 lb1 = -1.604410475e-15 wb1 = -3.961348637e-14 pb1 = 5.224266196e-21
+ keta = -7.798050099e-01 lketa = 9.928067751e-08 wketa = 4.295746201e-07 pketa = -5.665273047e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 8.437561931e-03 lpclm = 2.255302003e-08 wpclm = 1.287412004e-07 ppclm = -1.697851824e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.000000000e-08 lalpha0 = -9.147955830e-26 walpha0 = 2.270014417e-22 palpha0 = -2.993721485e-29
+ alpha1 = 0.85
+ beta0 = 1.390773688e+01 lbeta0 = -5.882291189e-09 wbeta0 = 4.115463526e-17 pbeta0 = -5.428546501e-24
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.998872496e-01 lkt1 = -4.184608273e-09 wkt1 = -8.445688593e-17 pkt1 = 1.113820147e-23
+ kt2 = -0.028878939
+ at = 5.372048694e+04 lat = 6.223330274e-12 wat = -2.680905163e-11 pat = 3.535533324e-18
+ ute = -1.119309967e+00 lute = -2.590799196e-08 wute = -2.297333057e-07 pute = 3.029745809e-14
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.153 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {0.4913699+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56800772
+ k2 = -0.040590746
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 2.78042
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.025731
+ ua = -1.0529435e-9
+ ub = 1.832e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 9.1484e-8
+ b1 = 1.6098e-9
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.154 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.471672731e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.819255524e-07 wvth0 = 1.524718189e-08 pvth0 = -3.042099587e-13
+ k1 = 8.566922029e-01 lk1 = -5.759798448e-06 wk1 = -1.321818023e-07 pk1 = 2.637275589e-12
+ k2 = -1.610472924e-01 lk2 = 2.403334679e-06 wk2 = 5.607514373e-08 pk2 = -1.118804595e-12
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.013776050e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.376726686e-07 wvoff = -1.776848878e-10 pvoff = 3.545147736e-15
+ nfactor = 3.864774810e+00 lnfactor = -2.163491814e-05 wnfactor = -4.677804086e-07 pnfactor = 9.333099047e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.058376774e-02 lu0 = 1.026969655e-07 wu0 = 1.845674936e-09 pu0 = -3.682468669e-14
+ ua = -1.676520142e-09 lua = 1.244152696e-14 wua = 2.356368865e-16 pua = -4.701399119e-21
+ ub = 2.292847676e-18 lub = -9.194777996e-24 wub = -1.844806717e-25 pub = 3.680736409e-30
+ uc = 6.321093241e-11 luc = -2.927725532e-16 wuc = 2.683584837e-20 puc = -5.354256531e-25
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.005405322e+00 la0 = 7.126705702e-06 wa0 = 2.083724697e-07 pa0 = -4.157422718e-12
+ ags = 3.183979180e-01 lags = 5.283673481e-07 wags = 1.373364005e-09 pags = -2.740119519e-14
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.376251231e-07 lb0 = -9.206021975e-13 wb0 = -2.615232352e-14 pb0 = 5.217880468e-19
+ b1 = 4.385568931e-09 lb1 = -5.538181139e-14 wb1 = -1.199120420e-15 pb1 = 2.392470792e-20
+ keta = -5.705121375e-03 lketa = 2.311468062e-08 wketa = 1.642985352e-09 pketa = -3.278064822e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.820098972e-02 lpclm = -1.024050039e-06 wpclm = -4.207861024e-08 ppclm = 8.395474241e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 3.656782392e-03 lpdiblc2 = -5.379934793e-08 wpdiblc2 = -1.678058385e-09 ppdiblc2 = 3.348042121e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -1.083126458e+08 lpscbe1 = 6.650214244e+03 wpscbe1 = 1.898571550e+01 ppscbe1 = -3.788007364e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.038984879e-01 lkt1 = 3.495267863e-07 wkt1 = 1.117634155e-08 pkt1 = -2.229890367e-13
+ kt2 = -6.617993721e-02 lkt2 = 7.314759852e-07 wkt2 = 1.661549918e-08 pkt2 = -3.315104624e-13
+ at = 2.419911516e+05 lat = -1.336599485e+00 wat = -2.367868973e-02 pat = 4.724343998e-7
+ ute = -5.417201598e-01 lute = -1.144599190e-05 wute = -2.565191388e-07 pute = 5.118039331e-12
+ ua1 = 1.702889580e-09 lua1 = -1.160979165e-14 wua1 = -3.637046743e-16 pua1 = 7.256592381e-21
+ ub1 = -9.727310539e-19 lub1 = 8.045816560e-24 wub1 = 3.186993780e-25 pub1 = -6.358652065e-30
+ uc1 = 1.840775064e-10 luc1 = -2.997952568e-15 wuc1 = -6.210524725e-17 puc1 = 1.239116503e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.155 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.175091453e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 3.225753551e-07 wvth0 = -4.049911288e-11 pvth0 = -1.826441386e-13
+ k1 = -3.109066945e-01 lk1 = 3.524809039e-06 wk1 = 4.045265681e-07 pk1 = -1.630565504e-12
+ k2 = 3.227172860e-01 lk2 = -1.443503680e-06 wk2 = -1.696409798e-07 pk2 = 6.760631593e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-8.298215126e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.839511273e-07 wvoff = -1.893147719e-08 pvoff = 1.526730724e-13
+ nfactor = -1.200015267e+00 lnfactor = 1.863968984e-05 wnfactor = 1.538009863e-06 pnfactor = -6.616706507e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.292991545e-02 lu0 = 4.521868088e-09 wu0 = -3.106288331e-09 pu0 = 2.552735932e-15
+ ua = 1.335033509e-10 lua = -1.951564464e-15 wua = -6.007883483e-16 pua = 1.949754814e-21
+ ub = 8.146667534e-19 lub = 2.559540799e-24 wub = 5.543881384e-25 pub = -2.194660444e-30
+ uc = -9.087236242e-11 luc = 9.324794714e-16 wuc = 5.437335560e-17 puc = -4.326924835e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 2.303990104e+00 la0 = -3.199485948e-06 wa0 = -4.839049878e-07 pa0 = 1.347485243e-12
+ ags = 1.613650989e-01 lags = 1.777073639e-06 wags = 1.079790350e-07 pags = -8.751168048e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -2.737004915e-07 lb0 = 2.350210142e-12 wb0 = 1.750627414e-13 pb0 = -1.078250205e-18
+ b1 = -1.641762318e-08 lb1 = 1.100426967e-13 wb1 = 7.979418042e-15 pb1 = -4.906193768e-20
+ keta = -9.589209499e-03 lketa = 5.400048717e-08 wketa = -4.224070720e-09 pketa = 1.387348348e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.220237848e+00 lpclm = 1.717334327e-05 wpclm = 8.273084310e-07 ppclm = -6.073714871e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -4.261137358e-03 lpdiblc2 = 9.163007692e-09 wpdiblc2 = 1.425870181e-09 ppdiblc2 = 8.798350618e-15
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 1.131145246e+09 lpscbe1 = -3.205807414e+03 wpscbe1 = -2.659445869e+02 ppscbe1 = 1.886931121e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.015955838e-01 lkt1 = 3.312143666e-07 wkt1 = 8.269852000e-09 pkt1 = -1.998769776e-13
+ kt2 = 2.885317634e-02 lkt2 = -2.421602487e-08 wkt2 = -2.093006291e-08 pkt2 = -3.295262060e-14
+ at = 8.605503920e+03 lat = 5.192554126e-01 wat = 7.103606920e-02 pat = -2.807260922e-7
+ ute = -3.093466952e+00 lute = 8.845194932e-06 wute = 1.006794284e-06 pute = -4.927678672e-12
+ ua1 = -2.333282128e-09 lua1 = 2.048536547e-14 wua1 = 2.080142285e-15 pua1 = -1.217658782e-20
+ ub1 = 1.873747470e-18 lub1 = -1.458904193e-23 wub1 = -1.567900949e-24 pub1 = 8.643369228e-30
+ uc1 = -3.312308027e-10 luc1 = 1.099717784e-15 wuc1 = 1.407496707e-16 puc1 = -3.739616654e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.156 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {6.234238611e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -9.598699806e-08 wvth0 = -5.275453823e-08 pvth0 = 2.567547103e-14
+ k1 = 7.211513646e-01 lk1 = -5.537615959e-07 wk1 = -8.753677852e-08 pk1 = 3.140102867e-13
+ k2 = -9.151387811e-02 lk2 = 1.934885867e-07 wk2 = 3.139629900e-08 pk2 = -1.184122430e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.142873993e+00 ldsub = -6.255329659e-06 wdsub = -6.974649334e-07 pdsub = 2.756298418e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.491011782e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 3.725314990e-07 wvoff = 6.060120558e-08 pvoff = -1.616306255e-13
+ nfactor = 5.136106937e+00 lnfactor = -6.399911105e-06 wnfactor = -1.047708141e-06 pnfactor = 3.601743345e-12
+ eta0 = 4.994616082e-01 leta0 = -1.657662360e-06 weta0 = -1.848282073e-07 peta0 = 7.304190809e-13
+ etab = -4.366991418e-01 letab = 1.449151371e-06 wetab = 1.615793762e-07 petab = -6.385424669e-13
+ u0 = 3.533449236e-02 lu0 = -4.980733695e-09 wu0 = -3.091539440e-09 pu0 = 2.494450069e-15
+ ua = -1.622843390e-09 lua = 4.989308853e-15 wua = 4.983567606e-16 pua = -2.393935859e-21
+ ub = 3.432101197e-18 lub = -7.784248646e-24 wub = -9.072087046e-25 pub = 3.581396350e-30
+ uc = 2.141712032e-10 luc = -2.730163997e-16 wuc = -9.650447488e-17 puc = 1.635587481e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.724208178e+05 lvsat = -1.155612274e+00 wvsat = -1.580920516e-01 pvsat = 6.247609748e-7
+ a0 = 4.945890435e+00 la0 = -1.363996167e-05 wa0 = -1.805688257e-06 pa0 = 6.571015429e-12
+ ags = -1.523668970e-01 lags = 3.016905152e-06 wags = 2.595401750e-07 pags = -1.474068394e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.081602306e-07 lb0 = 8.411420097e-13 wb0 = -1.538123254e-14 pb0 = -3.256382828e-19
+ b1 = 5.926001712e-08 lb1 = -1.890263321e-13 wb1 = -3.160353276e-14 pb1 = 1.073651735e-19
+ keta = 5.864766441e-02 lketa = -2.156635183e-07 wketa = -3.141195014e-08 pketa = 1.213167476e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 9.261102663e+00 lpclm = -2.819954815e-05 wpclm = -4.405336208e-06 ppclm = 1.460507406e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 1.596771646e-02 lpdiblc2 = -7.077901536e-08 wpdiblc2 = -7.279513782e-09 ppdiblc2 = 4.320099210e-14
+ pdiblcb = -9.095308305e-02 lpdiblcb = 2.606387358e-07 wpdiblcb = 2.906103889e-08 ppdiblcb = -1.148457674e-13
+ drout = 0.56
+ pscbe1 = -1.485804044e+08 lpscbe1 = 1.851516068e+03 wpscbe1 = 4.179748808e+02 ppscbe1 = -8.158372282e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.375267203e-02 lkt1 = -6.482313273e-07 wkt1 = -1.110546229e-07 pkt1 = 2.716791474e-13
+ kt2 = 1.686514935e-01 lkt2 = -5.766823382e-07 wkt2 = -9.926904010e-08 pkt2 = 2.766336949e-13
+ at = 3.016114347e+05 lat = -6.386691582e-01 wat = -7.121116970e-02 pat = 2.814180685e-7
+ ute = 2.345105303e+00 lute = -1.264739543e-05 wute = -1.742929961e-06 pute = 5.938904325e-12
+ ua1 = 1.287983896e-08 lua1 = -3.963507872e-14 wua1 = -5.813695179e-15 pua1 = 1.901891847e-20
+ ub1 = -8.224324439e-18 lub1 = 2.531733658e-23 wub1 = 3.648295973e-24 pub1 = -1.197042028e-29
+ uc1 = -2.086964770e-10 luc1 = 6.154767105e-16 wuc1 = 1.175374693e-16 puc1 = -2.822298076e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.157 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.816549309e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.807290833e-07 wvth0 = -1.738407931e-09 pvth0 = -7.390194440e-14
+ k1 = 4.581635978e-01 lk1 = -4.044077055e-08 wk1 = 7.186909385e-08 pk1 = 2.868993096e-15
+ k2 = -3.260792536e-02 lk2 = 7.851117676e-08 wk2 = -1.376619433e-08 pk2 = -3.026043038e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -2.320183686e+00 ldsub = 2.456027828e-06 wdsub = 1.394929867e-06 pdsub = -1.327807236e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {7.783411229e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.656072827e-07 wvoff = -7.758368570e-08 pvoff = 1.080898383e-13
+ nfactor = 2.903120190e+00 lnfactor = -2.041386702e-06 wnfactor = 1.788620444e-07 pnfactor = 1.207624305e-12
+ eta0 = -6.851821852e-01 leta0 = 6.546213524e-07 weta0 = 3.696564147e-07 peta0 = -3.518689177e-13
+ etab = 1.029664268e+00 letab = -1.413015508e-06 wetab = -5.137762403e-07 petab = 6.796713292e-13
+ u0 = 2.799688035e-02 lu0 = 9.341411774e-09 wu0 = 1.956968762e-09 pu0 = -7.359637170e-15
+ ua = 2.538813413e-09 lua = -3.133749990e-15 wua = -1.223773276e-15 pua = 9.674570386e-22
+ ub = -3.397676886e-18 lub = 5.546665427e-24 wub = 2.019423833e-24 pub = -2.131042094e-30
+ uc = 1.199030987e-10 luc = -8.901627767e-17 wuc = -3.158199786e-17 puc = 3.683779876e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.197689039e+05 lvsat = -1.949165077e-01 wvsat = 1.062435293e-01 pvsat = 1.088093770e-7
+ a0 = -3.870141616e+00 la0 = 3.567883785e-06 wa0 = 2.366256240e-06 pa0 = -1.572123768e-12
+ ags = -2.864834008e+00 lags = 8.311318169e-06 wags = 1.408322821e-06 pags = -3.716355414e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -7.733340500e-07 lb0 = 2.561713948e-12 wb0 = 4.785846827e-13 pb0 = -1.289800967e-18
+ b1 = -6.994816881e-08 lb1 = 6.317267105e-14 wb1 = 4.010129984e-14 pb1 = -3.259412684e-20
+ keta = 2.959942880e-01 lketa = -6.789358833e-07 wketa = -1.224711267e-07 pketa = 2.990534241e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.025912804e+01 lpclm = 9.901619287e-06 wpclm = 5.632097138e-06 ppclm = -4.986801378e-12
+ pdiblc1 = 1.409731587e+00 lpdiblc1 = -1.990394709e-06 wpdiblc1 = -5.329628678e-07 ppdiblc1 = 1.040280095e-12
+ pdiblc2 = -3.928374224e-02 lpdiblc2 = 3.706525711e-08 wpdiblc2 = 2.639887502e-08 ppdiblc2 = -2.253521512e-14
+ pdiblcb = -2.076266460e-02 lpdiblcb = 1.236353916e-07 wpdiblcb = -1.867105572e-09 ppdiblcb = -5.447770989e-14
+ drout = -8.958948241e-01 ldrout = 2.841733445e-06 wdrout = 6.019936659e-07 pdrout = -1.175019999e-12
+ pscbe1 = 1.140176721e+09 lpscbe1 = -6.639844782e+02 wpscbe1 = -1.498927489e+02 ppscbe1 = 2.925728086e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -2.822249135e-05 lalpha0 = 5.514550107e-11 walpha0 = 1.244895177e-11 palpha0 = -2.429887243e-17
+ alpha1 = 0.85
+ beta0 = -4.686808530e+00 lbeta0 = 3.620116318e-05 wbeta0 = 8.172317336e-06 pbeta0 = -1.595139093e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.811288910e-01 lkt1 = 3.811442944e-07 wkt1 = 1.032568056e-07 pkt1 = -1.466312580e-13
+ kt2 = -2.188761621e-01 lkt2 = 1.797255298e-07 wkt2 = 8.135968290e-08 pkt2 = -7.593207757e-14
+ at = 1.726950026e+05 lat = -3.870396237e-01 wat = -1.021217208e-02 pat = 1.623552840e-7
+ ute = -5.556134448e+00 lute = 2.774884315e-06 wute = 1.730833414e-06 pute = -8.414684031e-13
+ ua1 = -1.188656088e-08 lua1 = 8.705986572e-15 wua1 = 5.601467196e-15 pua1 = -3.262120083e-21
+ ub1 = 6.998076834e-18 lub1 = -4.394979236e-24 wub1 = -3.279135942e-24 pub1 = 1.551102455e-30
+ uc1 = 1.965415887e-10 luc1 = -1.754997703e-16 wuc1 = -6.765504760e-17 puc1 = 7.924394749e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.158 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {6.760090244e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.272885632e-09 wvth0 = -8.773516599e-08 pvth0 = 7.956735655e-15
+ k1 = 7.623533543e-01 lk1 = -3.299932202e-07 wk1 = -7.384074741e-08 pk1 = 1.415674225e-13
+ k2 = -4.385854157e-02 lk2 = 8.922042456e-08 wk2 = -6.892868728e-09 pk2 = -3.680301843e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.942889723e-01 ldsub = 6.254907872e-08 wdsub = 1.094528689e-08 pdsub = -1.041861063e-14
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.113151175e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 9.628375284e-09 wvoff = 4.582163286e-08 pvoff = -9.377339777e-15
+ nfactor = 4.908733100e-01 lnfactor = 2.547852711e-07 wnfactor = 1.797974002e-06 pnfactor = -3.335776037e-13
+ eta0 = -4.380244824e-01 leta0 = 4.193566311e-07 weta0 = -5.551115123e-23 peta0 = -4.076600169e-29
+ etab = -8.639860007e-01 letab = 3.895142035e-07 wetab = 3.805621820e-07 petab = -1.716324225e-13
+ u0 = 6.090244917e-02 lu0 = -2.198077398e-08 wu0 = -1.616623829e-08 pu0 = 9.891499282e-15
+ ua = 1.020357730e-09 lua = -1.688360876e-15 wua = -1.013963262e-15 pua = 7.677428735e-22
+ ub = 1.630857885e-18 lub = 7.600987209e-25 wub = 1.516769429e-25 pub = -3.531693167e-31
+ uc = -1.889255727e-10 luc = 2.049518669e-16 wuc = 1.171788108e-16 puc = -1.047647885e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -4.604561892e+05 lvsat = 1.293772462e-01 wvsat = 2.707948126e-01 pvsat = -4.782386315e-8
+ a0 = -1.023856506e+00 la0 = 8.585590683e-07 wa0 = 1.112091940e-06 pa0 = -3.783085994e-13
+ ags = 1.048301117e+01 lags = -4.394242047e-06 wags = -4.457252138e-06 pags = 1.866973944e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 5.035857133e-06 lb0 = -2.967944765e-12 wb0 = -2.417089252e-12 pb0 = 1.466536033e-18
+ b1 = 1.485216016e-08 lb1 = -1.754715090e-14 wb1 = -5.612205319e-16 pb1 = 6.111753716e-21
+ keta = -7.665833767e-01 lketa = 3.325116068e-07 wketa = 3.534047097e-07 pketa = -1.539237429e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.383932145e-01 lpclm = -3.763360469e-07 wpclm = 3.839559248e-07 ppclm = 8.804528095e-15
+ pdiblc1 = 5.314791804e-01 lpdiblc1 = -1.154402930e-06 wpdiblc1 = 6.125412354e-08 ppdiblc1 = 4.746562314e-13
+ pdiblc2 = 4.393337293e-03 lpdiblc2 = -4.510125042e-09 wpdiblc2 = 2.434015737e-09 ppdiblc2 = 2.764791015e-16
+ pdiblcb = 5.704305673e-01 lpdiblcb = -4.391102131e-07 wpdiblcb = -2.623657617e-07 ppdiblcb = 1.934860114e-13
+ drout = 3.074134857e+00 ldrout = -9.372623775e-07 wdrout = -1.203987547e-06 pdrout = 5.440592044e-13
+ pscbe1 = 1.893533116e+09 lpscbe1 = -1.381090117e+03 wpscbe1 = -4.818456838e+02 ppscbe1 = 6.085525003e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.989595066e-05 lalpha0 = -9.695149631e-12 walpha0 = -1.779320265e-11 palpha0 = 4.488059765e-18
+ alpha1 = 0.85
+ beta0 = 3.756665892e+01 lbeta0 = -4.019109669e-06 wbeta0 = -1.113882657e-05 pbeta0 = 2.430520037e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.989481820e-01 lkt1 = 1.735373893e-08 wkt1 = -3.883326428e-08 pkt1 = -1.137842012e-14
+ kt2 = -7.647180110e-02 lkt2 = 4.417352420e-08 wkt2 = 3.136503926e-08 pkt2 = -2.834312619e-14
+ at = -4.973709475e+05 lat = 2.507834229e-01 wat = 3.282091548e-01 pat = -1.597815470e-7
+ ute = -4.537414384e+00 lute = 1.805184042e-06 wute = 1.987251619e-06 pute = -1.085548021e-12
+ ua1 = -7.772818846e-09 lua1 = 4.790193690e-15 wua1 = 5.114908309e-15 pua1 = -2.798973923e-21
+ ub1 = 7.831139534e-18 lub1 = -5.187955792e-24 wub1 = -4.614985974e-24 pub1 = 2.822672719e-30
+ uc1 = 4.185163483e-10 luc1 = -3.867933265e-16 wuc1 = -1.868535015e-16 puc1 = 1.927066910e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.159 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {8.257382321e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.193266975e-08 wvth0 = -1.267564755e-07 pvth0 = 2.558972404e-14
+ k1 = -6.744845092e-01 lk1 = 3.192865104e-07 wk1 = 4.328007669e-07 pk1 = -8.737425162e-14
+ k2 = 3.868005265e-01 lk2 = -1.053862258e-07 wk2 = -1.596710994e-07 pk2 = 3.223456121e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.310235632e-01 ldsub = 4.594941508e-08 wdsub = -2.189057378e-08 pdsub = 4.419290925e-15
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.103590353e-03 lcdscd = -1.221701112e-09 wcdscd = 3.469446952e-24
+ cit = 0.0
+ voff = {-1.993167618e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 4.206546323e-09 wvoff = 4.531434201e-08 pvoff = -9.148104679e-15
+ nfactor = -3.365722895e-01 lnfactor = 6.286922160e-07 wnfactor = 1.915570744e-06 pnfactor = -3.867173375e-13
+ eta0 = 8.851262252e-01 leta0 = -1.785500338e-7
+ etab = 3.191082310e-02 letab = -1.532454912e-08 wetab = 1.345587289e-09 petab = -2.716485075e-16
+ u0 = -1.752454325e-03 lu0 = 6.331786462e-09 wu0 = 1.034513343e-08 pu0 = -2.088485882e-15
+ ua = -3.954370644e-09 lua = 5.596243562e-16 wua = 1.238208562e-15 pua = -2.499707827e-22
+ ub = 4.171248350e-18 lub = -3.878554630e-25 wub = -1.138517552e-24 pub = 2.298450619e-31
+ uc = 4.035755392e-10 luc = -6.278812807e-17 wuc = -2.072556413e-16 puc = 4.184097613e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -4.281925666e+05 lvsat = 1.147979281e-01 wvsat = 2.981726703e-01 pvsat = -6.019539685e-8
+ a0 = 3.723050666e-01 la0 = 2.276601808e-07 wa0 = 4.968984740e-07 pa0 = -1.003143608e-13
+ ags = 3.619210950e-01 lags = 1.792862574e-07 wags = -5.886944389e-07 pags = 1.188462220e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -2.769346431e-06 lb0 = 5.590784269e-13 wb0 = 1.497197300e-12 pb0 = -3.022556881e-19
+ b1 = -4.334296764e-08 lb1 = 8.750121651e-15 wb1 = 2.343259528e-14 pb1 = -4.730595768e-21
+ keta = 1.157258111e-02 lketa = -1.912228563e-08 wketa = 2.309252296e-08 pketa = -4.661941628e-15
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.248365317e-01 lpclm = 1.944934740e-07 wpclm = 7.292276614e-07 ppclm = -1.472172095e-13
+ pdiblc1 = -3.945213926e+00 lpdiblc1 = 8.685296273e-07 wpdiblc1 = 2.009343224e-06 ppdiblc1 = -4.056482194e-13
+ pdiblc2 = -1.688757484e-02 lpdiblc2 = 5.106314812e-09 wpdiblc2 = 5.505458267e-09 ppdiblc2 = -1.111447420e-15
+ pdiblcb = -6.419600984e-01 lpdiblcb = 1.087460933e-07 wpdiblcb = 2.997116346e-07 ppdiblcb = -6.050608451e-14
+ drout = 1.401074665e+00 ldrout = -1.812382651e-07 wdrout = 4.305879324e-13 pdrout = -8.692752229e-20
+ pscbe1 = -2.740844462e+09 lpscbe1 = 7.130970577e+02 wpscbe1 = 1.563262363e+03 ppscbe1 = -3.155929692e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.331484728e-05 lalpha0 = -6.721274054e-12 walpha0 = -1.420940177e-11 palpha0 = 2.868608239e-18
+ alpha1 = 0.85
+ beta0 = 4.026245524e+01 lbeta0 = -5.237288807e-06 wbeta0 = -1.041161621e-05 pbeta0 = 2.101907491e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -9.560707741e-02 lkt1 = -2.934414276e-08 wkt1 = -1.157057377e-07 pkt1 = 2.335879003e-14
+ kt2 = 6.178991731e-02 lkt2 = -1.830431938e-08 wkt2 = -5.667944352e-08 pkt2 = 1.144250274e-14
+ at = 8.093128452e+04 lat = -1.054036801e-02 wat = -4.588026373e-02 pat = 9.262353522e-9
+ ute = 8.440981305e-02 lute = -2.833304977e-07 wute = -7.501870888e-07 pute = 1.514485197e-13
+ ua1 = 5.130475444e-09 lua1 = -1.040559837e-15 wua1 = -1.950576165e-15 pua1 = 3.937842669e-22
+ ub1 = -7.168378183e-18 lub1 = 1.590041274e-24 wub1 = 2.948992969e-24 pub1 = -5.953456496e-31
+ uc1 = -9.095513914e-10 luc1 = 2.133352518e-16 wuc1 = 4.330845756e-16 puc1 = -8.743154720e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.160 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {2.764771980e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.895269710e-08 wvth0 = 1.819784314e-07 pvth0 = -3.673798772e-14
+ k1 = 9.070734896e-01 lk1 = 5.142908321e-17
+ k2 = -1.824697962e-01 lk2 = 9.538636231e-09 wk2 = 1.152739709e-08 pk2 = -2.327162452e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.829219179e+00 ldsub = -2.766959140e-07 wdsub = -7.409843688e-07 pdsub = 1.495906653e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999994e-03 lcdscd = 8.850576522e-19 wcdscd = 9.127889417e-19 pcdscd = -1.842744707e-25
+ cit = 0.0
+ voff = {-1.237493846e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.104907136e-08 wvoff = -1.195763488e-16 pvoff = 2.414018985e-23
+ nfactor = -8.852587839e+00 lnfactor = 2.347913951e-06 wnfactor = 6.129064766e-06 pnfactor = -1.237341724e-12
+ eta0 = 2.001907991e-03 leta0 = -2.640134585e-10 weta0 = 8.993474368e-16 peta0 = -1.815611599e-22
+ etab = -4.399800002e-02 letab = 2.220584827e-18
+ u0 = -1.200339756e-02 lu0 = 8.401257133e-09 wu0 = 2.227138455e-08 pu0 = -4.496169385e-15
+ ua = -1.124955223e-09 lua = -1.158085845e-17 wua = -5.360420252e-17 pua = 1.082167001e-23
+ ub = 2.968635726e-18 lub = -1.450708236e-25 wub = -4.677082392e-25 pub = 9.442140704e-32
+ uc = 2.418669184e-10 luc = -3.014222999e-17 wuc = -6.487540321e-17 puc = 1.309711128e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.995282079e+05 lvsat = -7.249126955e-02 wvsat = -1.984071985e-01 pvsat = 4.005464365e-8
+ a0 = 1.499999999e+00 la0 = 1.571058839e-16
+ ags = 1.250000000e+00 lags = 3.363753720e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 8.513050088e-06 lb0 = -1.718623065e-12 wb0 = -4.639722321e-12 pb0 = 9.366717818e-19
+ b1 = 1.364877983e-07 lb1 = -2.755429320e-14 wb1 = -7.373637243e-14 pb1 = 1.488597260e-20
+ keta = -5.324173871e-01 lketa = 9.069895314e-08 wketa = 1.856993897e-07 pketa = -3.748917848e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.640865481e-01 lpclm = -2.533940623e-08 wpclm = -7.638993597e-09 ppclm = 1.542167666e-15
+ pdiblc1 = 3.569721502e-01 lpdiblc1 = -2.689615197e-17
+ pdiblc2 = 8.406112095e-03 lpdiblc2 = 7.211453656e-19
+ pdiblcb = -1.032957700e-01 lpdiblcb = 2.135291943e-18
+ drout = 5.033266589e-01 ldrout = 1.424533824e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 1.407337189e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.850881889e-07 lalpha0 = -3.300515901e-14 walpha0 = -9.694283684e-14 palpha0 = 1.957091684e-20
+ alpha1 = 0.85
+ beta0 = 1.963757411e+01 lbeta0 = -1.073517178e-06 wbeta0 = -2.409505872e-06 pbeta0 = 4.864334550e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.700963859e-01 lkt1 = -1.430616667e-08 wkt1 = -4.782824173e-08 pkt1 = 9.655613269e-15
+ kt2 = -2.887893901e-02 lkt2 = 8.536088503e-19
+ at = -1.013955683e+05 lat = 2.626795935e-02 wat = 4.488094292e-02 pat = -9.060609638e-9
+ ute = -1.020424404e+00 lute = -6.028546117e-08 wute = -1.647872766e-07 pute = 3.326742019e-14
+ ua1 = -2.384733722e-11 lua1 = 1.610623275e-25
+ ub1 = 7.077531683e-19 lub1 = 2.287968181e-34
+ uc1 = 1.471862500e-10 luc1 = -3.312806654e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.161 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {1.805991071e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.627611220e-07 wvth0 = -5.282271796e-07 pvth0 = 5.692463847e-14
+ k1 = 0.90707349
+ k2 = -1.669940782e-01 lk2 = 7.497683066e-09 wk2 = -6.585896600e-09 pk2 = 6.163683312e-17
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -8.214264315e-01 ldsub = 7.287387975e-08 wdsub = 6.367821687e-07 pdsub = -3.211056338e-14
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000005e-03 lcdscd = -4.924515656e-19 wcdscd = -2.129837973e-18 pcdscd = 2.169900544e-25
+ cit = 0.0
+ voff = {-2.075300006e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 6.451184031e-17 wvoff = 2.790114806e-16 pvoff = -2.842598379e-23
+ nfactor = 2.576752691e+01 lnfactor = -2.217821402e-06 wnfactor = -1.263014566e-05 pnfactor = 1.236641707e-12
+ eta0 = -1.034739468e-02 leta0 = 1.364625037e-09 weta0 = 4.559393667e-09 peta0 = -6.012974591e-16
+ etab = -0.043998
+ u0 = 1.224977328e-01 lu0 = -9.336886445e-09 wu0 = -4.841977758e-08 pu0 = 4.826651768e-15
+ ua = -3.128056175e-09 lua = 2.525900982e-16 wua = 9.099774036e-16 pua = -1.162564358e-22
+ ub = 1.044798401e-17 lub = -1.131454754e-24 wub = -4.295374454e-24 pub = 5.992178552e-31
+ uc = -4.622848178e-10 luc = 6.272200513e-17 wuc = 2.787227266e-16 puc = -3.221695368e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -7.488089811e+05 lvsat = 9.214068726e-02 wvsat = 4.924190800e-01 pvsat = -5.105221679e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -2.957033937e-05 lb0 = 3.303852420e-12 wb0 = 1.547718299e-11 pb0 = -1.716365807e-18
+ b1 = -3.061265163e-07 lb1 = 3.081812522e-14 wb1 = 1.324371228e-13 pb1 = -1.230439412e-20
+ keta = 2.166194943e-02 lketa = 1.762641616e-08 wketa = -3.724065077e-09 pketa = -1.250782385e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.453138342e-02 lpclm = 2.591191519e-08 wpclm = 1.465652672e-07 ppclm = -1.879444445e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -3.883991170e-07 lalpha0 = 4.262692037e-14 walpha0 = 2.261999517e-13 palpha0 = -2.304547725e-20
+ alpha1 = 0.85
+ beta0 = 3.508462771e+00 lbeta0 = 1.053606154e-06 wbeta0 = 5.622180360e-06 pbeta0 = -5.727933570e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.063109003e-01 lkt1 = 1.684603971e-08 wkt1 = 1.115992310e-07 pkt1 = -1.136984127e-14
+ kt2 = -0.028878939
+ at = 2.474237824e+05 lat = -1.973468543e-02 wat = -1.047222000e-01 pat = 1.066920246e-8
+ ute = -1.814966711e+00 lute = 4.449957281e-08 wute = 1.463609909e-07 pute = -7.767124470e-15
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.162 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {0.4913699+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56800772
+ k2 = -0.040590746
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 2.78042
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.025731
+ ua = -1.0529435e-9
+ ub = 1.832e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 9.1484e-8
+ b1 = 1.6098e-9
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.163 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.817702567e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.915309403e-7
+ k1 = 5.567098995e-01 lk1 = 2.254127697e-7
+ k2 = -3.378657655e-02 lk2 = -1.357559791e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.017808550e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.296270710e-7
+ nfactor = 2.803162380e+00 lnfactor = -4.537532526e-07 wnfactor = 3.552713679e-21
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.477246701e-02 lu0 = 1.912453613e-8
+ ua = -1.141749888e-09 lua = 1.771854492e-15
+ ub = 1.874174789e-18 lub = -8.414663684e-25
+ uc = 6.327183549e-11 luc = -2.939876843e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.478299869e+00 la0 = -2.308430009e-6
+ ags = 3.215147230e-01 lags = 4.661812263e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 7.827327503e-08 lb0 = 2.635788125e-13
+ b1 = 1.664204119e-09 lb1 = -1.085464512e-15
+ keta = -1.976419529e-03 lketa = -5.127993490e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.729504833e-02 lpclm = 8.812755480e-07 ppclm = -2.220446049e-28
+ pdiblc1 = 0.39
+ pdiblc2 = -1.515165620e-04 lpdiblc2 = 2.218337962e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -6.522518163e+07 lpscbe1 = 5.790538287e+03 ppscbe1 = 3.814697266e-18
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.785341441e-01 lkt1 = -1.565395837e-7
+ kt2 = -2.847160196e-02 lkt2 = -2.087623258e-8
+ at = 1.882531350e+05 lat = -2.644249724e-1
+ ute = -1.123882006e+00 lute = 1.692319823e-7
+ ua1 = 8.774736444e-10 lua1 = 4.858808868e-15
+ ub1 = -2.494531757e-19 lub1 = -6.384937596e-24
+ uc1 = 4.313166665e-11 luc1 = -1.858179462e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.164 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.174172339e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -9.192958009e-8
+ k1 = 6.071532016e-01 lk1 = -1.757063659e-7
+ k2 = -6.227740302e-02 lk2 = 9.079968255e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.259465233e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 6.253544744e-8
+ nfactor = 2.290448121e+00 lnfactor = 3.623289522e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.588029506e-02 lu0 = 1.031521930e-8
+ ua = -1.229966275e-09 lua = 2.473340703e-15
+ ub = 2.072832611e-18 lub = -2.421169734e-24
+ uc = 3.252620055e-11 luc = -4.950205394e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.205783464e+00 la0 = -1.414119935e-7
+ ags = 4.064200086e-01 lags = -2.089755015e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.235987093e-07 lb0 = -9.684364686e-14
+ b1 = 1.691406670e-09 lb1 = -1.301775962e-15
+ keta = -1.917560068e-02 lketa = 8.548590692e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.426882576e-01 lpclm = 3.389244816e-06 wpclm = 2.220446049e-22 ppclm = -4.440892099e-28
+ pdiblc1 = 0.39
+ pdiblc2 = -1.025171335e-03 lpdiblc2 = 2.913057840e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 5.275926511e+08 lpscbe1 = 1.076521426e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.828274235e-01 lkt1 = -1.223999366e-7
+ kt2 = -1.864692104e-02 lkt2 = -9.900092610e-8
+ at = 1.698195537e+05 lat = -1.178433279e-1
+ ute = -8.085800536e-01 lute = -2.338011625e-6
+ ua1 = 2.387533168e-09 lua1 = -7.149004768e-15
+ ub1 = -1.684552764e-18 lub1 = 5.026803557e-24
+ uc1 = -1.180400046e-11 luc1 = 2.510239413e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.165 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.036991516e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.771735122e-8
+ k1 = 5.224894914e-01 lk1 = 1.588745419e-7
+ k2 = -2.026099817e-02 lk2 = -7.524414950e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.115687121e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 5.716048642e-9
+ nfactor = 2.758367370e+00 lnfactor = 1.774128331e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.831834410e-02 lu0 = 6.803396468e-10
+ ua = -4.918389228e-10 lua = -4.436507565e-16
+ ub = 1.373220533e-18 lub = 3.436139465e-25
+ uc = -4.842565427e-12 luc = 9.817486230e-17 puc = -5.169878828e-38
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.363604600e+04 lvsat = 2.622624489e-1
+ a0 = 8.479396350e-01 la0 = 1.272744237e-6
+ ags = 4.366510930e-01 lags = -3.284451492e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 7.325302338e-08 lb0 = 1.021165126e-13
+ b1 = -1.246317312e-08 lb1 = 5.463543899e-14 wb1 = 3.308722450e-30 pb1 = -1.323488980e-35
+ keta = -1.264073531e-02 lketa = 5.966089661e-08 wketa = 3.469446952e-24 pketa = 1.387778781e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.366646536e-01 lpclm = 4.946192650e-6
+ pdiblc1 = 0.39
+ pdiblc2 = -5.529034283e-04 lpdiblc2 = 2.726423184e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.057875285e-01 lkt1 = -3.166433390e-8
+ kt2 = -5.663636600e-02 lkt2 = 5.112883963e-8
+ at = 140000.0
+ ute = -1.610417584e+00 lute = 8.307548749e-7
+ ua1 = -3.141532565e-10 lua1 = 3.527738482e-15 pua1 = -1.654361225e-36
+ ub1 = 5.536467272e-20 lub1 = -1.849143105e-24
+ uc1 = 5.805098873e-11 luc1 = -2.503466317e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.166 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.777096706e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.301102283e-8
+ k1 = 6.212681700e-01 lk1 = -3.392968399e-8
+ k2 = -6.384985590e-02 lk2 = 9.836113722e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.455643000e-01 ldsub = -5.573875314e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-9.823954033e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.030090856e-8
+ nfactor = 3.309041785e+00 lnfactor = 6.992774020e-7
+ eta0 = 1.537410312e-01 leta0 = -1.439337178e-7
+ etab = -1.363342072e-01 letab = 1.294764787e-7
+ u0 = 3.243815733e-02 lu0 = -7.361045536e-9
+ ua = -2.385002539e-10 lua = -9.381376908e-16
+ ub = 1.185339856e-18 lub = 7.103346701e-25
+ uc = 4.822878123e-11 luc = -5.414090889e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.213473320e+05 lvsat = 5.202283627e-2
+ a0 = 1.5
+ ags = 3.313088529e-01 lags = -1.228296323e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.127983295e-07 lb0 = -3.654474191e-13 pb0 = 2.117582368e-34
+ b1 = 2.106042756e-08 lb1 = -1.079864024e-14
+ keta = 1.805004733e-02 lketa = -2.438589030e-10
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.522733322e+00 lpclm = -1.415764330e-6
+ pdiblc1 = 2.001896837e-01 lpdiblc1 = 3.704871499e-7
+ pdiblc2 = 2.062764645e-02 lpdiblc2 = -1.407768104e-8
+ pdiblcb = -0.025
+ drout = 4.703102312e-01 ldrout = 1.750637556e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.467909273e-01 lkt1 = 4.836942111e-8
+ kt2 = -3.423300662e-02 lkt2 = 7.400148129e-9
+ at = 1.495188100e+05 lat = -1.857958438e-2
+ ute = -1.628064281e+00 lute = 8.651991289e-7
+ ua1 = 8.257868283e-10 lua1 = 1.302711089e-15
+ ub1 = -4.438155885e-19 lub1 = -8.748026374e-25
+ uc1 = 4.300065746e-11 luc1 = 4.341792472e-18
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.167 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.768969173e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.378466728e-8
+ k1 = 5.947741785e-01 lk1 = -8.710556888e-9
+ k2 = -5.950168308e-02 lk2 = 5.697170628e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.191289451e-01 ldsub = 3.890438058e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.073244113e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.165319250e-8
+ nfactor = 4.571316858e+00 lnfactor = -5.022582567e-7
+ eta0 = -4.380244824e-01 leta0 = 4.193566311e-07 weta0 = 1.110223025e-22 peta0 = 8.153200337e-29
+ etab = -0.0003125
+ u0 = 2.421369690e-02 lu0 = 4.676620846e-10
+ ua = -1.280798932e-09 lua = 5.400661752e-17
+ ub = 1.975083776e-18 lub = -4.140756249e-26
+ uc = 7.700792919e-11 luc = -3.280841503e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.541038350e+05 lvsat = 2.084254342e-2
+ a0 = 1.5
+ ags = 3.674223382e-01 lags = -1.572053728e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -4.496483497e-07 lb0 = 3.603110884e-13 wb0 = -1.058791184e-28
+ b1 = 1.357848841e-08 lb1 = -3.676724520e-15
+ keta = 3.545712353e-02 lketa = -1.681332400e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.409768704e+00 lpclm = -3.563544566e-7
+ pdiblc1 = 6.704934226e-01 lpdiblc1 = -7.718604331e-08 wpdiblc1 = 8.881784197e-22
+ pdiblc2 = 9.917256884e-03 lpdiblc2 = -3.882664709e-9
+ pdiblcb = -0.025
+ drout = 3.417242576e-01 ldrout = 2.974623007e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -4.851443400e-07 lalpha0 = 4.903561095e-13 walpha0 = -5.293955920e-29 palpha0 = 1.852884572e-34
+ alpha1 = 0.85
+ beta0 = 1.228745412e+01 lbeta0 = 1.496876545e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.870790129e-01 lkt1 = -8.469215655e-9
+ kt2 = -5.289864105e-03 lkt2 = -2.015027931e-8
+ at = 2.474890600e+05 lat = -1.118356039e-1
+ ute = -2.741143519e-02 lute = -6.584319030e-7
+ ua1 = 3.835299287e-09 lua1 = -1.561986640e-15
+ ub1 = -2.642421110e-18 lub1 = 1.218008185e-24
+ uc1 = -5.541599185e-12 luc1 = 5.054824427e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.168 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {-7.528978819e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.695055709e-07 wvth0 = 5.688411126e-07 pvth0 = -2.570484908e-13
+ k1 = 3.077427633e-01 lk1 = 1.209934860e-07 wk1 = -6.585541001e-16 pk1 = 2.975879543e-22
+ k2 = 1.481502145e-01 lk2 = -8.813677649e-08 wk2 = -5.451413507e-08 pk2 = 2.463390187e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.006222508e+00 ldsub = -7.686492458e-07 wdsub = -8.041000353e-07 pdsub = 3.633575280e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.103590367e-03 lcdscd = -1.221701118e-09 wcdscd = -5.978099960e-18 pcdscd = 2.701391194e-24
+ cit = 0.0
+ voff = {-4.175720168e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.285418057e-07 wvoff = 1.414845915e-07 pvoff = -6.393419870e-14
+ nfactor = -9.362812576e+00 lnfactor = 5.794310086e-06 wnfactor = 5.892821054e-06 pnfactor = -2.662853871e-12
+ eta0 = 8.774537750e-01 leta0 = -1.750829993e-07 weta0 = 3.380727087e-09 peta0 = -1.527686337e-15
+ etab = 3.496458977e-02 letab = -1.594104660e-08 wetab = -2.843472549e-17 petab = 1.284910958e-23
+ u0 = -3.066102449e-02 lu0 = 2.526450606e-08 wu0 = 2.308317452e-08 pu0 = -1.043084799e-14
+ ua = -7.671291415e-10 lua = -1.781110013e-16 wua = -1.661920357e-16 pua = 7.509902330e-23
+ ub = 3.598876228e-18 lub = -7.751685193e-25 wub = -8.863120791e-25 pub = 4.005075886e-31
+ uc = -7.895394521e-11 luc = 3.766779274e-17 wuc = 5.362290449e-18 puc = -2.423117170e-24
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.835515690e+05 lvsat = -2.635929281e-01 wvsat = -2.357605717e-01 pvsat = 1.065357229e-7
+ a0 = 1.500000005e+00 la0 = -2.213846884e-15 wa0 = -2.011759648e-15 pa0 = 9.090759256e-22
+ ags = -9.741017958e-01 lags = 4.490038944e-07 wags = -4.307366130e-16 pags = 1.946417680e-22
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.245981073e-05 lb0 = -5.473228192e-12 wb0 = -5.213256680e-12 pb0 = 2.355771642e-18
+ b1 = 1.908543627e-07 lb1 = -8.378432385e-14 wb1 = -7.976224276e-14 pb1 = 3.604304202e-20
+ keta = 2.272577853e-01 lketa = -1.034843988e-07 wketa = -7.194527992e-08 pketa = 3.251070503e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.954487361e-01 lpclm = 1.471855649e-07 wpclm = 2.796573233e-07 ppclm = -1.263718309e-13
+ pdiblc1 = 6.149252006e-01 lpdiblc1 = -5.207581960e-08 wpdiblc1 = 3.444089458e-16 ppdiblc1 = -1.556319518e-22
+ pdiblc2 = -4.393116250e-03 lpdiblc2 = 2.583921013e-09 wpdiblc2 = -9.234389295e-18 ppdiblc2 = 4.172845229e-24
+ pdiblcb = 3.822571344e-02 lpdiblcb = -2.857049862e-08 wpdiblcb = -2.734246163e-17 ppdiblcb = 1.235547081e-23
+ drout = 1.401075647e+00 ldrout = -1.812384643e-07 wdrout = -1.824133733e-15 pdrout = 8.242913019e-22
+ pscbe1 = 8.069286533e+08 lpscbe1 = -3.130926765e+00 wpscbe1 = -1.802082062e-07 ppscbe1 = 8.143305779e-14
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.398667074e-06 lalpha0 = -3.609024762e-13 walpha0 = -1.461114530e-13 palpha0 = 6.602498948e-20
+ alpha1 = 0.85
+ beta0 = 1.751788458e+01 lbeta0 = -8.666555999e-07 wbeta0 = -3.896305449e-07 pbeta0 = 1.760666402e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.371340241e-01 lkt1 = -7.622650712e-08 wkt1 = -9.740763608e-08 pkt1 = 4.401666000e-14
+ kt2 = -6.684223721e-02 lkt2 = 7.664068600e-09 wkt2 = -1.093058977e-17 pkt2 = 4.939340603e-24
+ at = 1.426051150e+05 lat = -6.444054199e-02 wat = -7.305572702e-02 pat = 3.301249498e-8
+ ute = -1.175988471e+00 lute = -1.394117633e-07 wute = -1.948152720e-07 pute = 8.803331991e-14
+ ua1 = 7.037062506e-10 lua1 = -1.468792469e-16 wua1 = -2.062421829e-24 pua1 = 9.319688865e-31
+ ub1 = -4.757344987e-19 lub1 = 2.389236723e-25 wub1 = -2.929768350e-33 pub1 = 1.323906777e-39
+ uc1 = 7.331997411e-11 luc1 = 1.491219767e-17 wuc1 = 4.242113053e-26 puc1 = -1.916929031e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.169 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.300065666e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -6.524727630e-07 wvth0 = -2.031575402e-06 pvth0 = 2.679261956e-13
+ k1 = 9.070734843e-01 lk1 = 7.553753179e-16 wk1 = 2.351978168e-15 pk1 = -3.101812140e-22
+ k2 = -5.981589482e-01 lk2 = 6.252886358e-08 wk2 = 1.946933395e-07 pk2 = -2.567635231e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -6.369845367e+00 ldsub = 9.223197130e-07 wdsub = 2.871785840e-06 pdsub = -3.787339884e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999948e-03 lcdscd = 6.857008017e-18 wcdscd = 2.135035898e-17 pcdscd = -2.815706869e-24
+ cit = 0.0
+ voff = {1.023017333e+00+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.622858129e-07 wvoff = -5.053021125e-07 pvoff = 6.663974790e-14
+ nfactor = 5.281986048e+01 lnfactor = -6.759190132e-06 wnfactor = -2.104578948e-05 pnfactor = 2.775539762e-12
+ eta0 = 2.940352071e-02 leta0 = -3.877765327e-09 weta0 = -1.207402531e-08 peta0 = 1.592334532e-15
+ etab = -4.399800025e-02 letab = 3.261524384e-17 wetab = 1.015525442e-16 petab = -1.339285627e-23
+ u0 = 2.256354792e-01 lu0 = -2.647688840e-08 wu0 = -8.243990900e-08 pu0 = 1.087225764e-14
+ ua = -2.593634727e-09 lua = 1.906257729e-16 wua = 5.935429848e-16 pua = -7.827704238e-23
+ ub = -5.276585960e-18 lub = 1.016618663e-24 wub = 3.165400282e-24 pub = -4.174561546e-31
+ uc = 1.380969564e-10 luc = -6.150660329e-18 wuc = -1.915103732e-17 puc = 2.525657952e-24
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.861646742e+06 lvsat = 2.704223521e-01 wvsat = 8.420020418e-01 pvsat = -1.110440713e-7
+ a0 = 1.499999983e+00 la0 = 2.307531943e-15 wa0 = 7.184858930e-15 pa0 = -9.475460416e-22
+ ags = 1.249999996e+00 lags = 4.940634568e-16 wags = 1.538342786e-15 pags = -2.028786028e-22
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -4.427135090e-05 lb0 = 5.979715451e-12 wb0 = 1.861877386e-11 pb0 = -2.455462515e-18
+ b1 = -6.773467057e-07 lb1 = 9.148897603e-14 wb1 = 2.848651527e-13 pb1 = -3.756830120e-20
+ keta = -6.941124947e-01 lketa = 8.252275465e-08 wketa = 2.569474283e-07 pketa = -3.388648379e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.613440115e+00 lpclm = -3.207728527e-07 wpclm = -9.987761546e-07 ppclm = 1.317195980e-13
+ pdiblc1 = 3.569721530e-01 lpdiblc1 = -3.950444416e-16 wpdiblc1 = -1.230032076e-15 ppdiblc1 = 1.622177948e-22
+ pdiblc2 = 8.406112020e-03 lpdiblc2 = 1.059204113e-17 wpdiblc2 = 3.297997986e-17 ppdiblc2 = -4.349430538e-24
+ pdiblcb = -1.032957702e-01 lpdiblcb = 3.136224613e-17 wpdiblcb = 9.765144249e-17 ppdiblcb = -1.287833729e-23
+ drout = 5.033266441e-01 ldrout = 2.092319651e-15 wdrout = 6.514763840e-15 pdrout = -8.591736211e-22
+ pscbe1 = 7.914198784e+08 lpscbe1 = 2.067041397e-07 wpscbe1 = 6.436042786e-07 ppscbe1 = -8.487915993e-14
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.219188974e-06 lalpha0 = 1.675929206e-13 walpha0 = 5.218266178e-13 palpha0 = -6.881901618e-20
+ alpha1 = 0.85
+ beta0 = 1.101122937e+01 lbeta0 = 4.469144591e-07 wbeta0 = 1.391537660e-06 pbeta0 = -1.835173782e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.068153396e+00 lkt1 = 1.117286146e-07 wkt1 = 3.478844146e-07 pkt1 = -4.587934448e-14
+ kt2 = -2.887893910e-02 lkt2 = 1.253763759e-17 wkt2 = 3.903788404e-17 pkt2 = -5.148353965e-24
+ at = -5.916740043e+05 lat = 8.379646091e-02 wat = 2.609133108e-01 pat = -3.440950834e-8
+ ute = -2.973428510e+00 lute = 2.234572290e-07 wute = 6.957688284e-07 pute = -9.175868886e-14
+ ua1 = -2.384735394e-11 lua1 = 2.365640573e-24 wua1 = 7.365789721e-24 pua1 = -9.714077143e-31
+ ub1 = 7.077531445e-19 lub1 = 3.360506627e-33 wub1 = 1.046345875e-32 pub1 = -1.379931501e-39
+ uc1 = 1.471862504e-10 luc1 = -4.865786556e-26 wuc1 = -1.515039195e-25 puc1 = 1.998044430e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.170 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {-3.035229047e+00+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.467942390e-07 wvth0 = 1.604969324e-06 pvth0 = -2.116649594e-13
+ k1 = 0.90707349
+ k2 = -1.512266114e+00 lk2 = 1.830822307e-07 wk2 = 5.861840111e-07 pk2 = -7.730653357e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 3.213159080e+00 ldsub = -3.414964965e-07 wdsub = -1.140985314e-06 pdsub = 1.504742842e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = -6.688470453e+00 lnfactor = 1.088828059e-06 wnfactor = 1.671005367e-06 pnfactor = -2.203738588e-13
+ eta0 = 5.391586575e-04 leta0 = -7.110477581e-11 weta0 = -2.375705338e-10 peta0 = 3.133103957e-17
+ etab = -0.043998
+ u0 = 1.737752934e-01 lu0 = -1.963751524e-08 wu0 = -7.101431164e-08 pu0 = 9.365438434e-15
+ ua = -2.844196309e-09 lua = 2.236700849e-16 wua = 7.848996634e-16 pua = -1.035133525e-22
+ ub = 1.292471857e-17 lub = -1.383787580e-24 wub = -5.386702958e-24 pub = 7.104037728e-31
+ uc = -1.316563759e-10 luc = 2.942467889e-17 wuc = 1.330372550e-16 puc = -1.754508622e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.079825513e+05 lvsat = -5.527482872e-02 wvsat = -1.054266865e-01 pvsat = 1.390377685e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.001055089e-06 lb0 = 8.007095686e-13 wb0 = 4.651170118e-12 pb0 = -6.134009663e-19
+ b1 = 8.433993044e-08 lb1 = -8.963019229e-15 wb1 = -3.961488857e-14 pb1 = 5.224451119e-21
+ keta = -9.616951609e-01 lketa = 1.178118243e-07 wketa = 4.295745452e-07 pketa = -5.665272059e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.592040983e-02 lpclm = 2.179064358e-08 wpclm = 1.287409127e-07 ppclm = -1.697848030e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.249543125e-07 lalpha0 = -9.674040084e-15 walpha0 = 3.315074562e-21 palpha0 = -4.371953410e-28
+ alpha1 = 0.85
+ beta0 = 1.626781828e+01 lbeta0 = -2.463297428e-07 wbeta0 = 2.293410262e-14 pbeta0 = -3.024567263e-21
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.530400707e-01 lkt1 = -8.957445783e-09 wkt1 = -1.142115735e-15 pkt1 = 1.506234026e-22
+ kt2 = -0.028878939
+ at = 9.760154499e+03 lat = 4.478722611e-03 wat = -3.668076824e-10 pat = 4.837499000e-17
+ ute = -9.181979405e-01 lute = -4.758863367e-08 wute = -2.487840260e-07 pute = 3.280988613e-14
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.171 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {0.4913699+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56800772
+ k2 = -0.040590746
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.10827784+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 2.78042
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.025731
+ ua = -1.0529435e-9
+ ub = 1.832e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 9.1484e-8
+ b1 = 1.6098e-9
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.172 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.817702567e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.915309403e-7
+ k1 = 5.567098995e-01 lk1 = 2.254127697e-7
+ k2 = -3.378657655e-02 lk2 = -1.357559791e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.017808550e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.296270710e-7
+ nfactor = 2.803162380e+00 lnfactor = -4.537532526e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.477246701e-02 lu0 = 1.912453613e-8
+ ua = -1.141749888e-09 lua = 1.771854492e-15
+ ub = 1.874174789e-18 lub = -8.414663684e-25
+ uc = 6.327183549e-11 luc = -2.939876843e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.478299869e+00 la0 = -2.308430009e-6
+ ags = 3.215147230e-01 lags = 4.661812263e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 7.827327503e-08 lb0 = 2.635788125e-13
+ b1 = 1.664204119e-09 lb1 = -1.085464512e-15
+ keta = -1.976419529e-03 lketa = -5.127993490e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.729504833e-02 lpclm = 8.812755480e-07 ppclm = -2.220446049e-28
+ pdiblc1 = 0.39
+ pdiblc2 = -1.515165620e-04 lpdiblc2 = 2.218337962e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -6.522518163e+07 lpscbe1 = 5.790538287e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.785341441e-01 lkt1 = -1.565395837e-7
+ kt2 = -2.847160196e-02 lkt2 = -2.087623258e-8
+ at = 1.882531350e+05 lat = -2.644249724e-1
+ ute = -1.123882006e+00 lute = 1.692319823e-7
+ ua1 = 8.774736444e-10 lua1 = 4.858808868e-15
+ ub1 = -2.494531757e-19 lub1 = -6.384937596e-24
+ uc1 = 4.313166665e-11 luc1 = -1.858179462e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.173 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.174172339e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -9.192958009e-8
+ k1 = 6.071532016e-01 lk1 = -1.757063659e-7
+ k2 = -6.227740302e-02 lk2 = 9.079968255e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.259465233e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 6.253544744e-8
+ nfactor = 2.290448121e+00 lnfactor = 3.623289522e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.588029506e-02 lu0 = 1.031521930e-8
+ ua = -1.229966275e-09 lua = 2.473340703e-15
+ ub = 2.072832611e-18 lub = -2.421169734e-24
+ uc = 3.252620055e-11 luc = -4.950205394e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.205783465e+00 la0 = -1.414119935e-7
+ ags = 4.064200086e-01 lags = -2.089755015e-07 wags = -4.440892099e-22
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.235987093e-07 lb0 = -9.684364686e-14
+ b1 = 1.691406670e-09 lb1 = -1.301775962e-15
+ keta = -1.917560068e-02 lketa = 8.548590692e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.426882576e-01 lpclm = 3.389244816e-06 wpclm = 1.110223025e-22 ppclm = 8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = -1.025171335e-03 lpdiblc2 = 2.913057840e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 5.275926511e+08 lpscbe1 = 1.076521426e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.828274235e-01 lkt1 = -1.223999366e-7
+ kt2 = -1.864692104e-02 lkt2 = -9.900092610e-8
+ at = 1.698195537e+05 lat = -1.178433279e-1
+ ute = -8.085800536e-01 lute = -2.338011625e-6
+ ua1 = 2.387533168e-09 lua1 = -7.149004768e-15
+ ub1 = -1.684552764e-18 lub1 = 5.026803557e-24
+ uc1 = -1.180400046e-11 luc1 = 2.510239413e-16 puc1 = 1.033975766e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.174 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {5.036991516e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.771735122e-8
+ k1 = 5.224894914e-01 lk1 = 1.588745419e-7
+ k2 = -2.026099817e-02 lk2 = -7.524414950e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.115687121e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 5.716048642e-9
+ nfactor = 2.758367370e+00 lnfactor = 1.774128331e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.831834410e-02 lu0 = 6.803396468e-10
+ ua = -4.918389228e-10 lua = -4.436507565e-16
+ ub = 1.373220533e-18 lub = 3.436139465e-25
+ uc = -4.842565427e-12 luc = 9.817486230e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.363604600e+04 lvsat = 2.622624489e-1
+ a0 = 8.479396350e-01 la0 = 1.272744237e-6
+ ags = 4.366510930e-01 lags = -3.284451492e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 7.325302338e-08 lb0 = 1.021165126e-13
+ b1 = -1.246317312e-08 lb1 = 5.463543899e-14 wb1 = 3.308722450e-30 pb1 = -1.654361225e-35
+ keta = -1.264073531e-02 lketa = 5.966089661e-08 pketa = -6.938893904e-30
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.366646536e-01 lpclm = 4.946192650e-06 ppclm = 1.776356839e-27
+ pdiblc1 = 0.39
+ pdiblc2 = -5.529034283e-04 lpdiblc2 = 2.726423184e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.057875285e-01 lkt1 = -3.166433390e-8
+ kt2 = -5.663636600e-02 lkt2 = 5.112883963e-8
+ at = 140000.0
+ ute = -1.610417584e+00 lute = 8.307548749e-07 wute = -1.776356839e-21
+ ua1 = -3.141532565e-10 lua1 = 3.527738482e-15
+ ub1 = 5.536467273e-20 lub1 = -1.849143105e-24
+ uc1 = 5.805098873e-11 luc1 = -2.503466317e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.175 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-09*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.777096706e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.301102283e-8
+ k1 = 6.212681700e-01 lk1 = -3.392968399e-8
+ k2 = -6.384985590e-02 lk2 = 9.836113722e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.455643000e-01 ldsub = -5.573875314e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-9.823954033e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.030090856e-8
+ nfactor = 3.309041785e+00 lnfactor = 6.992774020e-7
+ eta0 = 1.537410312e-01 leta0 = -1.439337178e-7
+ etab = -1.363342072e-01 letab = 1.294764787e-7
+ u0 = 3.243815733e-02 lu0 = -7.361045536e-9
+ ua = -2.385002539e-10 lua = -9.381376908e-16
+ ub = 1.185339856e-18 lub = 7.103346701e-25
+ uc = 4.822878123e-11 luc = -5.414090889e-18 wuc = -5.169878828e-32
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.213473320e+05 lvsat = 5.202283627e-2
+ a0 = 1.5
+ ags = 3.313088529e-01 lags = -1.228296323e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.127983295e-07 lb0 = -3.654474191e-13
+ b1 = 2.106042756e-08 lb1 = -1.079864024e-14
+ keta = 1.805004733e-02 lketa = -2.438589030e-10
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.522733322e+00 lpclm = -1.415764330e-6
+ pdiblc1 = 2.001896837e-01 lpdiblc1 = 3.704871499e-7
+ pdiblc2 = 2.062764645e-02 lpdiblc2 = -1.407768104e-8
+ pdiblcb = -0.025
+ drout = 4.703102312e-01 ldrout = 1.750637556e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.467909273e-01 lkt1 = 4.836942111e-8
+ kt2 = -3.423300662e-02 lkt2 = 7.400148129e-9
+ at = 1.495188100e+05 lat = -1.857958438e-2
+ ute = -1.628064281e+00 lute = 8.651991289e-7
+ ua1 = 8.257868283e-10 lua1 = 1.302711089e-15
+ ub1 = -4.438155885e-19 lub1 = -8.748026374e-25
+ uc1 = 4.300065746e-11 luc1 = 4.341792472e-18
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.176 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {4.768969173e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.378466728e-8
+ k1 = 5.947741785e-01 lk1 = -8.710556888e-9
+ k2 = -5.950168308e-02 lk2 = 5.697170628e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.191289451e-01 ldsub = 3.890438058e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.073244113e-01+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.165319250e-8
+ nfactor = 4.571316858e+00 lnfactor = -5.022582567e-7
+ eta0 = -4.380244824e-01 leta0 = 4.193566311e-07 weta0 = 1.665334537e-22 peta0 = 1.734723476e-29
+ etab = -0.0003125
+ u0 = 2.421369690e-02 lu0 = 4.676620846e-10 wu0 = -2.775557562e-23
+ ua = -1.280798932e-09 lua = 5.400661752e-17
+ ub = 1.975083776e-18 lub = -4.140756249e-26
+ uc = 7.700792919e-11 luc = -3.280841503e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.541038350e+05 lvsat = 2.084254342e-2
+ a0 = 1.5
+ ags = 3.674223382e-01 lags = -1.572053728e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -4.496483497e-07 lb0 = 3.603110884e-13 pb0 = -5.293955920e-35
+ b1 = 1.357848841e-08 lb1 = -3.676724520e-15
+ keta = 3.545712353e-02 lketa = -1.681332400e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.409768704e+00 lpclm = -3.563544566e-7
+ pdiblc1 = 6.704934226e-01 lpdiblc1 = -7.718604331e-8
+ pdiblc2 = 9.917256884e-03 lpdiblc2 = -3.882664709e-9
+ pdiblcb = -0.025
+ drout = 3.417242576e-01 ldrout = 2.974623007e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -4.851443400e-07 lalpha0 = 4.903561095e-13 walpha0 = 1.058791184e-28 palpha0 = -2.117582368e-34
+ alpha1 = 0.85
+ beta0 = 1.228745412e+01 lbeta0 = 1.496876545e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.870790129e-01 lkt1 = -8.469215655e-9
+ kt2 = -5.289864105e-03 lkt2 = -2.015027931e-8
+ at = 2.474890600e+05 lat = -1.118356039e-1
+ ute = -2.741143519e-02 lute = -6.584319030e-7
+ ua1 = 3.835299287e-09 lua1 = -1.561986640e-15
+ ub1 = -2.642421110e-18 lub1 = 1.218008185e-24
+ uc1 = -5.541599185e-12 luc1 = 5.054824427e-17 puc1 = -2.584939414e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.177 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {6.323841045e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -5.647703838e-8
+ k1 = 3.077427617e-01 lk1 = 1.209934868e-7
+ k2 = 1.539354899e-02 lk2 = -2.814656173e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.802140521e-02 ldsub = 1.162246268e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.103590352e-03 lcdscd = -1.221701112e-9
+ cit = 0.0
+ voff = {-7.301876348e-02+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.715526294e-8
+ nfactor = 4.987800757e+00 lnfactor = -6.904594174e-7
+ eta0 = 8.856867600e-01 leta0 = -1.788033288e-7
+ etab = 3.496458970e-02 letab = -1.594104657e-08 wetab = -4.336808690e-25
+ u0 = 2.555274969e-02 lu0 = -1.374304279e-10
+ ua = -1.171851705e-09 lua = 4.775435517e-18
+ ub = 1.440466559e-18 lub = 2.001758002e-25
+ uc = -6.589531741e-11 luc = 3.176684695e-17 wuc = -6.462348536e-33 puc = -6.462348536e-39
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.094108014e+05 lvsat = -4.149623866e-3
+ a0 = 1.5
+ ags = -9.741017969e-01 lags = 4.490038949e-07 wags = -3.885780586e-22 pags = -9.714451465e-29
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -2.358795196e-07 lb0 = 2.637130157e-13
+ b1 = -3.388274940e-09 lb1 = 3.990233470e-15
+ keta = 5.205156677e-02 lketa = -2.431203761e-08 wketa = 1.734723476e-23 pketa = 3.035766083e-30
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 9.764899684e-01 lpclm = -1.605640282e-7
+ pdiblc1 = 6.149252015e-01 lpdiblc1 = -5.207581998e-8
+ pdiblc2 = -4.393116272e-03 lpdiblc2 = 2.583921023e-09 ppdiblc2 = -4.336808690e-31
+ pdiblcb = 3.822571337e-02 lpdiblcb = -2.857049858e-8
+ drout = 1.401075642e+00 ldrout = -1.812384623e-7
+ pscbe1 = 8.069286528e+08 lpscbe1 = -3.130926566e+0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.042846162e-06 lalpha0 = -2.001137663e-13
+ alpha1 = 0.85
+ beta0 = 1.656902880e+01 lbeta0 = -4.378857032e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.743479677e-01 lkt1 = 3.096596692e-8
+ kt2 = -6.684223724e-02 lkt2 = 7.664068612e-9
+ at = -3.530534254e+04 lat = 1.595381349e-2
+ ute = -1.650416358e+00 lute = 7.497318452e-8
+ ua1 = 7.037062456e-10 lua1 = -1.468792446e-16
+ ub1 = -4.757345058e-19 lub1 = 2.389236755e-25 wub1 = 9.629649722e-41 pub1 = 3.611118646e-47
+ uc1 = 7.331997422e-11 luc1 = 1.491219762e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.178 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {0.35263+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.90707349
+ k2 = -0.124028
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.62373
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = 1.56767
+ eta0 = 0.0
+ etab = -0.043998
+ u0 = 0.024872
+ ua = -1.148197e-9
+ ub = 2.43202e-18
+ uc = 9.1459e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 188856.0
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.0704e-6
+ b1 = 1.6377e-8
+ keta = -0.068376
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.18115
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 5.16e-8
+ alpha1 = 0.85
+ beta0 = 14.4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.22096074
+ kt2 = -0.028878939
+ at = 43720.487
+ ute = -1.2790432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8__model.179 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {3.932304e-09+sky130_fd_pr__nfet_01v8__toxe_slope_spectre*(4.148e-9*0.948*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = -1.0316e-8
+ lint = 2.40595e-8
+ vth0 = {-3.045170427e-01+sky130_fd_pr__nfet_01v8__vth0_slope_spectre*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.666520914e-08 wvth0 = 4.836515918e-07 pvth0 = -6.378445558e-14
+ k1 = 0.90707349
+ k2 = -4.744370369e-01 lk2 = 4.621229419e-08 wk2 = 1.600181815e-07 pk2 = -2.110335779e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 3.290138835e+00 ldsub = -3.516486635e-07 wdsub = -1.172595665e-06 pdsub = 1.546430889e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {-0.20753+sky130_fd_pr__nfet_01v8__voff_slope_spectre*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = -6.688470389e+00 lnfactor = 1.088828051e-06 wnfactor = 1.671005340e-06 pnfactor = -2.203738553e-13
+ eta0 = 8.627946104e-04 leta0 = -1.137862046e-10 weta0 = -3.704657991e-10 peta0 = 4.885740006e-17
+ etab = -0.043998
+ u0 = 7.747248961e-02 lu0 = -6.937005170e-09 wu0 = -3.146929871e-08 pu0 = 4.150202584e-15
+ ua = -2.844194477e-09 lua = 2.236698432e-16 wua = 7.848989109e-16 pua = -1.035132533e-22
+ ub = 1.292468824e-17 lub = -1.383783580e-24 wub = -5.386690503e-24 pub = 7.104021303e-31
+ uc = -1.406321093e-10 luc = 3.060840758e-17 wuc = 1.367229783e-16 puc = -1.803116311e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.059330551e+05 lvsat = -1.544023911e-02 wvsat = 1.860450219e-02 pvsat = -2.453580354e-9
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.001032725e-06 lb0 = 8.007066192e-13 wb0 = 4.651160935e-12 pb0 = -6.133997552e-19
+ b1 = 8.433660613e-08 lb1 = -8.962580816e-15 wb1 = -3.961352350e-14 pb1 = 5.224271092e-21
+ keta = -9.616948578e-01 lketa = 1.178117843e-07 wketa = 4.295744207e-07 pketa = -5.665270418e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.592022520e-02 lpclm = 2.179066793e-08 wpclm = 1.287409885e-07 ppclm = -1.697849030e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.249543199e-07 lalpha0 = -9.674041067e-15 walpha0 = 2.526371056e-22 palpha0 = -3.331806745e-29
+ alpha1 = 0.85
+ beta0 = 1.626781834e+01 lbeta0 = -2.463297501e-07 wbeta0 = 4.422417987e-17 pbeta0 = -5.826450433e-24
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 2.3267e-8
+ dwc = -3.2175e-8
+ xpart = 0.0
+ cgso = 2.4083264e-10
+ cgdo = 2.4083264e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.00104159201
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 2.856175336e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 1.852257592e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.530400733e-01 lkt1 = -8.957445446e-09 wkt1 = -9.402256751e-17 pkt1 = 1.239974790e-23
+ kt2 = -0.028878939
+ at = 9.760153678e+03 lat = 4.478722719e-03 wat = -2.983096056e-11 pat = 3.934124834e-18
+ ute = -9.014130388e-01 lute = -4.980224329e-08 wute = -2.556764437e-07 pute = 3.371886508e-14
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
.ends sky130_fd_pr__nfet_01v8
* Well Proximity Effect Parameters
