magic
tech sky130A
magscale 1 2
timestamp 1624884095
<< checkpaint >>
rect -1738 -1738 7260 8260
use sky130_fd_pr__genrivetdlring__example_559591418082  sky130_fd_pr__genrivetdlring__example_559591418082_0
timestamp 1624884095
transform 1 0 -478 0 1 -478
box 0 0 1 1
use sky130_fd_pr__gendlring__example_559591418081  sky130_fd_pr__gendlring__example_559591418081_0
timestamp 1624884095
transform 1 0 0 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 6000 6666 6000 6666 0 FreeSans 2000 0 0 0 HP
flabel comment s 6000 7000 6000 7000 0 FreeSans 2000 0 0 0 PLASTIC
flabel comment s 6000 7000 6000 7000 0 FreeSans 2000 0 0 0 PLASTIC
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 3925468
string GDS_START 3924600
<< end >>
