magic
tech sky130A
magscale 1 2
timestamp 1624884095
<< checkpaint >>
rect -1629 -2052 9937 4599
<< nwell >>
rect 1693 1097 4305 1263
rect 2517 555 2565 1097
rect 6085 979 6965 1730
<< mvnsubdiff >>
rect 1759 1163 1783 1197
rect 1817 1163 1852 1197
rect 1886 1163 1921 1197
rect 1955 1163 1990 1197
rect 2024 1163 2059 1197
rect 2093 1163 2128 1197
rect 2162 1163 2197 1197
rect 2231 1163 2266 1197
rect 2300 1163 2335 1197
rect 2369 1163 2404 1197
rect 2438 1163 2473 1197
rect 2507 1163 2542 1197
rect 2576 1163 2611 1197
rect 2645 1163 2680 1197
rect 2714 1163 2749 1197
rect 2783 1163 2818 1197
rect 2852 1163 2887 1197
rect 2921 1163 2956 1197
rect 2990 1163 3025 1197
rect 3059 1163 3093 1197
rect 3127 1163 3161 1197
rect 3195 1163 3229 1197
rect 3263 1163 3297 1197
rect 3331 1163 3365 1197
rect 3399 1163 3433 1197
rect 3467 1163 3501 1197
rect 3535 1163 3569 1197
rect 3603 1163 3637 1197
rect 3671 1163 3705 1197
rect 3739 1163 3773 1197
rect 3807 1163 3841 1197
rect 3875 1163 3909 1197
rect 3943 1163 3977 1197
rect 4011 1163 4045 1197
rect 4079 1163 4113 1197
rect 4147 1163 4181 1197
rect 4215 1163 4239 1197
<< mvnsubdiffcont >>
rect 1783 1163 1817 1197
rect 1852 1163 1886 1197
rect 1921 1163 1955 1197
rect 1990 1163 2024 1197
rect 2059 1163 2093 1197
rect 2128 1163 2162 1197
rect 2197 1163 2231 1197
rect 2266 1163 2300 1197
rect 2335 1163 2369 1197
rect 2404 1163 2438 1197
rect 2473 1163 2507 1197
rect 2542 1163 2576 1197
rect 2611 1163 2645 1197
rect 2680 1163 2714 1197
rect 2749 1163 2783 1197
rect 2818 1163 2852 1197
rect 2887 1163 2921 1197
rect 2956 1163 2990 1197
rect 3025 1163 3059 1197
rect 3093 1163 3127 1197
rect 3161 1163 3195 1197
rect 3229 1163 3263 1197
rect 3297 1163 3331 1197
rect 3365 1163 3399 1197
rect 3433 1163 3467 1197
rect 3501 1163 3535 1197
rect 3569 1163 3603 1197
rect 3637 1163 3671 1197
rect 3705 1163 3739 1197
rect 3773 1163 3807 1197
rect 3841 1163 3875 1197
rect 3909 1163 3943 1197
rect 3977 1163 4011 1197
rect 4045 1163 4079 1197
rect 4113 1163 4147 1197
rect 4181 1163 4215 1197
<< locali >>
rect 4876 3017 4982 3076
rect 4910 2983 4948 3017
rect 4876 2942 4982 2983
rect 5038 3013 5144 3074
rect 5072 2979 5110 3013
rect 5038 2940 5144 2979
rect 5213 3012 5319 3074
rect 5247 2978 5285 3012
rect 5213 2940 5319 2978
rect 6141 3003 6175 3041
rect 6287 3003 6321 3041
rect 6441 3003 6475 3041
rect 3394 2635 3454 2671
rect 2461 2570 2499 2604
rect 894 2527 928 2565
rect 2726 2495 2760 2538
rect 2843 2522 2877 2560
rect 3769 2491 3807 2525
rect 469 2342 507 2376
rect 663 2332 713 2428
rect 760 2375 803 2409
rect 1228 2396 1234 2430
rect 997 2360 1014 2378
rect 1048 2378 1054 2394
rect 1048 2360 1063 2378
rect 1342 2358 1380 2392
rect 1479 2373 1513 2413
rect 1583 2372 1617 2412
rect 1764 2396 1802 2430
rect 2009 2374 2043 2400
rect 2294 2399 2299 2433
rect 2481 2399 2490 2433
rect 2009 2359 2053 2374
rect 2588 2365 2626 2399
rect 3016 2365 3050 2404
rect 3131 2426 3165 2438
rect 2043 2325 2053 2359
rect 3215 2365 3249 2404
rect 3308 2418 3342 2428
rect 3516 2356 3550 2394
rect 3735 2332 3792 2428
rect 4082 2424 4116 2439
rect 4260 2424 4294 2439
rect 4396 2394 4434 2428
rect 3941 2340 3979 2374
rect 1103 2208 1137 2246
rect 4175 2229 4209 2267
rect 4550 2285 4584 2323
rect 1282 1969 1342 2005
rect 3394 1969 3454 2075
rect 951 1755 1039 1952
rect 1907 1767 1947 1801
rect 951 1746 989 1755
rect 986 1721 989 1746
rect 1023 1721 1039 1755
rect 906 1711 940 1712
rect 986 1683 1039 1721
rect 755 1622 768 1656
rect 986 1649 989 1683
rect 1023 1649 1039 1683
rect 1489 1690 1523 1728
rect 1387 1660 1421 1673
rect 986 1616 1039 1649
rect 1589 1690 1623 1700
rect 1873 1616 1927 1767
rect 2734 1725 2768 1763
rect 3041 1746 3151 1952
rect 3509 1861 3543 1899
rect 2009 1667 2047 1701
rect 2133 1637 2167 1675
rect 1190 1578 1224 1616
rect 2199 1616 2249 1712
rect 2433 1698 2467 1708
rect 2587 1667 2625 1701
rect 2997 1662 3031 1710
rect 2868 1622 2881 1656
rect 3098 1660 3151 1746
rect 3792 1861 3826 1899
rect 3307 1756 3341 1794
rect 3098 1626 3117 1660
rect 3151 1626 3189 1660
rect 3098 1616 3151 1626
rect 3729 1616 3791 1712
rect 3937 1651 3975 1685
rect 1660 1450 1705 1484
rect 1282 1373 1342 1409
rect 3394 1373 3454 1409
rect 1759 1163 1774 1197
rect 1817 1163 1847 1197
rect 1886 1163 1920 1197
rect 1955 1163 1990 1197
rect 2027 1163 2059 1197
rect 2100 1163 2128 1197
rect 2173 1163 2197 1197
rect 2246 1163 2266 1197
rect 2319 1163 2335 1197
rect 2392 1163 2404 1197
rect 2465 1163 2473 1197
rect 2538 1163 2542 1197
rect 2576 1163 2577 1197
rect 2645 1163 2650 1197
rect 2714 1163 2723 1197
rect 2783 1163 2796 1197
rect 2852 1163 2869 1197
rect 2921 1163 2942 1197
rect 2990 1163 3015 1197
rect 3059 1163 3088 1197
rect 3127 1163 3161 1197
rect 3195 1163 3229 1197
rect 3268 1163 3297 1197
rect 3341 1163 3365 1197
rect 3414 1163 3433 1197
rect 3487 1163 3501 1197
rect 3560 1163 3569 1197
rect 3632 1163 3637 1197
rect 3704 1163 3705 1197
rect 3739 1163 3742 1197
rect 3807 1163 3814 1197
rect 3875 1163 3886 1197
rect 3943 1163 3958 1197
rect 4011 1163 4030 1197
rect 4079 1163 4102 1197
rect 4147 1163 4181 1197
rect 4215 1163 4239 1197
rect 3180 918 3218 952
rect 2777 875 2791 909
rect 2825 875 2843 909
rect 2777 837 2843 875
rect 1888 802 1926 836
rect 2605 786 2625 820
rect 2659 786 2672 820
rect 1963 684 1979 718
rect 2013 684 2029 718
rect 1963 646 2029 684
rect 1963 612 1979 646
rect 2013 612 2029 646
rect 1963 573 2029 612
rect 2145 684 2162 718
rect 2196 684 2211 718
rect 2145 646 2211 684
rect 2246 690 2280 728
rect 2605 748 2672 786
rect 2605 714 2625 748
rect 2659 714 2672 748
rect 2145 612 2162 646
rect 2196 612 2211 646
rect 2145 573 2211 612
rect 2316 573 2333 582
rect 1802 501 1836 539
rect 2367 573 2382 582
rect 2333 510 2367 548
rect 2605 471 2672 714
rect 2777 803 2791 837
rect 2825 803 2843 837
rect 2777 573 2843 803
rect 3242 764 3264 798
rect 3298 764 3308 798
rect 3242 726 3308 764
rect 3242 692 3264 726
rect 3298 692 3308 726
rect 3105 573 3137 598
rect 3242 573 3308 692
rect 3748 622 3786 656
rect 3936 652 3970 690
rect 3537 573 3554 598
rect 3071 526 3105 564
rect 3588 573 3603 598
rect 3554 526 3588 564
rect 3741 498 3775 536
rect 2708 452 2742 490
rect 4030 493 4064 531
rect 4197 511 4231 549
rect 4536 513 4682 1246
rect 7815 1114 8309 1126
rect 4787 1080 4825 1114
rect 7849 1080 7887 1114
rect 7921 1080 8309 1114
rect 7815 1074 8309 1080
rect 7815 959 8309 971
rect 4787 925 4825 959
rect 7849 925 7887 959
rect 7921 925 8309 959
rect 7815 917 8309 925
rect 7815 809 8309 815
rect 4787 775 4825 809
rect 7844 775 7882 809
rect 7916 775 8309 809
rect 7815 767 8309 775
rect 7815 653 8309 659
rect 4787 619 4825 653
rect 7815 619 7816 653
rect 7850 619 7888 653
rect 7922 619 8309 653
rect 7815 612 8309 619
rect 4536 460 4882 513
<< viali >>
rect 4876 2983 4910 3017
rect 4948 2983 4982 3017
rect 5038 2979 5072 3013
rect 5110 2979 5144 3013
rect 5213 2978 5247 3012
rect 5285 2978 5319 3012
rect 6141 3041 6175 3075
rect 6141 2969 6175 3003
rect 6287 3041 6321 3075
rect 6287 2969 6321 3003
rect 6441 3041 6475 3075
rect 6441 2969 6475 3003
rect 894 2565 928 2599
rect 2427 2570 2461 2604
rect 2499 2570 2533 2604
rect 894 2493 928 2527
rect 2726 2538 2760 2572
rect 2726 2461 2760 2495
rect 2843 2560 2877 2594
rect 2843 2488 2877 2522
rect 3735 2491 3769 2525
rect 3807 2491 3841 2525
rect 435 2342 469 2376
rect 507 2342 541 2376
rect 726 2375 760 2409
rect 803 2375 837 2409
rect 1194 2396 1228 2430
rect 1479 2413 1513 2447
rect 1014 2360 1048 2394
rect 1308 2358 1342 2392
rect 1380 2358 1414 2392
rect 1479 2339 1513 2373
rect 1583 2412 1617 2446
rect 1730 2396 1764 2430
rect 1802 2396 1836 2430
rect 2009 2400 2043 2434
rect 1583 2338 1617 2372
rect 2260 2399 2294 2433
rect 2447 2399 2481 2433
rect 3016 2404 3050 2438
rect 2554 2365 2588 2399
rect 2626 2365 2660 2399
rect 3131 2392 3165 2426
rect 3215 2404 3249 2438
rect 2009 2325 2043 2359
rect 3016 2331 3050 2365
rect 3308 2384 3342 2418
rect 3516 2394 3550 2428
rect 3215 2331 3249 2365
rect 3516 2322 3550 2356
rect 4082 2390 4116 2424
rect 4260 2390 4294 2424
rect 4362 2394 4396 2428
rect 4434 2394 4468 2428
rect 3907 2340 3941 2374
rect 3979 2340 4013 2374
rect 4550 2323 4584 2357
rect 1103 2246 1137 2280
rect 1103 2174 1137 2208
rect 4175 2267 4209 2301
rect 4550 2251 4584 2285
rect 4175 2195 4209 2229
rect 1873 1767 1907 1801
rect 1947 1767 1981 1801
rect 989 1721 1023 1755
rect 906 1677 940 1711
rect 721 1622 755 1656
rect 989 1649 1023 1683
rect 1489 1728 1523 1762
rect 1190 1616 1224 1650
rect 1387 1626 1421 1660
rect 1489 1656 1523 1690
rect 1589 1656 1623 1690
rect 2734 1763 2768 1797
rect 3509 1899 3543 1933
rect 1975 1667 2009 1701
rect 2047 1667 2081 1701
rect 2133 1675 2167 1709
rect 2133 1603 2167 1637
rect 2433 1664 2467 1698
rect 2553 1667 2587 1701
rect 2625 1667 2659 1701
rect 2734 1691 2768 1725
rect 2834 1622 2868 1656
rect 2997 1628 3031 1662
rect 3307 1794 3341 1828
rect 3509 1827 3543 1861
rect 3792 1899 3826 1933
rect 3792 1827 3826 1861
rect 3307 1722 3341 1756
rect 3117 1626 3151 1660
rect 3189 1626 3223 1660
rect 3903 1651 3937 1685
rect 3975 1651 4009 1685
rect 1190 1544 1224 1578
rect 1705 1450 1739 1484
rect 1774 1163 1783 1197
rect 1783 1163 1808 1197
rect 1847 1163 1852 1197
rect 1852 1163 1881 1197
rect 1920 1163 1921 1197
rect 1921 1163 1954 1197
rect 1993 1163 2024 1197
rect 2024 1163 2027 1197
rect 2066 1163 2093 1197
rect 2093 1163 2100 1197
rect 2139 1163 2162 1197
rect 2162 1163 2173 1197
rect 2212 1163 2231 1197
rect 2231 1163 2246 1197
rect 2285 1163 2300 1197
rect 2300 1163 2319 1197
rect 2358 1163 2369 1197
rect 2369 1163 2392 1197
rect 2431 1163 2438 1197
rect 2438 1163 2465 1197
rect 2504 1163 2507 1197
rect 2507 1163 2538 1197
rect 2577 1163 2611 1197
rect 2650 1163 2680 1197
rect 2680 1163 2684 1197
rect 2723 1163 2749 1197
rect 2749 1163 2757 1197
rect 2796 1163 2818 1197
rect 2818 1163 2830 1197
rect 2869 1163 2887 1197
rect 2887 1163 2903 1197
rect 2942 1163 2956 1197
rect 2956 1163 2976 1197
rect 3015 1163 3025 1197
rect 3025 1163 3049 1197
rect 3088 1163 3093 1197
rect 3093 1163 3122 1197
rect 3161 1163 3195 1197
rect 3234 1163 3263 1197
rect 3263 1163 3268 1197
rect 3307 1163 3331 1197
rect 3331 1163 3341 1197
rect 3380 1163 3399 1197
rect 3399 1163 3414 1197
rect 3453 1163 3467 1197
rect 3467 1163 3487 1197
rect 3526 1163 3535 1197
rect 3535 1163 3560 1197
rect 3598 1163 3603 1197
rect 3603 1163 3632 1197
rect 3670 1163 3671 1197
rect 3671 1163 3704 1197
rect 3742 1163 3773 1197
rect 3773 1163 3776 1197
rect 3814 1163 3841 1197
rect 3841 1163 3848 1197
rect 3886 1163 3909 1197
rect 3909 1163 3920 1197
rect 3958 1163 3977 1197
rect 3977 1163 3992 1197
rect 4030 1163 4045 1197
rect 4045 1163 4064 1197
rect 4102 1163 4113 1197
rect 4113 1163 4136 1197
rect 3146 918 3180 952
rect 3218 918 3252 952
rect 2791 875 2825 909
rect 1854 802 1888 836
rect 1926 802 1960 836
rect 2625 786 2659 820
rect 2246 728 2280 762
rect 1979 684 2013 718
rect 1979 612 2013 646
rect 2162 684 2196 718
rect 2246 656 2280 690
rect 2625 714 2659 748
rect 2162 612 2196 646
rect 1802 539 1836 573
rect 1802 467 1836 501
rect 2333 548 2367 582
rect 2333 476 2367 510
rect 2791 803 2825 837
rect 3264 764 3298 798
rect 3264 692 3298 726
rect 3071 564 3105 598
rect 3936 690 3970 724
rect 3714 622 3748 656
rect 3786 622 3820 656
rect 3936 618 3970 652
rect 2708 490 2742 524
rect 3071 492 3105 526
rect 3554 564 3588 598
rect 3554 492 3588 526
rect 3741 536 3775 570
rect 3741 464 3775 498
rect 4030 531 4064 565
rect 4030 459 4064 493
rect 4197 549 4231 583
rect 4197 477 4231 511
rect 4753 1080 4787 1114
rect 4825 1080 4859 1114
rect 7815 1080 7849 1114
rect 7887 1080 7921 1114
rect 4753 925 4787 959
rect 4825 925 4859 959
rect 7815 925 7849 959
rect 7887 925 7921 959
rect 4753 775 4787 809
rect 4825 775 4859 809
rect 7810 775 7844 809
rect 7882 775 7916 809
rect 4753 619 4787 653
rect 4825 619 4859 653
rect 7816 619 7850 653
rect 7888 619 7922 653
rect 2708 418 2742 452
<< metal1 >>
rect 235 3186 2723 3214
tri 235 3162 259 3186 nw
tri 2693 3162 2717 3186 ne
rect 2717 3162 2723 3186
rect 2775 3162 2787 3214
rect 2839 3162 2845 3214
rect 3107 3148 3113 3200
rect 3165 3148 3177 3200
rect 3229 3194 3235 3200
tri 3235 3194 3241 3200 sw
rect 3229 3171 5474 3194
tri 5474 3171 5497 3194 sw
rect 3229 3160 5497 3171
rect 3229 3148 3235 3160
tri 3235 3148 3247 3160 nw
tri 5454 3148 5466 3160 ne
rect 5466 3148 5497 3160
tri 5497 3148 5520 3171 sw
tri 5466 3138 5476 3148 ne
rect 5476 3138 5520 3148
tri 5520 3138 5530 3148 sw
rect 2479 3086 2485 3138
rect 2537 3086 2549 3138
rect 2601 3120 2607 3138
tri 2607 3120 2625 3138 sw
tri 5476 3120 5494 3138 ne
rect 5494 3120 5530 3138
tri 5530 3120 5548 3138 sw
rect 2601 3099 5416 3120
tri 5416 3099 5437 3120 sw
tri 5494 3117 5497 3120 ne
rect 5497 3117 5548 3120
tri 5548 3117 5551 3120 sw
rect 2601 3086 5437 3099
tri 5497 3087 5527 3117 ne
rect 5527 3087 6021 3117
rect 5383 3052 5437 3086
tri 5527 3083 5531 3087 ne
rect 5531 3083 6021 3087
rect 4861 2974 4867 3026
rect 4919 2974 4936 3026
rect 4988 2974 4994 3026
rect 5026 2970 5032 3022
rect 5084 2970 5098 3022
rect 5150 2970 5156 3022
rect 5201 2969 5207 3021
rect 5259 2969 5273 3021
rect 5325 2969 5331 3021
rect 5967 2987 6021 3083
rect 6132 3081 6184 3087
rect 6132 3015 6184 3029
rect 6132 2957 6184 2963
rect 6278 3081 6330 3087
rect 6278 3015 6330 3029
rect 6278 2957 6330 2963
rect 6432 3081 6484 3087
rect 6432 3015 6484 3029
rect 6432 2957 6484 2963
rect 2560 2838 2566 2890
rect 2618 2838 2630 2890
rect 2682 2838 2688 2890
rect 2974 2872 2980 2924
rect 3032 2872 3044 2924
rect 3096 2872 3469 2924
rect 3521 2872 3533 2924
rect 3585 2872 3591 2924
rect 187 2765 1220 2817
rect 1272 2765 1284 2817
rect 1336 2765 1342 2817
rect 1419 2765 1425 2817
rect 1477 2765 1489 2817
rect 1541 2765 1861 2817
rect 1913 2765 1925 2817
rect 1977 2765 1983 2817
rect 2051 2765 2057 2817
rect 2109 2765 2121 2817
rect 2173 2793 2179 2817
tri 2179 2793 2203 2817 sw
rect 3241 2793 3247 2817
rect 2173 2765 3247 2793
rect 3299 2765 3311 2817
rect 3363 2765 3369 2817
rect 3602 2649 3630 2677
rect 888 2599 934 2611
rect 888 2565 894 2599
rect 928 2565 934 2599
rect 888 2527 934 2565
rect 2415 2604 2545 2610
rect 2415 2570 2427 2604
rect 2533 2570 2545 2604
rect 2837 2594 4648 2607
rect 2415 2564 2447 2570
tri 2415 2538 2441 2564 ne
rect 2441 2552 2447 2564
rect 2499 2564 2545 2570
rect 2717 2578 2769 2584
rect 2499 2552 2505 2564
rect 2441 2540 2505 2552
rect 2441 2538 2447 2540
tri 2441 2532 2447 2538 ne
rect 888 2493 894 2527
rect 928 2515 934 2527
rect 928 2495 2268 2515
tri 2268 2495 2288 2515 sw
rect 928 2493 2288 2495
rect 888 2487 2288 2493
rect 888 2481 934 2487
tri 2200 2481 2206 2487 ne
rect 2206 2481 2288 2487
tri 2206 2472 2215 2481 ne
rect 2215 2472 2288 2481
tri 2288 2472 2311 2495 sw
rect 2499 2538 2505 2540
tri 2505 2538 2531 2564 nw
tri 2499 2532 2505 2538 nw
rect 2447 2482 2499 2488
rect 2717 2507 2769 2526
tri 2215 2461 2226 2472 ne
rect 2226 2461 2311 2472
tri 2226 2459 2228 2461 ne
rect 2228 2459 2311 2461
tri 953 2447 962 2456 se
rect 962 2447 1214 2456
tri 1214 2447 1223 2456 sw
rect 1390 2449 1442 2455
tri 942 2436 953 2447 se
rect 953 2436 1223 2447
tri 1223 2436 1234 2447 sw
tri 936 2430 942 2436 se
rect 942 2430 1246 2436
tri 922 2416 936 2430 se
rect 936 2428 1194 2430
rect 936 2416 962 2428
tri 962 2416 974 2428 nw
tri 1148 2416 1160 2428 ne
rect 1160 2416 1194 2428
tri 921 2415 922 2416 se
rect 922 2415 961 2416
tri 961 2415 962 2416 nw
tri 1160 2415 1161 2416 ne
rect 1161 2415 1194 2416
rect 714 2409 946 2415
rect 423 2376 553 2382
rect 423 2342 435 2376
rect 469 2342 507 2376
rect 541 2342 553 2376
rect 714 2375 726 2409
rect 760 2375 803 2409
rect 837 2400 946 2409
tri 946 2400 961 2415 nw
tri 1161 2400 1176 2415 ne
rect 1176 2400 1194 2415
rect 837 2396 942 2400
tri 942 2396 946 2400 nw
rect 1002 2396 1132 2400
tri 1132 2396 1136 2400 sw
tri 1176 2396 1180 2400 ne
rect 1180 2396 1194 2400
rect 1228 2396 1246 2430
tri 1371 2413 1390 2432 se
tri 1370 2412 1371 2413 se
rect 1371 2412 1390 2413
tri 1356 2398 1370 2412 se
rect 1370 2398 1390 2412
rect 837 2394 940 2396
tri 940 2394 942 2396 nw
rect 1002 2394 1136 2396
tri 1136 2394 1138 2396 sw
tri 1180 2394 1182 2396 ne
rect 837 2375 915 2394
rect 714 2369 915 2375
tri 915 2369 940 2394 nw
rect 1002 2360 1014 2394
rect 1048 2392 1138 2394
tri 1138 2392 1140 2394 sw
rect 1048 2360 1140 2392
rect 1002 2359 1140 2360
tri 1140 2359 1173 2392 sw
rect 1182 2390 1246 2396
rect 1296 2397 1390 2398
rect 1296 2392 1442 2397
rect 1002 2358 1173 2359
tri 1173 2358 1174 2359 sw
rect 1296 2358 1308 2392
rect 1342 2358 1380 2392
rect 1414 2385 1442 2392
rect 1002 2354 1174 2358
tri 1174 2354 1178 2358 sw
rect 423 2336 553 2342
tri 1123 2339 1138 2354 ne
rect 1138 2339 1178 2354
tri 1178 2339 1193 2354 sw
rect 1296 2352 1390 2358
tri 1365 2339 1378 2352 ne
rect 1378 2339 1390 2352
tri 1138 2338 1139 2339 ne
rect 1139 2338 1193 2339
tri 1193 2338 1194 2339 sw
tri 1378 2338 1379 2339 ne
rect 1379 2338 1390 2339
tri 1139 2336 1141 2338 ne
rect 1141 2336 1194 2338
tri 1141 2325 1152 2336 ne
rect 1152 2325 1194 2336
tri 1194 2325 1207 2338 sw
tri 1379 2327 1390 2338 ne
rect 1390 2327 1442 2333
rect 1470 2452 1522 2459
rect 1470 2385 1522 2400
rect 1470 2327 1522 2333
rect 1574 2452 1626 2458
rect 1735 2453 1787 2459
rect 1574 2388 1626 2400
rect 1718 2430 1735 2436
tri 2228 2446 2241 2459 ne
rect 2241 2446 2311 2459
rect 2837 2560 2843 2594
rect 2877 2563 4648 2594
rect 2877 2560 2909 2563
rect 2837 2555 2909 2560
tri 2909 2555 2917 2563 nw
tri 4634 2555 4642 2563 ne
rect 4642 2555 4648 2563
rect 4700 2555 4712 2607
rect 4764 2555 4770 2607
rect 5606 2567 5634 2595
rect 2837 2534 2888 2555
tri 2888 2534 2909 2555 nw
rect 2837 2522 2883 2534
tri 2883 2529 2888 2534 nw
tri 3243 2529 3248 2534 se
rect 3248 2531 3594 2534
tri 3594 2531 3597 2534 sw
rect 3248 2529 3597 2531
tri 3239 2525 3243 2529 se
rect 3243 2525 3597 2529
tri 3597 2525 3603 2531 sw
rect 3723 2525 4300 2531
rect 2837 2488 2843 2522
rect 2877 2488 2883 2522
tri 3225 2511 3239 2525 se
rect 3239 2511 3603 2525
tri 3603 2511 3617 2525 sw
rect 2837 2476 2883 2488
rect 3122 2505 3174 2511
rect 2912 2480 2964 2486
rect 2717 2449 2769 2455
rect 1787 2430 1848 2436
rect 1718 2396 1730 2430
rect 1787 2401 1802 2430
rect 1764 2396 1802 2401
rect 1836 2396 1848 2430
rect 1718 2390 1848 2396
rect 2003 2434 2049 2446
tri 2241 2439 2248 2446 ne
rect 2003 2400 2009 2434
rect 2043 2400 2049 2434
rect 1574 2326 1626 2336
rect 1735 2387 1787 2390
rect 2003 2359 2049 2400
rect 2248 2433 2311 2446
rect 2248 2399 2260 2433
rect 2294 2399 2311 2433
rect 2248 2393 2311 2399
rect 2435 2433 2502 2439
tri 2911 2438 2912 2439 se
rect 2435 2399 2447 2433
rect 2481 2399 2502 2433
tri 2878 2405 2911 2438 se
rect 2911 2428 2912 2438
rect 2911 2416 2964 2428
rect 2911 2405 2912 2416
tri 2415 2365 2435 2385 se
rect 2435 2365 2502 2399
tri 2412 2362 2415 2365 se
rect 2415 2362 2502 2365
tri 2409 2359 2412 2362 se
rect 2412 2359 2499 2362
tri 2499 2359 2502 2362 nw
rect 2542 2399 2912 2405
rect 2542 2365 2554 2399
rect 2588 2365 2626 2399
rect 2660 2365 2912 2399
rect 2542 2364 2912 2365
rect 2542 2359 2964 2364
tri 1881 2354 1886 2359 se
rect 1886 2354 2009 2359
rect 1735 2329 1787 2335
tri 1856 2329 1881 2354 se
rect 1881 2329 2009 2354
tri 1853 2326 1856 2329 se
rect 1856 2326 2009 2329
tri 1852 2325 1853 2326 se
rect 1853 2325 2009 2326
rect 2043 2331 2471 2359
tri 2471 2331 2499 2359 nw
tri 2911 2358 2912 2359 ne
rect 2912 2358 2964 2359
rect 3007 2444 3059 2450
rect 3007 2377 3059 2392
rect 3122 2441 3174 2453
rect 3122 2380 3174 2389
tri 3209 2495 3225 2511 se
rect 3225 2495 3617 2511
rect 3209 2492 3617 2495
rect 3209 2491 3285 2492
tri 3285 2491 3286 2492 nw
tri 3578 2491 3579 2492 ne
rect 3579 2491 3617 2492
tri 3617 2491 3637 2511 sw
rect 3723 2491 3735 2525
rect 3769 2491 3807 2525
rect 3841 2491 4300 2525
rect 3209 2480 3274 2491
tri 3274 2480 3285 2491 nw
tri 3579 2480 3590 2491 ne
rect 3590 2485 3637 2491
tri 3637 2485 3643 2491 sw
rect 3723 2485 4300 2491
rect 3590 2480 3643 2485
tri 3643 2480 3648 2485 sw
rect 3209 2438 3255 2480
tri 3255 2461 3274 2480 nw
tri 3590 2476 3594 2480 ne
rect 3594 2476 3648 2480
tri 3594 2464 3606 2476 ne
rect 3209 2404 3215 2438
rect 3249 2404 3255 2438
rect 3209 2365 3255 2404
tri 3179 2331 3209 2361 se
rect 3209 2331 3215 2365
rect 3249 2331 3255 2365
rect 2043 2325 2462 2331
tri 1152 2322 1155 2325 ne
rect 1155 2324 1207 2325
tri 1207 2324 1208 2325 sw
tri 1851 2324 1852 2325 se
rect 1852 2324 2462 2325
rect 1155 2322 1208 2324
tri 1208 2322 1210 2324 sw
tri 1849 2322 1851 2324 se
rect 1851 2322 2462 2324
tri 2462 2322 2471 2331 nw
tri 3175 2327 3179 2331 se
rect 3179 2327 3255 2331
tri 1155 2301 1176 2322 ne
rect 1176 2313 1210 2322
tri 1210 2313 1219 2322 sw
tri 1840 2313 1849 2322 se
rect 1849 2313 2453 2322
tri 2453 2313 2462 2322 nw
rect 3007 2319 3059 2325
rect 1176 2309 1219 2313
tri 1219 2309 1223 2313 sw
tri 1836 2309 1840 2313 se
rect 1840 2309 1876 2313
tri 1876 2309 1880 2313 nw
rect 1176 2301 1223 2309
tri 1223 2301 1231 2309 sw
tri 1828 2301 1836 2309 se
rect 1836 2301 1868 2309
tri 1868 2301 1876 2309 nw
tri 1176 2299 1178 2301 ne
rect 1178 2299 1231 2301
tri 1231 2299 1233 2301 sw
tri 1826 2299 1828 2301 se
rect 1828 2299 1866 2301
tri 1866 2299 1868 2301 nw
tri 1178 2292 1185 2299 ne
rect 1185 2297 1233 2299
tri 1233 2297 1235 2299 sw
tri 1824 2297 1826 2299 se
rect 1826 2297 1852 2299
rect 1185 2292 1852 2297
rect 1097 2280 1143 2292
rect 1097 2246 1103 2280
rect 1137 2246 1143 2280
tri 1185 2269 1208 2292 ne
rect 1208 2285 1852 2292
tri 1852 2285 1866 2299 nw
rect 1208 2269 1836 2285
tri 1836 2269 1852 2285 nw
tri 1883 2269 1899 2285 se
rect 1899 2269 2969 2285
tri 2969 2269 2985 2285 sw
rect 3136 2281 3255 2327
rect 3302 2418 3348 2440
rect 3302 2384 3308 2418
rect 3342 2384 3348 2418
tri 3296 2281 3302 2287 se
rect 3302 2281 3348 2384
rect 3510 2428 3556 2440
rect 3510 2394 3516 2428
rect 3550 2394 3556 2428
rect 3510 2356 3556 2394
rect 3510 2322 3516 2356
rect 3550 2322 3556 2356
tri 3284 2269 3296 2281 se
rect 3296 2269 3348 2281
tri 1881 2267 1883 2269 se
rect 1883 2267 2985 2269
tri 2985 2267 2987 2269 sw
tri 3282 2267 3284 2269 se
rect 3284 2267 3348 2269
tri 3348 2267 3368 2287 sw
tri 3490 2267 3510 2287 se
rect 3510 2267 3556 2322
tri 3600 2301 3606 2307 se
rect 3606 2301 3648 2476
tri 4220 2457 4248 2485 ne
rect 4248 2457 4300 2485
tri 4835 2489 4841 2495 se
rect 4835 2483 4887 2489
tri 4503 2475 4505 2477 se
rect 4505 2475 4711 2477
tri 4711 2475 4713 2477 sw
rect 4073 2451 4125 2457
tri 4248 2451 4254 2457 ne
rect 4073 2390 4082 2399
rect 4116 2390 4125 2399
rect 4073 2387 4125 2390
rect 3895 2374 4025 2380
rect 3895 2340 3907 2374
rect 3941 2340 3979 2374
rect 4013 2340 4025 2374
rect 3895 2334 4025 2340
rect 4254 2424 4300 2457
tri 4462 2434 4503 2475 se
rect 4503 2434 4713 2475
rect 4254 2390 4260 2424
rect 4294 2390 4300 2424
rect 4254 2378 4300 2390
rect 4350 2431 4713 2434
rect 4350 2428 4505 2431
rect 4350 2394 4362 2428
rect 4396 2394 4434 2428
rect 4468 2411 4505 2428
tri 4505 2411 4525 2431 nw
tri 4691 2411 4711 2431 ne
rect 4711 2411 4713 2431
rect 4468 2410 4504 2411
tri 4504 2410 4505 2411 nw
tri 4711 2410 4712 2411 ne
rect 4712 2410 4713 2411
rect 4468 2409 4503 2410
tri 4503 2409 4504 2410 nw
tri 4712 2409 4713 2410 ne
tri 4713 2409 4779 2475 sw
rect 4468 2394 4482 2409
rect 4350 2388 4482 2394
tri 4482 2388 4503 2409 nw
tri 4713 2389 4733 2409 ne
tri 4532 2357 4544 2369 se
rect 4544 2357 4590 2369
tri 4521 2346 4532 2357 se
rect 4532 2346 4550 2357
rect 4073 2329 4125 2335
tri 4157 2301 4169 2313 se
rect 4169 2301 4215 2313
tri 1867 2253 1881 2267 se
rect 1881 2257 2987 2267
rect 1881 2253 1908 2257
tri 1908 2253 1912 2257 nw
tri 2949 2253 2953 2257 ne
rect 2953 2253 2987 2257
tri 2987 2253 3001 2267 sw
tri 3268 2253 3282 2267 se
rect 3282 2253 3368 2267
tri 3368 2253 3382 2267 sw
tri 3476 2253 3490 2267 se
rect 3490 2253 3556 2267
tri 1865 2251 1867 2253 se
rect 1867 2251 1906 2253
tri 1906 2251 1908 2253 nw
tri 2953 2251 2955 2253 ne
rect 2955 2251 3556 2253
rect 1097 2214 1143 2246
tri 1858 2244 1865 2251 se
rect 1865 2244 1899 2251
tri 1899 2244 1906 2251 nw
tri 2955 2244 2962 2251 ne
rect 2962 2244 3556 2251
tri 1855 2241 1858 2244 se
rect 1858 2241 1896 2244
tri 1896 2241 1899 2244 nw
tri 2962 2241 2965 2244 ne
rect 2965 2241 3556 2244
rect 1097 2208 1224 2214
rect 1097 2174 1103 2208
rect 1137 2201 1224 2208
tri 1224 2201 1237 2214 sw
rect 1137 2195 1237 2201
tri 1237 2195 1243 2201 sw
rect 1137 2189 1243 2195
tri 1243 2189 1249 2195 sw
rect 1688 2189 1694 2241
rect 1746 2189 1758 2241
rect 1810 2229 1884 2241
tri 1884 2229 1896 2241 nw
tri 2965 2237 2969 2241 ne
rect 2969 2237 3556 2241
tri 2969 2229 2977 2237 ne
rect 2977 2229 3556 2237
rect 1810 2225 1880 2229
tri 1880 2225 1884 2229 nw
tri 2977 2225 2981 2229 ne
rect 2981 2225 3556 2229
tri 3596 2297 3600 2301 se
rect 3600 2297 3648 2301
rect 3596 2291 3648 2297
tri 4132 2276 4157 2301 se
rect 4157 2276 4175 2301
rect 3596 2227 3648 2239
rect 1810 2213 1868 2225
tri 1868 2213 1880 2225 nw
rect 1810 2189 1816 2213
rect 1137 2174 1249 2189
rect 1097 2162 1249 2174
tri 1202 2127 1237 2162 ne
rect 1237 2151 1249 2162
tri 1249 2151 1287 2189 sw
rect 3596 2169 3648 2175
rect 3908 2270 4175 2276
rect 3960 2267 4175 2270
rect 4209 2267 4215 2301
rect 4462 2294 4468 2346
rect 4520 2294 4532 2346
rect 4584 2294 4590 2357
tri 4510 2285 4519 2294 ne
rect 4519 2285 4590 2294
rect 3960 2229 4215 2267
tri 4519 2260 4544 2285 ne
rect 4544 2251 4550 2285
rect 4584 2251 4590 2285
rect 4544 2239 4590 2251
tri 4684 2239 4733 2288 se
rect 4733 2268 4779 2409
rect 4835 2419 4887 2431
rect 4835 2361 4887 2367
tri 4835 2355 4841 2361 ne
rect 3960 2218 4175 2229
rect 3908 2204 4175 2218
rect 3960 2195 4175 2204
rect 4209 2195 4215 2229
tri 4670 2225 4684 2239 se
rect 4684 2225 4733 2239
tri 4667 2222 4670 2225 se
rect 4670 2222 4733 2225
tri 4733 2222 4779 2268 nw
tri 4658 2213 4667 2222 se
rect 4667 2213 4720 2222
rect 3960 2183 4215 2195
tri 4654 2209 4658 2213 se
rect 4658 2209 4720 2213
tri 4720 2209 4733 2222 nw
rect 1237 2127 1287 2151
tri 1287 2127 1311 2151 sw
tri 2779 2127 2803 2151 se
rect 2803 2127 2809 2151
tri 1237 2099 1265 2127 ne
rect 1265 2099 2809 2127
rect 2861 2099 2873 2151
rect 2925 2099 2931 2151
rect 3908 2146 3960 2152
tri 3960 2146 3997 2183 nw
rect 3602 2033 3630 2061
rect 1574 1893 1580 1945
rect 1632 1893 1644 1945
rect 1696 1936 3549 1945
rect 1696 1893 3122 1936
tri 3088 1863 3118 1893 ne
rect 3118 1884 3122 1893
rect 3174 1933 3549 1936
rect 3174 1899 3509 1933
rect 3543 1899 3549 1933
rect 3174 1893 3549 1899
rect 3174 1884 3176 1893
rect 3118 1872 3176 1884
rect 3118 1863 3122 1872
tri 1198 1861 1200 1863 se
rect 1200 1861 2429 1863
tri 1165 1828 1198 1861 se
rect 1198 1835 2429 1861
rect 1198 1828 1215 1835
tri 1215 1828 1222 1835 nw
tri 2399 1828 2406 1835 ne
rect 2406 1828 2429 1835
tri 1152 1815 1165 1828 se
rect 1165 1815 1202 1828
tri 1202 1815 1215 1828 nw
tri 2406 1815 2419 1828 ne
rect 2419 1815 2429 1828
tri 1150 1813 1152 1815 se
rect 1152 1813 1200 1815
tri 1200 1813 1202 1815 nw
tri 2419 1813 2421 1815 ne
rect 2421 1813 2429 1815
tri 1138 1801 1150 1813 se
rect 1150 1801 1188 1813
tri 1188 1801 1200 1813 nw
tri 2421 1811 2423 1813 ne
rect 2423 1811 2429 1813
rect 2481 1811 2493 1863
rect 2545 1811 2551 1863
tri 3118 1861 3120 1863 ne
rect 3120 1861 3122 1863
tri 3120 1859 3122 1861 ne
rect 3174 1861 3176 1872
tri 3176 1861 3208 1893 nw
tri 3469 1861 3501 1893 ne
rect 3501 1861 3549 1893
tri 3174 1859 3176 1861 nw
rect 3122 1814 3174 1820
rect 3297 1855 3349 1861
tri 3501 1859 3503 1861 ne
rect 1861 1801 2253 1807
tri 1104 1767 1138 1801 se
rect 1138 1767 1154 1801
tri 1154 1767 1188 1801 nw
rect 982 1759 1034 1767
tri 1100 1763 1104 1767 se
rect 1104 1763 1150 1767
tri 1150 1763 1154 1767 nw
tri 1099 1762 1100 1763 se
rect 1100 1762 1149 1763
tri 1149 1762 1150 1763 nw
rect 1483 1762 1529 1774
rect 900 1711 946 1724
rect 900 1677 906 1711
rect 940 1677 946 1711
rect 709 1656 780 1662
rect 709 1622 721 1656
rect 755 1649 780 1656
tri 780 1649 787 1656 sw
rect 755 1622 787 1649
rect 709 1616 787 1622
tri 787 1616 820 1649 sw
rect 900 1632 946 1677
rect 982 1695 1034 1707
rect 982 1637 1034 1643
tri 1072 1735 1099 1762 se
rect 1099 1737 1124 1762
tri 1124 1737 1149 1762 nw
rect 1099 1735 1122 1737
tri 1122 1735 1124 1737 nw
tri 1165 1735 1167 1737 se
rect 1167 1735 1280 1737
tri 1280 1735 1282 1737 sw
rect 1072 1728 1115 1735
tri 1115 1728 1122 1735 nw
tri 1158 1728 1165 1735 se
rect 1165 1728 1282 1735
tri 1282 1728 1289 1735 sw
rect 1483 1728 1489 1762
rect 1523 1728 1529 1762
rect 1072 1725 1112 1728
tri 1112 1725 1115 1728 nw
tri 1155 1725 1158 1728 se
rect 1158 1725 1289 1728
tri 1289 1725 1292 1728 sw
rect 1072 1721 1108 1725
tri 1108 1721 1112 1725 nw
tri 1151 1721 1155 1725 se
rect 1155 1721 1292 1725
tri 1292 1721 1296 1725 sw
tri 946 1632 947 1633 sw
rect 900 1628 947 1632
tri 900 1616 912 1628 ne
rect 912 1616 947 1628
tri 947 1616 963 1632 sw
tri 1056 1616 1072 1632 se
rect 1072 1616 1100 1721
tri 1100 1713 1108 1721 nw
tri 1143 1713 1151 1721 se
rect 1151 1713 1296 1721
tri 1296 1713 1304 1721 sw
tri 1139 1709 1143 1713 se
rect 1143 1709 1304 1713
tri 1304 1709 1308 1713 sw
tri 1131 1701 1139 1709 se
rect 1139 1701 1177 1709
tri 1177 1701 1185 1709 nw
tri 1242 1701 1250 1709 ne
rect 1250 1701 1308 1709
tri 1308 1701 1316 1709 sw
tri 754 1609 761 1616 ne
rect 761 1609 820 1616
tri 820 1609 827 1616 sw
tri 912 1609 919 1616 ne
rect 919 1614 963 1616
tri 963 1614 965 1616 sw
tri 1054 1614 1056 1616 se
rect 1056 1614 1100 1616
rect 919 1609 965 1614
tri 761 1603 767 1609 ne
rect 767 1603 827 1609
tri 827 1603 833 1609 sw
tri 919 1603 925 1609 ne
rect 925 1603 965 1609
tri 965 1603 976 1614 sw
tri 1043 1603 1054 1614 se
rect 1054 1610 1100 1614
rect 1054 1603 1093 1610
tri 1093 1603 1100 1610 nw
tri 1128 1698 1131 1701 se
rect 1131 1698 1174 1701
tri 1174 1698 1177 1701 nw
tri 1250 1698 1253 1701 ne
rect 1253 1698 1316 1701
rect 1128 1690 1166 1698
tri 1166 1690 1174 1698 nw
tri 1253 1690 1261 1698 ne
rect 1261 1690 1316 1698
tri 1316 1690 1327 1701 sw
rect 1483 1690 1529 1728
rect 1128 1685 1161 1690
tri 1161 1685 1166 1690 nw
tri 1261 1685 1266 1690 ne
rect 1266 1685 1327 1690
tri 1327 1685 1332 1690 sw
tri 767 1590 780 1603 ne
rect 780 1600 833 1603
tri 833 1600 836 1603 sw
tri 925 1600 928 1603 ne
rect 928 1600 976 1603
tri 976 1600 979 1603 sw
tri 1040 1600 1043 1603 se
rect 1043 1600 1090 1603
tri 1090 1600 1093 1603 nw
rect 780 1591 836 1600
tri 836 1591 845 1600 sw
tri 928 1591 937 1600 ne
rect 937 1591 1081 1600
tri 1081 1591 1090 1600 nw
rect 780 1590 845 1591
tri 780 1578 792 1590 ne
rect 792 1588 845 1590
tri 845 1588 848 1591 sw
tri 937 1588 940 1591 ne
rect 940 1588 1078 1591
tri 1078 1588 1081 1591 nw
rect 792 1582 848 1588
tri 848 1582 854 1588 sw
tri 940 1582 946 1588 ne
rect 946 1582 1072 1588
tri 1072 1582 1078 1588 nw
rect 792 1578 854 1582
tri 854 1578 858 1582 sw
tri 946 1578 950 1582 ne
rect 950 1578 1068 1582
tri 1068 1578 1072 1582 nw
tri 1126 1578 1128 1580 se
rect 1128 1578 1156 1685
tri 1156 1680 1161 1685 nw
tri 1266 1680 1271 1685 ne
rect 1271 1680 1427 1685
tri 1271 1671 1280 1680 ne
rect 1280 1671 1427 1680
tri 1280 1662 1289 1671 ne
rect 1289 1662 1427 1671
tri 792 1544 826 1578 ne
rect 826 1572 858 1578
tri 858 1572 864 1578 sw
tri 950 1572 956 1578 ne
rect 956 1572 1062 1578
tri 1062 1572 1068 1578 nw
tri 1120 1572 1126 1578 se
rect 1126 1572 1156 1578
rect 826 1544 864 1572
tri 864 1544 892 1572 sw
tri 1092 1544 1120 1572 se
rect 1120 1564 1156 1572
rect 1120 1544 1136 1564
tri 1136 1544 1156 1564 nw
rect 1184 1650 1230 1662
tri 1289 1660 1291 1662 ne
rect 1291 1660 1427 1662
rect 1184 1616 1190 1650
rect 1224 1616 1230 1650
tri 1291 1626 1325 1660 ne
rect 1325 1626 1387 1660
rect 1421 1637 1427 1660
rect 1483 1656 1489 1690
rect 1523 1656 1529 1690
tri 1427 1637 1440 1650 sw
rect 1483 1644 1529 1656
rect 1580 1768 1632 1774
rect 1861 1767 1873 1801
rect 1907 1767 1947 1801
rect 1981 1767 2201 1801
rect 1861 1761 2201 1767
tri 2175 1756 2180 1761 ne
rect 2180 1756 2201 1761
tri 2180 1735 2201 1756 ne
rect 2728 1797 2774 1809
rect 2613 1783 2665 1789
rect 2201 1737 2253 1749
rect 1580 1702 1632 1716
rect 2127 1709 2173 1721
rect 1963 1701 2093 1707
rect 1963 1667 1975 1701
rect 2009 1667 2047 1701
rect 2081 1667 2093 1701
rect 1963 1661 2093 1667
rect 2127 1675 2133 1709
rect 2167 1675 2173 1709
rect 2201 1679 2253 1685
rect 2424 1775 2476 1781
rect 2424 1710 2476 1723
rect 2613 1719 2665 1731
rect 1580 1644 1632 1650
tri 2122 1644 2127 1649 se
rect 2127 1644 2173 1675
rect 2541 1701 2613 1707
rect 2728 1763 2734 1797
rect 2768 1763 2774 1797
rect 3503 1827 3509 1861
rect 3543 1827 3549 1861
rect 3503 1815 3549 1827
rect 3786 1933 4023 1945
rect 3786 1899 3792 1933
rect 3826 1899 4023 1933
rect 3786 1893 4023 1899
rect 4075 1893 4087 1945
rect 4139 1893 4145 1945
rect 3786 1861 3832 1893
rect 3786 1827 3792 1861
rect 3826 1827 3832 1861
tri 3832 1859 3866 1893 nw
rect 3786 1815 3832 1827
rect 3297 1794 3307 1803
rect 3341 1794 3349 1803
rect 3297 1791 3349 1794
rect 2728 1725 2774 1763
rect 3202 1780 3254 1786
rect 2541 1667 2553 1701
rect 2587 1667 2613 1701
rect 2665 1667 2671 1707
rect 2728 1691 2734 1725
rect 2768 1691 2774 1725
rect 2728 1679 2774 1691
rect 2985 1738 3037 1744
rect 3202 1716 3254 1728
rect 2541 1661 2671 1667
rect 2985 1674 3037 1686
tri 3187 1685 3202 1700 se
tri 3168 1666 3187 1685 se
rect 3187 1666 3202 1685
rect 2424 1652 2476 1658
rect 2822 1656 2893 1662
tri 2115 1637 2122 1644 se
rect 2122 1637 2173 1644
rect 1421 1626 1440 1637
rect 1184 1588 1230 1616
tri 1325 1614 1337 1626 ne
rect 1337 1616 1440 1626
tri 1440 1616 1461 1637 sw
tri 2094 1616 2115 1637 se
rect 2115 1616 2133 1637
rect 1337 1614 2133 1616
tri 1337 1603 1348 1614 ne
rect 1348 1603 2133 1614
rect 2167 1623 2173 1637
tri 2173 1623 2200 1650 sw
tri 2795 1623 2822 1650 se
rect 2822 1623 2834 1656
rect 2167 1622 2460 1623
tri 2460 1622 2461 1623 sw
tri 2794 1622 2795 1623 se
rect 2795 1622 2834 1623
rect 2868 1622 2893 1656
rect 2167 1616 2461 1622
tri 2461 1616 2467 1622 sw
tri 2788 1616 2794 1622 se
rect 2794 1616 2893 1622
rect 2985 1616 3037 1622
rect 3105 1664 3202 1666
rect 3297 1722 3307 1739
rect 3341 1722 3349 1739
rect 3297 1710 3349 1722
rect 3425 1776 3477 1782
rect 3425 1712 3477 1724
rect 3105 1660 3254 1664
rect 3105 1626 3117 1660
rect 3151 1626 3189 1660
rect 3223 1626 3254 1660
rect 3425 1654 3477 1660
rect 3891 1685 4021 1691
rect 3891 1651 3903 1685
rect 3937 1651 3975 1685
rect 4009 1651 4021 1685
rect 3891 1645 4021 1651
rect 3105 1620 3254 1626
rect 2167 1603 2893 1616
tri 1230 1588 1236 1594 sw
rect 1348 1591 2893 1603
rect 1348 1588 2140 1591
tri 2140 1588 2143 1591 nw
tri 2421 1588 2424 1591 ne
rect 2424 1588 2893 1591
tri 4633 1588 4654 1609 se
rect 4654 1588 4708 2209
tri 4708 2197 4720 2209 nw
rect 5870 1654 5876 1706
rect 5928 1654 5940 1706
rect 5992 1654 5998 1706
rect 1184 1578 1236 1588
rect 1184 1544 1190 1578
rect 1224 1560 1236 1578
tri 1236 1560 1264 1588 sw
tri 4606 1561 4633 1588 se
rect 4633 1587 4708 1588
rect 4633 1561 4654 1587
tri 2152 1560 2153 1561 se
rect 2153 1560 2205 1561
rect 1224 1555 2205 1560
rect 1224 1544 2153 1555
tri 826 1543 827 1544 ne
rect 827 1543 892 1544
tri 892 1543 893 1544 sw
tri 1091 1543 1092 1544 se
rect 1092 1543 1135 1544
tri 1135 1543 1136 1544 nw
tri 827 1515 855 1543 ne
rect 855 1515 1107 1543
tri 1107 1515 1135 1543 nw
rect 1184 1532 2153 1544
tri 2119 1515 2136 1532 ne
rect 2136 1515 2153 1532
tri 2136 1498 2153 1515 ne
tri 4588 1543 4606 1561 se
rect 4606 1543 4654 1561
tri 4578 1533 4588 1543 se
rect 4588 1533 4654 1543
tri 4654 1533 4708 1587 nw
tri 4560 1515 4578 1533 se
rect 4578 1515 4606 1533
rect 2153 1491 2205 1503
rect 1444 1484 1751 1490
rect 1444 1450 1705 1484
rect 1739 1450 1751 1484
rect 1444 1444 1751 1450
tri 4535 1490 4560 1515 se
rect 4560 1490 4606 1515
tri 4530 1485 4535 1490 se
rect 4535 1485 4606 1490
tri 4606 1485 4654 1533 nw
rect 2153 1433 2205 1439
rect 4397 1433 4403 1485
rect 4455 1433 4467 1485
rect 4519 1444 4565 1485
tri 4565 1444 4606 1485 nw
rect 4519 1433 4554 1444
tri 4554 1433 4565 1444 nw
rect 3602 1370 3630 1398
rect 5233 1323 5261 1351
rect 7694 1295 7700 1347
rect 7752 1295 7764 1347
rect 7816 1313 8247 1347
tri 8247 1313 8281 1347 sw
rect 7816 1295 8281 1313
tri 8183 1272 8206 1295 ne
rect 8206 1272 8281 1295
tri 6385 1249 6408 1272 ne
rect 6408 1249 6665 1272
tri 6665 1249 6688 1272 nw
tri 8206 1249 8229 1272 ne
tri 6408 1238 6419 1249 ne
rect 6419 1238 6654 1249
tri 6654 1238 6665 1249 nw
rect 1762 1201 4148 1203
rect 1762 1197 4331 1201
rect 1762 1163 1774 1197
rect 1808 1163 1847 1197
rect 1881 1163 1920 1197
rect 1954 1163 1993 1197
rect 2027 1163 2066 1197
rect 2100 1163 2139 1197
rect 2173 1163 2212 1197
rect 2246 1163 2285 1197
rect 2319 1163 2358 1197
rect 2392 1163 2431 1197
rect 2465 1163 2504 1197
rect 2538 1163 2577 1197
rect 2611 1163 2650 1197
rect 2684 1163 2723 1197
rect 2757 1163 2796 1197
rect 2830 1163 2869 1197
rect 2903 1163 2942 1197
rect 2976 1163 3015 1197
rect 3049 1163 3088 1197
rect 3122 1163 3161 1197
rect 3195 1163 3234 1197
rect 3268 1163 3307 1197
rect 3341 1163 3380 1197
rect 3414 1163 3453 1197
rect 3487 1163 3526 1197
rect 3560 1163 3598 1197
rect 3632 1163 3670 1197
rect 3704 1163 3742 1197
rect 3776 1163 3814 1197
rect 3848 1163 3886 1197
rect 3920 1163 3958 1197
rect 3992 1163 4030 1197
rect 4064 1163 4102 1197
rect 4136 1163 4331 1197
rect 1762 1157 4331 1163
rect 2489 999 2572 1157
rect 2499 998 2572 999
rect 3432 998 4331 1157
rect 4913 1155 4919 1207
rect 4971 1155 4983 1207
rect 5035 1155 5041 1207
rect 6419 1154 6631 1238
tri 6631 1215 6654 1238 nw
rect 7043 1155 7049 1207
rect 7101 1155 7123 1207
rect 7175 1155 7181 1207
tri 7181 1201 7187 1207 sw
tri 4731 1080 4741 1090 se
rect 4741 1080 4747 1124
tri 4725 1074 4731 1080 se
rect 4731 1074 4747 1080
tri 4723 1072 4725 1074 se
rect 4725 1072 4747 1074
rect 4799 1072 4813 1124
rect 4865 1072 4871 1124
rect 7803 1073 7809 1125
rect 7861 1073 7875 1125
rect 7927 1073 7933 1125
tri 4687 1036 4723 1072 se
rect 4723 1036 4753 1072
tri 4753 1036 4789 1072 nw
tri 4649 998 4687 1036 se
rect 4687 998 4715 1036
tri 4715 998 4753 1036 nw
tri 4621 970 4649 998 se
rect 4649 970 4687 998
tri 4687 970 4715 998 nw
tri 4615 964 4621 970 se
rect 4621 969 4686 970
tri 4686 969 4687 970 nw
rect 4621 968 4685 969
tri 4685 968 4686 969 nw
rect 4621 964 4681 968
tri 4681 964 4685 968 nw
tri 4734 964 4738 968 se
rect 4738 964 4747 968
rect 3782 958 3788 964
rect 3134 952 3788 958
rect 2785 909 2831 921
rect 3134 918 3146 952
rect 3180 918 3218 952
rect 3252 918 3788 952
rect 3134 912 3788 918
rect 3840 912 3852 964
rect 3904 958 3910 964
tri 4610 959 4615 964 se
rect 4615 959 4676 964
tri 4676 959 4681 964 nw
tri 4729 959 4734 964 se
rect 4734 959 4747 964
tri 4609 958 4610 959 se
rect 4610 958 4675 959
tri 4675 958 4676 959 nw
tri 4728 958 4729 959 se
rect 4729 958 4747 959
rect 3904 912 4073 958
tri 4576 925 4609 958 se
rect 4609 925 4642 958
tri 4642 925 4675 958 nw
tri 4695 925 4728 958 se
rect 4728 925 4747 958
tri 4563 912 4576 925 se
rect 4576 917 4634 925
tri 4634 917 4642 925 nw
tri 4687 917 4695 925 se
rect 4695 917 4747 925
rect 4576 916 4633 917
tri 4633 916 4634 917 nw
tri 4686 916 4687 917 se
rect 4687 916 4747 917
rect 4799 916 4813 968
rect 4865 916 4871 968
rect 7803 917 7809 969
rect 7861 917 7875 969
rect 7927 917 7933 969
rect 4576 912 4629 916
tri 4629 912 4633 916 nw
tri 4682 912 4686 916 se
rect 4686 912 4748 916
tri 4748 912 4752 916 nw
rect 2785 875 2791 909
rect 2825 884 2831 909
tri 4555 904 4563 912 se
rect 4563 904 4621 912
tri 4621 904 4629 912 nw
tri 4674 904 4682 912 se
rect 4682 904 4732 912
tri 4535 884 4555 904 se
rect 4555 896 4613 904
tri 4613 896 4621 904 nw
tri 4666 896 4674 904 se
rect 4674 896 4732 904
tri 4732 896 4748 912 nw
rect 4555 884 4601 896
tri 4601 884 4613 896 nw
tri 4654 884 4666 896 se
rect 4666 884 4720 896
tri 4720 884 4732 896 nw
rect 8229 891 8281 1272
rect 2825 875 4568 884
rect 2785 851 4568 875
tri 4568 851 4601 884 nw
tri 4621 851 4654 884 se
rect 4654 851 4674 884
rect 1842 836 1972 842
rect 1842 802 1854 836
rect 1888 802 1926 836
rect 1960 802 1972 836
rect 2785 838 4555 851
tri 4555 838 4568 851 nw
tri 4608 838 4621 851 se
rect 4621 838 4674 851
tri 4674 838 4720 884 nw
rect 2785 837 2831 838
rect 1842 796 1972 802
rect 2619 820 2665 832
rect 2619 786 2625 820
rect 2659 786 2665 820
rect 2785 803 2791 837
rect 2825 803 2831 837
tri 4600 830 4608 838 se
rect 4608 830 4666 838
tri 4666 830 4674 838 nw
tri 4580 810 4600 830 se
rect 4600 815 4651 830
tri 4651 815 4666 830 nw
rect 8229 827 8281 839
rect 4600 810 4646 815
tri 4646 810 4651 815 nw
rect 2785 791 2831 803
rect 3258 809 4645 810
tri 4645 809 4646 810 nw
rect 3258 798 4611 809
rect 2240 762 2286 774
rect 1973 728 2019 730
rect 2156 728 2202 730
rect 2240 728 2246 762
rect 2280 728 2286 762
rect 1970 722 2022 728
rect 1970 658 2022 670
rect 1970 600 2022 606
rect 2153 722 2205 728
rect 2153 658 2205 670
rect 2240 690 2286 728
rect 2619 748 2665 786
rect 2619 714 2625 748
rect 2659 714 2665 748
rect 3258 764 3264 798
rect 3298 775 4611 798
tri 4611 775 4645 809 nw
rect 3298 769 4605 775
tri 4605 769 4611 775 nw
rect 3298 764 4600 769
tri 4600 764 4605 769 nw
rect 4741 766 4747 818
rect 4799 766 4813 818
rect 4865 766 4871 818
tri 2733 729 2747 743 se
rect 2747 729 3154 743
tri 3154 729 3168 743 sw
tri 2730 726 2733 729 se
rect 2733 726 3168 729
tri 3168 726 3171 729 sw
rect 3258 726 3337 764
rect 7798 763 7804 815
rect 7856 763 7875 815
rect 7927 763 7933 815
rect 8229 769 8281 775
rect 2619 702 2665 714
tri 2707 703 2730 726 se
rect 2730 715 3171 726
rect 2730 703 2747 715
tri 2747 703 2759 715 nw
tri 3142 703 3154 715 ne
rect 3154 703 3171 715
tri 2706 702 2707 703 se
rect 2707 702 2736 703
tri 2696 692 2706 702 se
rect 2706 692 2736 702
tri 2736 692 2747 703 nw
tri 3154 692 3165 703 ne
rect 3165 692 3171 703
tri 3171 692 3205 726 sw
rect 3258 692 3264 726
rect 3298 692 3337 726
tri 3478 724 3490 736 se
rect 3490 724 3976 736
tri 3450 696 3478 724 se
rect 3478 708 3936 724
rect 3478 696 3490 708
tri 3490 696 3502 708 nw
tri 2694 690 2696 692 se
rect 2696 690 2734 692
tri 2734 690 2736 692 nw
tri 3165 690 3167 692 ne
rect 3167 690 3205 692
tri 3205 690 3207 692 sw
rect 2240 656 2246 690
rect 2280 656 2286 690
tri 2693 689 2694 690 se
rect 2694 689 2733 690
tri 2733 689 2734 690 nw
tri 3167 689 3168 690 ne
rect 3168 689 3207 690
tri 3207 689 3208 690 sw
tri 2667 663 2693 689 se
rect 2693 687 2731 689
tri 2731 687 2733 689 nw
tri 3168 687 3170 689 ne
rect 3170 687 3208 689
rect 2693 663 2707 687
tri 2707 663 2731 687 nw
tri 2757 673 2771 687 se
rect 2771 673 3130 687
tri 3130 673 3144 687 sw
tri 3170 673 3184 687 ne
rect 3184 680 3208 687
tri 3208 680 3217 689 sw
rect 3258 680 3337 692
tri 3444 690 3450 696 se
rect 3450 690 3484 696
tri 3484 690 3490 696 nw
rect 3930 690 3936 708
rect 3970 690 3976 724
tri 3434 680 3444 690 se
rect 3444 680 3474 690
tri 3474 680 3484 690 nw
rect 3184 673 3217 680
tri 2747 663 2757 673 se
rect 2757 663 3144 673
tri 3144 663 3154 673 sw
tri 3184 663 3194 673 ne
rect 3194 663 3217 673
tri 2660 656 2667 663 se
rect 2667 656 2700 663
tri 2700 656 2707 663 nw
tri 2740 656 2747 663 se
rect 2747 659 3154 663
rect 2747 656 2780 659
tri 2780 656 2783 659 nw
tri 3118 656 3121 659 ne
rect 3121 656 3154 659
tri 3154 656 3161 663 sw
tri 3194 656 3201 663 ne
rect 3201 659 3217 663
tri 3217 659 3238 680 sw
tri 3413 659 3434 680 se
rect 3434 659 3453 680
tri 3453 659 3474 680 nw
tri 3493 659 3514 680 se
rect 3514 659 3832 680
rect 3201 656 3238 659
tri 3238 656 3241 659 sw
tri 3410 656 3413 659 se
rect 3413 656 3450 659
tri 3450 656 3453 659 nw
tri 3490 656 3493 659 se
rect 3493 656 3832 659
rect 2240 644 2286 656
tri 2654 650 2660 656 se
rect 2660 650 2694 656
tri 2694 650 2700 656 nw
tri 2734 650 2740 656 se
rect 2740 650 2771 656
rect 2327 649 2693 650
tri 2693 649 2694 650 nw
tri 2733 649 2734 650 se
rect 2734 649 2771 650
rect 2327 647 2691 649
tri 2691 647 2693 649 nw
tri 2731 647 2733 649 se
rect 2733 647 2771 649
tri 2771 647 2780 656 nw
tri 3121 647 3130 656 ne
rect 3130 650 3161 656
tri 3161 650 3167 656 sw
tri 3201 650 3207 656 ne
rect 3207 650 3241 656
rect 3130 649 3167 650
tri 3167 649 3168 650 sw
tri 3207 649 3208 650 ne
rect 3208 649 3241 650
tri 3241 649 3248 656 sw
tri 3403 649 3410 656 se
rect 3410 649 3443 656
tri 3443 649 3450 656 nw
tri 3483 649 3490 656 se
rect 3490 652 3714 656
rect 3490 649 3514 652
rect 3130 647 3168 649
rect 2153 600 2205 606
rect 2327 622 2666 647
tri 2666 622 2691 647 nw
tri 2717 633 2731 647 se
rect 2731 633 2757 647
tri 2757 633 2771 647 nw
tri 3130 633 3144 647 ne
rect 3144 633 3168 647
tri 3168 633 3184 649 sw
tri 3208 633 3224 649 ne
rect 3224 640 3434 649
tri 3434 640 3443 649 nw
tri 3474 640 3483 649 se
rect 3483 640 3514 649
tri 3514 640 3526 652 nw
rect 3224 633 3416 640
tri 2706 622 2717 633 se
rect 2717 622 2746 633
tri 2746 622 2757 633 nw
tri 3144 622 3155 633 ne
rect 3155 622 3184 633
tri 3184 622 3195 633 sw
tri 3224 622 3235 633 ne
rect 3235 622 3416 633
tri 3416 622 3434 640 nw
tri 3456 622 3474 640 se
rect 3474 622 3496 640
tri 3496 622 3514 640 nw
rect 3702 622 3714 652
rect 3748 622 3786 656
rect 3820 622 3832 656
rect 1796 573 1842 585
rect 1796 539 1802 573
rect 1836 539 1842 573
rect 1796 501 1842 539
rect 1796 467 1802 501
rect 1836 467 1842 501
rect 1796 434 1842 467
rect 2327 582 2373 622
tri 2702 618 2706 622 se
rect 2706 618 2742 622
tri 2742 618 2746 622 nw
tri 3155 618 3159 622 ne
rect 3159 621 3195 622
tri 3195 621 3196 622 sw
tri 3235 621 3236 622 ne
rect 3236 621 3415 622
tri 3415 621 3416 622 nw
tri 3455 621 3456 622 se
rect 3456 621 3492 622
rect 3159 618 3196 621
tri 3196 618 3199 621 sw
tri 3452 618 3455 621 se
rect 3455 618 3492 621
tri 3492 618 3496 622 nw
tri 2694 610 2702 618 se
rect 2702 610 2734 618
tri 2734 610 2742 618 nw
tri 3159 610 3167 618 ne
rect 3167 610 3199 618
tri 3199 610 3207 618 sw
tri 3444 610 3452 618 se
rect 3452 610 3484 618
tri 3484 610 3492 618 nw
rect 3702 616 3832 622
rect 3930 652 3976 690
rect 3930 618 3936 652
rect 3970 618 3976 652
tri 2691 607 2694 610 se
rect 2694 607 2731 610
tri 2731 607 2734 610 nw
tri 2682 598 2691 607 se
rect 2691 598 2722 607
tri 2722 598 2731 607 nw
rect 3002 598 3111 610
tri 3167 598 3179 610 ne
rect 3179 600 3207 610
tri 3207 600 3217 610 sw
tri 3434 600 3444 610 se
rect 3444 600 3474 610
tri 3474 600 3484 610 nw
rect 3179 598 3217 600
tri 3217 598 3219 600 sw
tri 3432 598 3434 600 se
rect 3434 598 3472 600
tri 3472 598 3474 600 nw
rect 3548 598 3594 610
rect 3930 606 3976 618
rect 4741 611 4747 663
rect 4799 611 4813 663
rect 4865 611 4871 663
rect 7804 607 7810 659
rect 7862 607 7880 659
rect 7932 607 7938 659
rect 2327 548 2333 582
rect 2367 548 2373 582
tri 2651 567 2682 598 se
rect 2682 567 2691 598
tri 2691 567 2722 598 nw
tri 2648 564 2651 567 se
rect 2651 564 2688 567
tri 2688 564 2691 567 nw
rect 3002 564 3071 598
rect 3105 564 3111 598
tri 3179 593 3184 598 ne
rect 3184 593 3219 598
tri 3219 593 3224 598 sw
tri 3427 593 3432 598 se
rect 3432 593 3467 598
tri 3467 593 3472 598 nw
tri 3111 574 3130 593 sw
tri 3184 574 3203 593 ne
rect 3203 574 3439 593
tri 3203 565 3212 574 ne
rect 3212 565 3439 574
tri 3439 565 3467 593 nw
rect 2327 510 2373 548
tri 2620 536 2648 564 se
rect 2648 536 2660 564
tri 2660 536 2688 564 nw
tri 2615 531 2620 536 se
rect 2620 531 2655 536
tri 2655 531 2660 536 nw
tri 2611 527 2615 531 se
rect 2615 527 2651 531
tri 2651 527 2655 531 nw
tri 2610 526 2611 527 se
rect 2611 526 2650 527
tri 2650 526 2651 527 nw
tri 2608 524 2610 526 se
rect 2610 524 2648 526
tri 2648 524 2650 526 nw
rect 2702 524 2748 536
rect 2327 476 2333 510
rect 2367 476 2373 510
tri 2574 490 2608 524 se
rect 2608 490 2614 524
tri 2614 490 2648 524 nw
rect 2702 490 2708 524
rect 2742 490 2748 524
tri 2571 487 2574 490 se
rect 2574 487 2611 490
tri 2611 487 2614 490 nw
rect 2327 464 2373 476
tri 2548 464 2571 487 se
rect 2571 464 2588 487
tri 2588 464 2611 487 nw
tri 2543 459 2548 464 se
rect 2548 459 2583 464
tri 2583 459 2588 464 nw
tri 2536 452 2543 459 se
rect 2543 452 2576 459
tri 2576 452 2583 459 nw
rect 2702 452 2748 490
rect 3002 526 3111 564
rect 3002 492 3071 526
rect 3105 492 3111 526
rect 3548 564 3554 598
rect 3588 564 3594 598
rect 4191 583 4237 595
rect 3548 526 3594 564
tri 3111 503 3130 522 nw
rect 3002 480 3111 492
rect 3548 492 3554 526
rect 3588 492 3594 526
rect 3548 480 3594 492
rect 3735 570 3782 582
rect 3735 536 3741 570
rect 3775 536 3782 570
rect 3735 498 3782 536
rect 3735 464 3741 498
rect 3775 464 3782 498
rect 3735 452 3782 464
rect 4021 575 4073 581
rect 4021 511 4073 523
rect 4191 549 4197 583
rect 4231 549 4237 583
rect 4191 511 4237 549
rect 8186 571 8238 577
rect 4191 477 4197 511
rect 4231 477 4237 511
tri 8152 503 8186 537 se
rect 8186 507 8238 519
rect 4191 465 4237 477
rect 4021 453 4073 459
tri 2531 447 2536 452 se
rect 2536 447 2571 452
tri 2571 447 2576 452 nw
tri 2518 434 2531 447 se
rect 2531 434 2558 447
tri 2558 434 2571 447 nw
rect 1796 418 2542 434
tri 2542 418 2558 434 nw
rect 2702 418 2708 452
rect 2742 418 3782 452
rect 4024 447 4070 453
rect 4752 451 4758 503
rect 4810 451 4822 503
rect 4874 451 4880 503
tri 8238 503 8272 537 sw
rect 8186 449 8238 455
rect 1796 406 2530 418
tri 2530 406 2542 418 nw
rect 2702 406 3782 418
rect -369 205 -317 211
tri -317 163 -275 205 sw
rect 2493 164 2499 374
rect 3433 163 4325 378
rect 4331 163 5080 378
tri 5325 341 5359 375 nw
tri 5080 163 5081 164 nw
rect -317 153 -275 163
rect -369 141 -275 153
rect -317 135 -275 141
tri -275 135 -247 163 sw
rect -317 89 878 135
rect -369 83 878 89
rect 930 83 942 135
rect 994 83 1000 135
tri 6461 22 6485 46 sw
rect 6433 16 6485 22
rect 6433 -48 6485 -36
rect 6433 -106 6485 -100
rect 6433 -158 6485 -152
rect 6433 -222 6485 -210
rect 6433 -280 6485 -274
tri 6461 -304 6485 -280 nw
<< via1 >>
rect 2723 3162 2775 3214
rect 2787 3162 2839 3214
rect 3113 3148 3165 3200
rect 3177 3148 3229 3200
rect 2485 3086 2537 3138
rect 2549 3086 2601 3138
rect 4867 3017 4919 3026
rect 4867 2983 4876 3017
rect 4876 2983 4910 3017
rect 4910 2983 4919 3017
rect 4867 2974 4919 2983
rect 4936 3017 4988 3026
rect 4936 2983 4948 3017
rect 4948 2983 4982 3017
rect 4982 2983 4988 3017
rect 4936 2974 4988 2983
rect 5032 3013 5084 3022
rect 5032 2979 5038 3013
rect 5038 2979 5072 3013
rect 5072 2979 5084 3013
rect 5032 2970 5084 2979
rect 5098 3013 5150 3022
rect 5098 2979 5110 3013
rect 5110 2979 5144 3013
rect 5144 2979 5150 3013
rect 5098 2970 5150 2979
rect 5207 3012 5259 3021
rect 5207 2978 5213 3012
rect 5213 2978 5247 3012
rect 5247 2978 5259 3012
rect 5207 2969 5259 2978
rect 5273 3012 5325 3021
rect 5273 2978 5285 3012
rect 5285 2978 5319 3012
rect 5319 2978 5325 3012
rect 5273 2969 5325 2978
rect 6132 3075 6184 3081
rect 6132 3041 6141 3075
rect 6141 3041 6175 3075
rect 6175 3041 6184 3075
rect 6132 3029 6184 3041
rect 6132 3003 6184 3015
rect 6132 2969 6141 3003
rect 6141 2969 6175 3003
rect 6175 2969 6184 3003
rect 6132 2963 6184 2969
rect 6278 3075 6330 3081
rect 6278 3041 6287 3075
rect 6287 3041 6321 3075
rect 6321 3041 6330 3075
rect 6278 3029 6330 3041
rect 6278 3003 6330 3015
rect 6278 2969 6287 3003
rect 6287 2969 6321 3003
rect 6321 2969 6330 3003
rect 6278 2963 6330 2969
rect 6432 3075 6484 3081
rect 6432 3041 6441 3075
rect 6441 3041 6475 3075
rect 6475 3041 6484 3075
rect 6432 3029 6484 3041
rect 6432 3003 6484 3015
rect 6432 2969 6441 3003
rect 6441 2969 6475 3003
rect 6475 2969 6484 3003
rect 6432 2963 6484 2969
rect 2566 2838 2618 2890
rect 2630 2838 2682 2890
rect 2980 2872 3032 2924
rect 3044 2872 3096 2924
rect 3469 2872 3521 2924
rect 3533 2872 3585 2924
rect 1220 2765 1272 2817
rect 1284 2765 1336 2817
rect 1425 2765 1477 2817
rect 1489 2765 1541 2817
rect 1861 2765 1913 2817
rect 1925 2765 1977 2817
rect 2057 2765 2109 2817
rect 2121 2765 2173 2817
rect 3247 2765 3299 2817
rect 3311 2765 3363 2817
rect 2447 2570 2461 2604
rect 2461 2570 2499 2604
rect 2447 2552 2499 2570
rect 2717 2572 2769 2578
rect 2447 2488 2499 2540
rect 2717 2538 2726 2572
rect 2726 2538 2760 2572
rect 2760 2538 2769 2572
rect 2717 2526 2769 2538
rect 2717 2495 2769 2507
rect 1390 2397 1442 2449
rect 1390 2358 1414 2385
rect 1414 2358 1442 2385
rect 1390 2333 1442 2358
rect 1470 2447 1522 2452
rect 1470 2413 1479 2447
rect 1479 2413 1513 2447
rect 1513 2413 1522 2447
rect 1470 2400 1522 2413
rect 1470 2373 1522 2385
rect 1470 2339 1479 2373
rect 1479 2339 1513 2373
rect 1513 2339 1522 2373
rect 1470 2333 1522 2339
rect 1574 2446 1626 2452
rect 1574 2412 1583 2446
rect 1583 2412 1617 2446
rect 1617 2412 1626 2446
rect 1574 2400 1626 2412
rect 1735 2430 1787 2453
rect 2717 2461 2726 2495
rect 2726 2461 2760 2495
rect 2760 2461 2769 2495
rect 4648 2555 4700 2607
rect 4712 2555 4764 2607
rect 2717 2455 2769 2461
rect 1735 2401 1764 2430
rect 1764 2401 1787 2430
rect 1574 2372 1626 2388
rect 1574 2338 1583 2372
rect 1583 2338 1617 2372
rect 1617 2338 1626 2372
rect 1574 2336 1626 2338
rect 1735 2335 1787 2387
rect 2912 2428 2964 2480
rect 3122 2453 3174 2505
rect 2912 2364 2964 2416
rect 3007 2438 3059 2444
rect 3007 2404 3016 2438
rect 3016 2404 3050 2438
rect 3050 2404 3059 2438
rect 3007 2392 3059 2404
rect 3122 2426 3174 2441
rect 3122 2392 3131 2426
rect 3131 2392 3165 2426
rect 3165 2392 3174 2426
rect 3122 2389 3174 2392
rect 3007 2365 3059 2377
rect 3007 2331 3016 2365
rect 3016 2331 3050 2365
rect 3050 2331 3059 2365
rect 3007 2325 3059 2331
rect 4073 2424 4125 2451
rect 4073 2399 4082 2424
rect 4082 2399 4116 2424
rect 4116 2399 4125 2424
rect 4073 2335 4125 2387
rect 1694 2189 1746 2241
rect 1758 2189 1810 2241
rect 3596 2239 3648 2291
rect 3596 2175 3648 2227
rect 3908 2218 3960 2270
rect 4468 2294 4520 2346
rect 4532 2323 4550 2346
rect 4550 2323 4584 2346
rect 4532 2294 4584 2323
rect 4835 2431 4887 2483
rect 4835 2367 4887 2419
rect 3908 2152 3960 2204
rect 2809 2099 2861 2151
rect 2873 2099 2925 2151
rect 1580 1893 1632 1945
rect 1644 1893 1696 1945
rect 3122 1884 3174 1936
rect 2429 1811 2481 1863
rect 2493 1811 2545 1863
rect 3122 1820 3174 1872
rect 3297 1828 3349 1855
rect 982 1755 1034 1759
rect 982 1721 989 1755
rect 989 1721 1023 1755
rect 1023 1721 1034 1755
rect 982 1707 1034 1721
rect 982 1683 1034 1695
rect 982 1649 989 1683
rect 989 1649 1023 1683
rect 1023 1649 1034 1683
rect 982 1643 1034 1649
rect 1580 1716 1632 1768
rect 2201 1749 2253 1801
rect 1580 1690 1632 1702
rect 1580 1656 1589 1690
rect 1589 1656 1623 1690
rect 1623 1656 1632 1690
rect 2201 1685 2253 1737
rect 2424 1723 2476 1775
rect 2424 1698 2476 1710
rect 2613 1731 2665 1783
rect 1580 1650 1632 1656
rect 2424 1664 2433 1698
rect 2433 1664 2467 1698
rect 2467 1664 2476 1698
rect 2424 1658 2476 1664
rect 2613 1701 2665 1719
rect 3297 1803 3307 1828
rect 3307 1803 3341 1828
rect 3341 1803 3349 1828
rect 4023 1893 4075 1945
rect 4087 1893 4139 1945
rect 2613 1667 2625 1701
rect 2625 1667 2659 1701
rect 2659 1667 2665 1701
rect 2985 1686 3037 1738
rect 3202 1728 3254 1780
rect 2985 1662 3037 1674
rect 2985 1628 2997 1662
rect 2997 1628 3031 1662
rect 3031 1628 3037 1662
rect 2985 1622 3037 1628
rect 3202 1664 3254 1716
rect 3297 1756 3349 1791
rect 3297 1739 3307 1756
rect 3307 1739 3341 1756
rect 3341 1739 3349 1756
rect 3425 1724 3477 1776
rect 3425 1660 3477 1712
rect 5876 1654 5928 1706
rect 5940 1654 5992 1706
rect 2153 1503 2205 1555
rect 2153 1439 2205 1491
rect 4403 1433 4455 1485
rect 4467 1433 4519 1485
rect 7700 1295 7752 1347
rect 7764 1295 7816 1347
rect 4919 1155 4971 1207
rect 4983 1155 5035 1207
rect 7049 1155 7101 1207
rect 7123 1155 7175 1207
rect 4747 1114 4799 1124
rect 4747 1080 4753 1114
rect 4753 1080 4787 1114
rect 4787 1080 4799 1114
rect 4747 1072 4799 1080
rect 4813 1114 4865 1124
rect 4813 1080 4825 1114
rect 4825 1080 4859 1114
rect 4859 1080 4865 1114
rect 4813 1072 4865 1080
rect 7809 1114 7861 1125
rect 7809 1080 7815 1114
rect 7815 1080 7849 1114
rect 7849 1080 7861 1114
rect 7809 1073 7861 1080
rect 7875 1114 7927 1125
rect 7875 1080 7887 1114
rect 7887 1080 7921 1114
rect 7921 1080 7927 1114
rect 7875 1073 7927 1080
rect 3788 912 3840 964
rect 3852 912 3904 964
rect 4747 959 4799 968
rect 4747 925 4753 959
rect 4753 925 4787 959
rect 4787 925 4799 959
rect 4747 916 4799 925
rect 4813 959 4865 968
rect 4813 925 4825 959
rect 4825 925 4859 959
rect 4859 925 4865 959
rect 4813 916 4865 925
rect 7809 959 7861 969
rect 7809 925 7815 959
rect 7815 925 7849 959
rect 7849 925 7861 959
rect 7809 917 7861 925
rect 7875 959 7927 969
rect 7875 925 7887 959
rect 7887 925 7921 959
rect 7921 925 7927 959
rect 7875 917 7927 925
rect 8229 839 8281 891
rect 1970 718 2022 722
rect 1970 684 1979 718
rect 1979 684 2013 718
rect 2013 684 2022 718
rect 1970 670 2022 684
rect 1970 646 2022 658
rect 1970 612 1979 646
rect 1979 612 2013 646
rect 2013 612 2022 646
rect 1970 606 2022 612
rect 2153 718 2205 722
rect 2153 684 2162 718
rect 2162 684 2196 718
rect 2196 684 2205 718
rect 2153 670 2205 684
rect 2153 646 2205 658
rect 2153 612 2162 646
rect 2162 612 2196 646
rect 2196 612 2205 646
rect 4747 809 4799 818
rect 4747 775 4753 809
rect 4753 775 4787 809
rect 4787 775 4799 809
rect 4747 766 4799 775
rect 4813 809 4865 818
rect 4813 775 4825 809
rect 4825 775 4859 809
rect 4859 775 4865 809
rect 4813 766 4865 775
rect 7804 809 7856 815
rect 7804 775 7810 809
rect 7810 775 7844 809
rect 7844 775 7856 809
rect 7804 763 7856 775
rect 7875 809 7927 815
rect 7875 775 7882 809
rect 7882 775 7916 809
rect 7916 775 7927 809
rect 7875 763 7927 775
rect 8229 775 8281 827
rect 2153 606 2205 612
rect 4747 653 4799 663
rect 4747 619 4753 653
rect 4753 619 4787 653
rect 4787 619 4799 653
rect 4747 611 4799 619
rect 4813 653 4865 663
rect 4813 619 4825 653
rect 4825 619 4859 653
rect 4859 619 4865 653
rect 4813 611 4865 619
rect 7810 653 7862 659
rect 7810 619 7816 653
rect 7816 619 7850 653
rect 7850 619 7862 653
rect 7810 607 7862 619
rect 7880 653 7932 659
rect 7880 619 7888 653
rect 7888 619 7922 653
rect 7922 619 7932 653
rect 7880 607 7932 619
rect 4021 565 4073 575
rect 4021 531 4030 565
rect 4030 531 4064 565
rect 4064 531 4073 565
rect 4021 523 4073 531
rect 4021 493 4073 511
rect 4021 459 4030 493
rect 4030 459 4064 493
rect 4064 459 4073 493
rect 8186 519 8238 571
rect 4758 451 4810 503
rect 4822 451 4874 503
rect 8186 455 8238 507
rect -369 153 -317 205
rect -369 89 -317 141
rect 878 83 930 135
rect 942 83 994 135
rect 6433 -36 6485 16
rect 6433 -100 6485 -48
rect 6433 -210 6485 -158
rect 6433 -274 6485 -222
<< metal2 >>
tri 1985 3324 2000 3339 se
rect 2000 3324 2442 3339
tri 2442 3324 2457 3339 sw
tri 1946 3285 1985 3324 se
rect 1985 3302 2457 3324
rect 1985 3285 2000 3302
tri 2000 3285 2017 3302 nw
tri 2405 3285 2422 3302 ne
rect 2422 3285 2457 3302
tri 1931 3270 1946 3285 se
rect 1946 3270 1985 3285
tri 1985 3270 2000 3285 nw
tri 2422 3270 2437 3285 ne
rect 2437 3270 2457 3285
tri 1346 2924 1377 2955 se
rect 1377 2924 1555 2955
tri 1555 2924 1586 2955 sw
tri 1312 2890 1346 2924 se
rect 1346 2903 1586 2924
rect 1346 2890 1386 2903
tri 1386 2890 1399 2903 nw
tri 1533 2890 1546 2903 ne
rect 1546 2890 1586 2903
tri 1586 2890 1620 2924 sw
tri 1304 2882 1312 2890 se
rect 1312 2882 1378 2890
tri 1378 2882 1386 2890 nw
tri 1546 2882 1554 2890 ne
rect 1554 2882 1620 2890
tri 1620 2882 1628 2890 sw
tri 1303 2881 1304 2882 se
rect 1304 2881 1377 2882
tri 1377 2881 1378 2882 nw
tri 1554 2881 1555 2882 ne
rect 1555 2881 1628 2882
tri 1273 2851 1303 2881 se
rect 1303 2851 1347 2881
tri 1347 2851 1377 2881 nw
tri 1555 2860 1576 2881 ne
tri 1260 2838 1273 2851 se
rect 1273 2838 1342 2851
tri 1342 2846 1347 2851 nw
tri 1239 2817 1260 2838 se
rect 1260 2817 1342 2838
rect 1214 2765 1220 2817
rect 1272 2765 1284 2817
rect 1336 2765 1342 2817
rect 1419 2765 1425 2817
rect 1477 2765 1489 2817
rect 1541 2765 1547 2817
tri 1398 2607 1419 2628 se
rect 1419 2607 1471 2765
tri 1471 2731 1505 2765 nw
tri 1566 2661 1576 2671 se
rect 1576 2661 1628 2881
tri 1918 2838 1931 2851 se
rect 1931 2838 1983 3270
tri 1983 3268 1985 3270 nw
tri 2437 3268 2439 3270 ne
rect 2439 3268 2457 3270
tri 2439 3250 2457 3268 ne
tri 2457 3250 2531 3324 sw
tri 2684 3283 2703 3302 se
rect 2703 3283 3238 3302
tri 3238 3283 3257 3302 sw
tri 2655 3254 2684 3283 se
rect 2684 3268 3257 3283
rect 2684 3254 2703 3268
tri 2703 3254 2717 3268 nw
tri 3224 3254 3238 3268 ne
rect 3238 3254 3257 3268
tri 2457 3228 2479 3250 ne
rect 2479 3162 2531 3250
tri 2654 3253 2655 3254 se
rect 2655 3253 2702 3254
tri 2702 3253 2703 3254 nw
tri 3238 3253 3239 3254 ne
rect 3239 3253 3257 3254
tri 2531 3162 2541 3172 sw
rect 2479 3148 2541 3162
tri 2541 3148 2555 3162 sw
rect 2479 3138 2555 3148
tri 2555 3138 2565 3148 sw
rect 2479 3086 2485 3138
rect 2537 3086 2549 3138
rect 2601 3086 2607 3138
tri 2653 2924 2654 2925 se
rect 2654 2924 2688 3253
tri 2688 3239 2702 3253 nw
tri 3239 3239 3253 3253 ne
rect 3253 3239 3257 3253
tri 3253 3235 3257 3239 ne
tri 3257 3235 3305 3283 sw
tri 3257 3225 3267 3235 ne
rect 3267 3225 3305 3235
tri 3267 3221 3271 3225 ne
tri 2619 2890 2653 2924 se
rect 2653 2890 2688 2924
rect 2560 2838 2566 2890
rect 2618 2838 2630 2890
rect 2682 2838 2688 2890
tri 1897 2817 1918 2838 se
rect 1918 2817 1983 2838
tri 2579 2817 2600 2838 ne
rect 2600 2817 2667 2838
tri 2667 2817 2688 2838 nw
rect 2717 3162 2723 3214
rect 2775 3162 2787 3214
rect 2839 3162 2845 3214
rect 2717 3148 2794 3162
tri 2794 3148 2808 3162 nw
rect 3107 3148 3113 3200
rect 3165 3148 3177 3200
rect 3229 3148 3235 3200
rect 1855 2765 1861 2817
rect 1913 2765 1925 2817
rect 1977 2765 1983 2817
rect 2051 2765 2057 2817
rect 2109 2765 2121 2817
rect 2173 2765 2179 2817
tri 2600 2804 2613 2817 ne
rect 2051 2728 2125 2765
tri 2125 2728 2162 2765 nw
tri 1512 2607 1566 2661 se
rect 1566 2610 1577 2661
tri 1577 2610 1628 2661 nw
tri 1977 2654 2051 2728 se
tri 2051 2654 2125 2728 nw
tri 1970 2647 1977 2654 se
rect 1977 2647 2044 2654
tri 2044 2647 2051 2654 nw
rect 1566 2607 1574 2610
tri 1574 2607 1577 2610 nw
tri 1395 2604 1398 2607 se
rect 1398 2606 1471 2607
rect 1398 2604 1469 2606
tri 1469 2604 1471 2606 nw
tri 1509 2604 1512 2607 se
rect 1512 2604 1571 2607
tri 1571 2604 1574 2607 nw
tri 1390 2599 1395 2604 se
rect 1395 2599 1464 2604
tri 1464 2599 1469 2604 nw
tri 1504 2599 1509 2604 se
rect 1509 2599 1566 2604
tri 1566 2599 1571 2604 nw
tri 1345 2554 1390 2599 se
rect 1390 2566 1431 2599
tri 1431 2566 1464 2599 nw
tri 1471 2566 1504 2599 se
rect 1504 2566 1519 2599
rect 1390 2554 1419 2566
tri 1419 2554 1431 2566 nw
tri 1459 2554 1471 2566 se
rect 1471 2554 1519 2566
tri 1343 2552 1345 2554 se
rect 1345 2552 1417 2554
tri 1417 2552 1419 2554 nw
tri 1457 2552 1459 2554 se
rect 1459 2552 1519 2554
tri 1519 2552 1566 2599 nw
tri 1331 2540 1343 2552 se
rect 1343 2540 1405 2552
tri 1405 2540 1417 2552 nw
tri 1445 2540 1457 2552 se
rect 1457 2540 1507 2552
tri 1507 2540 1519 2552 nw
tri 1328 2537 1331 2540 se
rect 1331 2537 1402 2540
tri 1402 2537 1405 2540 nw
tri 1442 2537 1445 2540 se
rect 1445 2537 1504 2540
tri 1504 2537 1507 2540 nw
tri 1279 2488 1328 2537 se
rect 1328 2514 1379 2537
tri 1379 2514 1402 2537 nw
tri 1419 2514 1442 2537 se
rect 1442 2514 1455 2537
rect 1328 2488 1353 2514
tri 1353 2488 1379 2514 nw
tri 1393 2488 1419 2514 se
rect 1419 2488 1455 2514
tri 1455 2488 1504 2537 nw
tri 1271 2480 1279 2488 se
rect 1279 2480 1345 2488
tri 1345 2480 1353 2488 nw
tri 1390 2485 1393 2488 se
rect 1393 2485 1449 2488
rect 1390 2482 1449 2485
tri 1449 2482 1455 2488 nw
tri 1246 2455 1271 2480 se
rect 1271 2455 1320 2480
tri 1320 2455 1345 2480 nw
tri 1244 2453 1246 2455 se
rect 1246 2453 1318 2455
tri 1318 2453 1320 2455 nw
tri 1243 2452 1244 2453 se
rect 1244 2452 1317 2453
tri 1317 2452 1318 2453 nw
tri 1240 2449 1243 2452 se
rect 1243 2449 1314 2452
tri 1314 2449 1317 2452 nw
rect 1390 2449 1442 2482
tri 1442 2475 1449 2482 nw
tri 1197 2406 1240 2449 se
rect 1240 2406 1271 2449
tri 1271 2406 1314 2449 nw
tri 1188 2397 1197 2406 se
rect 1197 2397 1262 2406
tri 1262 2397 1271 2406 nw
tri 1179 2388 1188 2397 se
rect 1188 2388 1253 2397
tri 1253 2388 1262 2397 nw
tri 1176 2385 1179 2388 se
rect 1179 2385 1250 2388
tri 1250 2385 1253 2388 nw
rect 1390 2385 1442 2397
tri 1160 2369 1176 2385 se
rect 1176 2369 1234 2385
tri 1234 2369 1250 2385 nw
tri 1152 2141 1160 2149 se
rect 1160 2141 1212 2369
tri 1212 2347 1234 2369 nw
rect 1390 2327 1442 2333
rect 1470 2452 1522 2458
rect 1470 2385 1522 2400
tri 1447 2152 1470 2175 se
rect 1470 2153 1522 2333
rect 1470 2152 1521 2153
tri 1521 2152 1522 2153 nw
rect 1574 2452 1626 2458
rect 1574 2388 1626 2400
tri 1446 2151 1447 2152 se
rect 1447 2151 1520 2152
tri 1520 2151 1521 2152 nw
tri 1436 2141 1446 2151 se
rect 1446 2141 1510 2151
tri 1510 2141 1520 2151 nw
tri 1110 2099 1152 2141 se
rect 1152 2127 1212 2141
tri 1264 2127 1278 2141 se
rect 1278 2127 1468 2141
rect 1152 2099 1184 2127
tri 1184 2099 1212 2127 nw
tri 1236 2099 1264 2127 se
rect 1264 2099 1468 2127
tri 1468 2099 1510 2141 nw
tri 1086 2075 1110 2099 se
rect 1110 2075 1160 2099
tri 1160 2075 1184 2099 nw
tri 1212 2075 1236 2099 se
rect 1236 2089 1458 2099
tri 1458 2089 1468 2099 nw
rect 1236 2075 1278 2089
tri 1078 2067 1086 2075 se
rect 1086 2067 1152 2075
tri 1152 2067 1160 2075 nw
tri 1204 2067 1212 2075 se
rect 1212 2067 1278 2075
tri 1278 2067 1300 2089 nw
tri 1012 2001 1078 2067 se
rect 1078 2023 1108 2067
tri 1108 2023 1152 2067 nw
tri 1160 2023 1204 2067 se
rect 1204 2023 1206 2067
rect 1078 2001 1086 2023
tri 1086 2001 1108 2023 nw
tri 1138 2001 1160 2023 se
rect 1160 2001 1206 2023
tri 982 1971 1012 2001 se
rect 1012 1971 1056 2001
tri 1056 1971 1086 2001 nw
tri 1132 1995 1138 2001 se
rect 1138 1995 1206 2001
tri 1206 1995 1278 2067 nw
rect 982 1759 1034 1971
tri 1034 1949 1056 1971 nw
rect 982 1695 1034 1707
rect 982 1637 1034 1643
tri 1068 1555 1132 1619 se
rect 1132 1597 1184 1995
tri 1184 1973 1206 1995 nw
rect 1574 1945 1626 2336
rect 1735 2453 1787 2459
rect 1735 2387 1787 2401
rect 1735 2241 1787 2335
rect 1688 2189 1694 2241
rect 1746 2189 1758 2241
rect 1810 2189 1816 2241
rect 1574 1893 1580 1945
rect 1632 1893 1644 1945
rect 1696 1893 1702 1945
rect 1132 1555 1142 1597
tri 1142 1555 1184 1597 nw
rect 1580 1768 1632 1774
rect 1580 1702 1632 1716
tri 1058 1545 1068 1555 se
rect 1068 1545 1132 1555
tri 1132 1545 1142 1555 nw
tri 1016 1503 1058 1545 se
rect 1058 1503 1113 1545
tri 1113 1526 1132 1545 nw
tri 1004 1491 1016 1503 se
rect 1016 1491 1113 1503
tri 998 1485 1004 1491 se
rect 1004 1485 1113 1491
rect 1580 247 1632 1650
rect 1970 722 2022 2647
tri 2022 2625 2044 2647 nw
rect 2447 2604 2499 2610
rect 2447 2540 2499 2552
tri 2444 1884 2447 1887 se
rect 2447 1884 2499 2488
tri 2499 1884 2512 1897 sw
tri 2432 1872 2444 1884 se
rect 2444 1872 2512 1884
tri 2512 1872 2524 1884 sw
tri 2423 1863 2432 1872 se
rect 2432 1863 2524 1872
tri 2524 1863 2533 1872 sw
rect 2197 1809 2253 1818
rect 2423 1811 2429 1863
rect 2481 1811 2493 1863
rect 2545 1811 2551 1863
rect 2613 1783 2665 2817
tri 2665 2815 2667 2817 nw
rect 2717 2578 2769 3148
tri 2769 3123 2794 3148 nw
tri 3107 3124 3131 3148 ne
rect 3131 3123 3210 3148
tri 3210 3123 3235 3148 nw
rect 2974 2872 2980 2924
rect 3032 2872 3044 2924
rect 3096 2872 3102 2924
rect 2974 2846 3076 2872
tri 3076 2846 3102 2872 nw
rect 2974 2809 3068 2846
tri 3068 2838 3076 2846 nw
rect 2974 2789 3048 2809
tri 3048 2789 3068 2809 nw
tri 2957 2772 2974 2789 se
rect 2974 2772 3031 2789
tri 3031 2772 3048 2789 nw
tri 2950 2765 2957 2772 se
rect 2957 2765 3024 2772
tri 3024 2765 3031 2772 nw
rect 2717 2507 2769 2526
rect 2717 2449 2769 2455
tri 2912 2727 2950 2765 se
rect 2950 2727 2986 2765
tri 2986 2727 3024 2765 nw
rect 2912 2480 2964 2727
tri 2964 2705 2986 2727 nw
rect 3131 2647 3183 3123
tri 3183 3096 3210 3123 nw
rect 3271 2970 3305 3225
rect 6132 3081 6184 3087
rect 4861 2974 4867 3026
rect 4919 2974 4936 3026
rect 4988 2974 4994 3026
tri 3305 2970 3307 2972 sw
rect 3271 2969 3307 2970
tri 3307 2969 3308 2970 sw
rect 3271 2968 3308 2969
tri 3308 2968 3309 2969 sw
rect 3271 2963 3309 2968
tri 3309 2963 3314 2968 sw
rect 3271 2958 3314 2963
tri 3271 2924 3305 2958 ne
rect 3305 2924 3314 2958
tri 3314 2924 3353 2963 sw
tri 3305 2920 3309 2924 ne
rect 3309 2920 3353 2924
tri 3353 2920 3357 2924 sw
tri 3309 2872 3357 2920 ne
tri 3357 2872 3405 2920 sw
rect 3463 2872 3469 2924
rect 3521 2872 3533 2924
rect 3585 2920 3998 2924
tri 3998 2920 4002 2924 sw
rect 3585 2872 4002 2920
tri 3357 2824 3405 2872 ne
tri 3405 2846 3431 2872 sw
tri 3976 2846 4002 2872 ne
tri 4002 2846 4076 2920 sw
rect 4920 2882 4972 2974
rect 5026 2970 5032 3022
rect 5084 2970 5098 3022
rect 5150 2970 5156 3022
rect 5026 2957 5156 2970
rect 5201 2969 5207 3021
rect 5259 2969 5273 3021
rect 5325 2969 5331 3021
rect 6132 3015 6184 3029
tri 5156 2957 5158 2959 sw
rect 6132 2957 6184 2963
rect 6278 3081 6330 3087
rect 6278 3015 6330 3029
rect 5026 2955 5158 2957
tri 5158 2955 5160 2957 sw
tri 5026 2924 5057 2955 ne
rect 5057 2952 5160 2955
tri 5160 2952 5163 2955 sw
rect 5057 2924 5163 2952
tri 5057 2920 5061 2924 ne
rect 5061 2922 5163 2924
tri 5163 2922 5193 2952 sw
tri 6248 2922 6278 2952 se
rect 6278 2922 6330 2963
rect 5061 2920 6330 2922
tri 5061 2904 5077 2920 ne
rect 5077 2908 6330 2920
rect 5077 2904 6294 2908
tri 4972 2882 4994 2904 sw
tri 5077 2882 5099 2904 ne
rect 5099 2882 6294 2904
tri 4920 2872 4930 2882 ne
rect 4930 2872 4994 2882
tri 4994 2872 5004 2882 sw
tri 5099 2872 5109 2882 ne
rect 5109 2872 6294 2882
tri 6294 2872 6330 2908 nw
rect 6432 3081 6484 3087
rect 6432 3015 6484 3029
tri 6410 2884 6432 2906 se
rect 6432 2884 6484 2963
tri 6398 2872 6410 2884 se
rect 6410 2872 6472 2884
tri 6472 2872 6484 2884 nw
tri 4930 2846 4956 2872 ne
rect 4956 2866 5004 2872
tri 5004 2866 5010 2872 sw
tri 6392 2866 6398 2872 se
rect 6398 2866 6466 2872
tri 6466 2866 6472 2872 nw
rect 4956 2846 5010 2866
rect 3405 2824 3431 2846
tri 3431 2824 3453 2846 sw
tri 4002 2824 4024 2846 ne
rect 4024 2824 4076 2846
tri 3405 2817 3412 2824 ne
rect 3412 2817 3958 2824
tri 3958 2817 3965 2824 sw
tri 4024 2817 4031 2824 ne
rect 4031 2817 4076 2824
rect 3241 2765 3247 2817
rect 3299 2765 3311 2817
rect 3363 2765 3369 2817
tri 3412 2790 3439 2817 ne
rect 3439 2790 3965 2817
tri 3944 2778 3956 2790 ne
rect 3956 2778 3965 2790
tri 3965 2778 4004 2817 sw
tri 4031 2778 4070 2817 ne
rect 4070 2778 4076 2817
tri 3956 2776 3958 2778 ne
rect 3958 2776 4004 2778
tri 3958 2765 3969 2776 ne
rect 3969 2772 4004 2776
tri 4004 2772 4010 2778 sw
tri 4070 2772 4076 2778 ne
tri 4076 2772 4150 2846 sw
tri 4956 2808 4994 2846 ne
rect 4994 2844 5010 2846
tri 5010 2844 5032 2866 sw
tri 6370 2844 6392 2866 se
rect 6392 2844 6408 2866
rect 4994 2808 6408 2844
tri 6408 2808 6466 2866 nw
tri 4994 2792 5010 2808 ne
rect 5010 2792 6392 2808
tri 6392 2792 6408 2808 nw
rect 3969 2765 4010 2772
tri 4010 2765 4017 2772 sw
tri 4076 2765 4083 2772 ne
rect 4083 2765 4150 2772
tri 3131 2607 3171 2647 ne
rect 3171 2607 3183 2647
tri 3183 2607 3245 2669 sw
tri 3171 2598 3180 2607 ne
rect 3180 2598 3245 2607
tri 3245 2598 3254 2607 sw
tri 3180 2595 3183 2598 ne
rect 3183 2595 3254 2598
tri 3183 2576 3202 2595 ne
rect 2912 2416 2964 2428
rect 2912 2358 2964 2364
rect 3007 2563 3063 2572
rect 3007 2483 3063 2507
rect 3059 2392 3063 2427
rect 3007 2377 3063 2392
rect 3059 2325 3063 2377
rect 3007 2319 3063 2325
rect 3122 2505 3174 2511
rect 3122 2441 3174 2453
rect 2803 2099 2809 2151
rect 2861 2099 2873 2151
rect 2925 2099 2931 2151
tri 2833 2058 2874 2099 ne
rect 2874 1967 2931 2099
tri 2874 1952 2889 1967 ne
rect 2889 1952 2931 1967
tri 2931 1952 2963 1984 sw
tri 2889 1945 2896 1952 ne
rect 2896 1945 2963 1952
tri 2963 1945 2970 1952 sw
tri 2896 1936 2905 1945 ne
rect 2905 1936 2970 1945
tri 2970 1936 2979 1945 sw
rect 3122 1936 3174 2389
tri 2905 1910 2931 1936 ne
rect 2931 1910 2979 1936
tri 2931 1884 2957 1910 ne
rect 2957 1884 2979 1910
tri 2979 1884 3031 1936 sw
tri 2957 1878 2963 1884 ne
rect 2963 1878 3031 1884
tri 3031 1878 3037 1884 sw
tri 2963 1872 2969 1878 ne
rect 2969 1872 3037 1878
tri 2969 1856 2985 1872 ne
rect 2197 1749 2201 1753
rect 2197 1737 2253 1749
rect 2197 1729 2201 1737
rect 2197 1664 2253 1673
rect 2424 1775 2480 1781
rect 2476 1772 2480 1775
rect 2424 1710 2480 1716
rect 2476 1692 2480 1710
rect 2613 1719 2665 1731
rect 2613 1661 2665 1667
rect 2985 1738 3037 1872
rect 3122 1872 3174 1884
rect 3122 1814 3174 1820
rect 2985 1674 3037 1686
rect 2424 1627 2480 1636
rect 3202 1780 3254 2595
tri 3297 1861 3308 1872 se
rect 3308 1861 3336 2765
tri 3969 2730 4004 2765 ne
rect 4004 2730 4017 2765
tri 4017 2730 4052 2765 sw
tri 4083 2730 4118 2765 ne
rect 4118 2730 4150 2765
tri 4004 2682 4052 2730 ne
tri 4052 2698 4084 2730 sw
tri 4118 2698 4150 2730 ne
tri 4150 2698 4224 2772 sw
rect 4052 2682 4084 2698
tri 4084 2682 4100 2698 sw
tri 4150 2682 4166 2698 ne
rect 4166 2682 4224 2698
tri 4052 2634 4100 2682 ne
tri 4100 2634 4148 2682 sw
tri 4166 2634 4214 2682 ne
rect 4214 2634 4224 2682
tri 4100 2607 4127 2634 ne
rect 4127 2624 4148 2634
tri 4148 2624 4158 2634 sw
tri 4214 2624 4224 2634 ne
tri 4224 2624 4298 2698 sw
rect 4127 2607 4158 2624
tri 4158 2607 4175 2624 sw
tri 4224 2607 4241 2624 ne
rect 4241 2607 4298 2624
tri 4298 2607 4315 2624 sw
tri 4127 2586 4148 2607 ne
rect 4148 2586 4175 2607
tri 4175 2586 4196 2607 sw
tri 4241 2586 4262 2607 ne
rect 4262 2586 4315 2607
tri 4148 2563 4171 2586 ne
rect 4171 2563 4196 2586
tri 4196 2563 4219 2586 sw
tri 4262 2563 4285 2586 ne
rect 4285 2563 4315 2586
rect 3529 2507 3538 2563
rect 3594 2507 3618 2563
rect 3674 2560 4127 2563
tri 4127 2560 4130 2563 sw
tri 4171 2560 4174 2563 ne
rect 4174 2560 4219 2563
tri 4219 2560 4222 2563 sw
tri 4285 2560 4288 2563 ne
rect 4288 2560 4315 2563
rect 3674 2555 4130 2560
tri 4130 2555 4135 2560 sw
tri 4174 2555 4179 2560 ne
rect 4179 2555 4222 2560
tri 4222 2555 4227 2560 sw
tri 4288 2555 4293 2560 ne
rect 4293 2555 4315 2560
tri 4315 2555 4367 2607 sw
rect 4642 2555 4648 2607
rect 4700 2555 4712 2607
rect 4764 2598 5978 2607
tri 5978 2598 5987 2607 sw
rect 4764 2555 5987 2598
rect 3674 2550 4135 2555
tri 4135 2550 4140 2555 sw
tri 4179 2550 4184 2555 ne
rect 4184 2550 4227 2555
tri 4227 2550 4232 2555 sw
tri 4293 2550 4298 2555 ne
rect 4298 2550 4367 2555
tri 4367 2550 4372 2555 sw
tri 5956 2550 5961 2555 ne
rect 5961 2550 5987 2555
tri 5987 2550 6035 2598 sw
rect 3674 2542 4140 2550
tri 4140 2542 4148 2550 sw
tri 4184 2542 4192 2550 ne
rect 4192 2542 4232 2550
rect 3674 2538 4148 2542
tri 4148 2538 4152 2542 sw
tri 4192 2538 4196 2542 ne
rect 4196 2538 4232 2542
tri 4232 2538 4244 2550 sw
tri 4298 2538 4310 2550 ne
rect 4310 2538 4372 2550
rect 3674 2511 4152 2538
tri 4152 2511 4179 2538 sw
tri 4196 2511 4223 2538 ne
rect 4223 2511 4244 2538
tri 4244 2511 4271 2538 sw
tri 4310 2511 4337 2538 ne
rect 4337 2511 4372 2538
tri 4372 2511 4411 2550 sw
tri 5961 2524 5987 2550 ne
rect 5987 2524 6035 2550
tri 6035 2524 6061 2550 sw
tri 5987 2511 6000 2524 ne
rect 6000 2511 6061 2524
tri 6061 2511 6074 2524 sw
rect 3674 2507 4179 2511
tri 4179 2507 4183 2511 sw
tri 4223 2507 4227 2511 ne
rect 4227 2507 4271 2511
tri 4271 2507 4275 2511 sw
tri 4337 2507 4341 2511 ne
rect 4341 2507 4411 2511
tri 4117 2494 4130 2507 ne
rect 4130 2494 4183 2507
tri 4183 2494 4196 2507 sw
tri 4227 2494 4240 2507 ne
rect 4240 2494 4275 2507
tri 4275 2494 4288 2507 sw
tri 4341 2494 4354 2507 ne
rect 4354 2494 4411 2507
tri 4130 2483 4141 2494 ne
rect 4141 2490 4196 2494
tri 4196 2490 4200 2494 sw
tri 4240 2490 4244 2494 ne
rect 4244 2490 4288 2494
tri 4288 2490 4292 2494 sw
tri 4354 2490 4358 2494 ne
rect 4358 2490 4411 2494
rect 4141 2483 4200 2490
tri 4200 2483 4207 2490 sw
tri 4244 2483 4251 2490 ne
rect 4251 2483 4292 2490
tri 4292 2483 4299 2490 sw
tri 4358 2483 4365 2490 ne
rect 4365 2489 4411 2490
tri 4411 2489 4433 2511 sw
tri 6000 2489 6022 2511 ne
rect 6022 2489 6074 2511
tri 6074 2489 6096 2511 sw
rect 4365 2483 4433 2489
tri 4433 2483 4439 2489 sw
tri 4829 2483 4835 2489 se
rect 4835 2483 4887 2489
tri 4141 2457 4167 2483 ne
rect 4167 2476 4207 2483
tri 4207 2476 4214 2483 sw
tri 4251 2476 4258 2483 ne
rect 4258 2476 4299 2483
tri 4299 2476 4306 2483 sw
tri 4365 2476 4372 2483 ne
rect 4372 2476 4439 2483
tri 4439 2476 4446 2483 sw
tri 4822 2476 4829 2483 se
rect 4829 2476 4835 2483
rect 4167 2457 4214 2476
tri 4214 2457 4233 2476 sw
tri 4258 2457 4277 2476 ne
rect 4277 2457 4306 2476
tri 4306 2457 4325 2476 sw
tri 4372 2457 4391 2476 ne
rect 4391 2457 4835 2476
rect 4073 2451 4125 2457
tri 4167 2431 4193 2457 ne
rect 4193 2446 4233 2457
tri 4233 2446 4244 2457 sw
tri 4277 2446 4288 2457 ne
rect 4288 2446 4325 2457
rect 4193 2442 4244 2446
tri 4244 2442 4248 2446 sw
tri 4288 2442 4292 2446 ne
rect 4292 2442 4325 2446
tri 4325 2442 4340 2457 sw
tri 4391 2442 4406 2457 ne
rect 4406 2442 4835 2457
rect 4193 2431 4248 2442
tri 4248 2431 4259 2442 sw
tri 4292 2431 4303 2442 ne
rect 4303 2431 4340 2442
tri 4340 2431 4351 2442 sw
tri 4406 2431 4417 2442 ne
rect 4417 2431 4835 2442
tri 6022 2450 6061 2489 ne
rect 6061 2450 6096 2489
tri 6096 2450 6135 2489 sw
tri 4193 2428 4196 2431 ne
rect 4196 2428 4259 2431
tri 4259 2428 4262 2431 sw
tri 4303 2428 4306 2431 ne
rect 4306 2428 4351 2431
tri 4351 2428 4354 2431 sw
tri 4417 2428 4420 2431 ne
rect 4420 2428 4887 2431
tri 4196 2419 4205 2428 ne
rect 4205 2424 4262 2428
tri 4262 2424 4266 2428 sw
tri 4306 2424 4310 2428 ne
rect 4310 2424 4354 2428
tri 4354 2424 4358 2428 sw
tri 4420 2424 4424 2428 ne
rect 4424 2424 4887 2428
rect 4205 2419 4266 2424
tri 4266 2419 4271 2424 sw
tri 4310 2419 4315 2424 ne
rect 4315 2419 4358 2424
tri 4358 2419 4363 2424 sw
tri 4801 2419 4806 2424 ne
rect 4806 2419 4887 2424
rect 3827 2388 3883 2397
rect 4073 2387 4125 2399
tri 3883 2335 3901 2353 sw
tri 4205 2367 4257 2419 ne
rect 4257 2398 4271 2419
tri 4271 2398 4292 2419 sw
tri 4315 2398 4336 2419 ne
rect 4336 2398 4363 2419
rect 4257 2394 4292 2398
tri 4292 2394 4296 2398 sw
tri 4336 2394 4340 2398 ne
rect 4340 2394 4363 2398
tri 4363 2394 4388 2419 sw
tri 4806 2394 4831 2419 ne
rect 4831 2394 4835 2419
rect 4257 2390 4296 2394
tri 4296 2390 4300 2394 sw
tri 4340 2390 4344 2394 ne
rect 4344 2390 4388 2394
tri 4388 2390 4392 2394 sw
tri 4831 2390 4835 2394 ne
rect 4257 2367 4300 2390
tri 4300 2367 4323 2390 sw
tri 4344 2367 4367 2390 ne
rect 4367 2367 4392 2390
tri 4392 2367 4415 2390 sw
tri 6061 2376 6135 2450 ne
tri 6135 2376 6209 2450 sw
tri 4257 2362 4262 2367 ne
rect 4262 2362 4323 2367
tri 4323 2362 4328 2367 sw
tri 4367 2362 4372 2367 ne
rect 4372 2362 4415 2367
tri 4415 2362 4420 2367 sw
tri 4262 2346 4278 2362 ne
rect 4278 2361 4328 2362
tri 4328 2361 4329 2362 sw
tri 4372 2361 4373 2362 ne
rect 4373 2361 4420 2362
tri 4420 2361 4421 2362 sw
rect 4835 2361 4887 2367
tri 6135 2361 6150 2376 ne
rect 6150 2361 6209 2376
tri 6209 2361 6224 2376 sw
rect 4278 2350 4329 2361
tri 4329 2350 4340 2361 sw
tri 4373 2350 4384 2361 ne
rect 4384 2350 4421 2361
rect 4278 2346 4340 2350
tri 4340 2346 4344 2350 sw
tri 4384 2346 4388 2350 ne
rect 4388 2346 4421 2350
tri 4421 2346 4436 2361 sw
tri 6150 2346 6165 2361 ne
rect 6165 2346 6224 2361
rect 3883 2332 3901 2335
rect 3827 2308 3901 2332
rect 3494 2241 3503 2297
rect 3559 2241 3583 2297
rect 3639 2291 3648 2297
tri 3546 2239 3548 2241 ne
rect 3548 2239 3596 2241
tri 3548 2227 3560 2239 ne
rect 3560 2227 3648 2239
tri 3560 2191 3596 2227 ne
rect 3596 2169 3648 2175
rect 3883 2294 3901 2308
tri 3901 2294 3942 2335 sw
rect 3883 2276 3942 2294
tri 3942 2276 3960 2294 sw
rect 3883 2270 3960 2276
rect 3883 2252 3908 2270
rect 3827 2218 3908 2252
rect 3827 2204 3960 2218
rect 3408 2113 3417 2169
rect 3473 2113 3497 2169
rect 3553 2113 3562 2169
rect 3827 2152 3908 2204
rect 3827 2146 3960 2152
tri 3408 2096 3425 2113 ne
rect 3425 2096 3545 2113
tri 3545 2096 3562 2113 nw
tri 3336 1861 3349 1874 sw
rect 3297 1855 3349 1861
rect 3297 1791 3349 1803
rect 3297 1733 3349 1739
rect 3425 1776 3477 2096
tri 3477 2028 3545 2096 nw
rect 4073 1945 4125 2335
tri 4278 2296 4328 2346 ne
rect 4328 2302 4344 2346
tri 4344 2302 4388 2346 sw
tri 4388 2312 4422 2346 ne
rect 4422 2312 4468 2346
tri 4444 2302 4454 2312 ne
rect 4454 2302 4468 2312
rect 4328 2296 4388 2302
tri 4388 2296 4394 2302 sw
tri 4454 2296 4460 2302 ne
rect 4460 2296 4468 2302
tri 4328 2294 4330 2296 ne
rect 4330 2294 4394 2296
tri 4394 2294 4396 2296 sw
tri 4460 2294 4462 2296 ne
rect 4462 2294 4468 2296
rect 4520 2294 4532 2346
rect 4584 2294 4590 2346
tri 6165 2302 6209 2346 ne
rect 6209 2302 6224 2346
tri 6224 2302 6283 2361 sw
tri 6209 2294 6217 2302 ne
rect 6217 2294 6283 2302
tri 4330 2230 4394 2294 ne
rect 4394 2280 4396 2294
tri 4396 2280 4410 2294 sw
tri 6217 2280 6231 2294 ne
rect 4394 2230 4410 2280
tri 4410 2230 4460 2280 sw
tri 4394 2174 4450 2230 ne
rect 4450 2174 6097 2230
tri 6075 2153 6096 2174 ne
rect 6096 2153 6097 2174
tri 6097 2153 6174 2230 sw
tri 6096 2152 6097 2153 ne
rect 6097 2152 6174 2153
tri 6097 2131 6118 2152 ne
rect 4017 1893 4023 1945
rect 4075 1893 4087 1945
rect 4139 1893 4145 1945
rect 3202 1716 3254 1728
rect 3202 1658 3254 1664
tri 3477 1733 3484 1740 sw
rect 3477 1724 3484 1733
rect 3425 1712 3484 1724
rect 3477 1706 3484 1712
tri 3484 1706 3511 1733 sw
rect 3477 1660 5876 1706
rect 3425 1654 5876 1660
rect 5928 1654 5940 1706
rect 5992 1654 5998 1706
rect 2985 1616 3037 1622
rect 1970 658 2022 670
rect 1970 600 2022 606
rect 2153 1555 2205 1561
rect 2153 1491 2205 1503
rect 2153 722 2205 1439
rect 4397 1433 4403 1485
rect 4455 1433 4467 1485
rect 4519 1461 4525 1485
tri 4525 1461 4549 1485 sw
rect 4519 1433 4948 1461
rect 2427 1385 2483 1394
rect 2427 1305 2483 1329
rect 2427 1207 2483 1249
tri 2483 1207 2497 1221 sw
rect 4920 1207 4948 1433
rect 6118 1363 6174 2152
rect 6231 1433 6283 2294
tri 6283 1433 6297 1447 sw
rect 6231 1425 6297 1433
tri 6231 1421 6235 1425 ne
rect 6235 1421 6297 1425
tri 6297 1421 6309 1433 sw
tri 6235 1373 6283 1421 ne
rect 6283 1373 6309 1421
tri 6283 1368 6288 1373 ne
rect 6288 1368 6309 1373
tri 6174 1363 6179 1368 sw
tri 6288 1363 6293 1368 ne
rect 6293 1363 6309 1368
rect 6118 1347 6179 1363
tri 6179 1347 6195 1363 sw
tri 6293 1347 6309 1363 ne
tri 6309 1347 6383 1421 sw
rect 6118 1346 6195 1347
tri 6118 1295 6169 1346 ne
rect 6169 1295 6195 1346
tri 6195 1295 6247 1347 sw
tri 6309 1295 6361 1347 ne
rect 6361 1295 7700 1347
rect 7752 1295 7764 1347
rect 7816 1295 7822 1347
tri 6169 1285 6179 1295 ne
rect 6179 1285 6247 1295
tri 6247 1285 6257 1295 sw
tri 6179 1207 6257 1285 ne
tri 6257 1207 6335 1285 sw
rect 2427 1199 2497 1207
tri 2427 1184 2442 1199 ne
rect 2442 1184 2497 1199
tri 2497 1184 2520 1207 sw
tri 2442 1155 2471 1184 ne
rect 2471 1155 2520 1184
tri 2520 1155 2549 1184 sw
rect 4913 1155 4919 1207
rect 4971 1155 4983 1207
rect 5035 1155 5041 1207
tri 6257 1155 6309 1207 ne
rect 6309 1155 7049 1207
rect 7101 1155 7123 1207
rect 7175 1155 7181 1207
tri 2471 1143 2483 1155 ne
rect 2483 1143 2549 1155
tri 2483 1125 2501 1143 ne
rect 2501 1125 2549 1143
tri 2549 1125 2579 1155 sw
tri 2501 1124 2502 1125 ne
rect 2502 1124 2579 1125
tri 2579 1124 2580 1125 sw
tri 7609 1124 7610 1125 se
rect 7610 1124 7809 1125
tri 2502 1106 2520 1124 ne
rect 2520 1106 2580 1124
tri 2580 1106 2598 1124 sw
tri 2520 1072 2554 1106 ne
rect 2554 1097 3213 1106
rect 2554 1072 3157 1097
tri 2554 1050 2576 1072 ne
rect 2576 1050 3157 1072
tri 3109 1002 3157 1050 ne
rect 4741 1072 4747 1124
rect 4799 1072 4813 1124
rect 4865 1073 7809 1124
rect 7861 1073 7875 1125
rect 7927 1073 7933 1125
rect 4865 1072 7631 1073
tri 7631 1072 7632 1073 nw
rect 3157 1017 3213 1041
tri 7489 968 7490 969 se
rect 7490 968 7809 969
rect 3157 952 3213 961
rect 3782 912 3788 964
rect 3840 912 3852 964
rect 3904 912 3910 964
rect 4741 916 4747 968
rect 4799 916 4813 968
rect 4865 917 7809 968
rect 7861 917 7875 969
rect 7927 917 7933 969
rect 4865 916 7623 917
tri 7623 916 7624 917 nw
rect 2153 658 2205 670
rect 2153 600 2205 606
rect 3858 553 3910 912
rect 8229 891 8281 897
rect 8229 827 8281 839
rect 4741 766 4747 818
rect 4799 766 4813 818
rect 4865 815 7615 818
tri 7615 815 7618 818 sw
rect 4865 766 7804 815
tri 7593 763 7596 766 ne
rect 7596 763 7804 766
rect 7856 763 7875 815
rect 7927 763 7933 815
rect 8229 696 8281 775
tri 8229 690 8235 696 ne
rect 8235 690 8281 696
tri 8281 690 8309 718 sw
tri 8235 663 8262 690 ne
rect 8262 663 8309 690
tri 8309 663 8336 690 sw
rect 4741 611 4747 663
rect 4799 611 4813 663
rect 4865 659 7687 663
tri 7687 659 7691 663 sw
tri 8262 659 8266 663 ne
rect 8266 659 8336 663
tri 8336 659 8340 663 sw
rect 4865 611 7810 659
tri 7665 607 7669 611 ne
rect 7669 607 7810 611
rect 7862 607 7880 659
rect 7932 607 7938 659
tri 8266 644 8281 659 ne
rect 8281 644 8340 659
tri 8281 616 8309 644 ne
rect 8309 616 8340 644
tri 8340 616 8383 659 sw
tri 8309 607 8318 616 ne
rect 8318 607 8578 616
tri 8578 607 8587 616 sw
tri 8318 591 8334 607 ne
rect 8334 591 8587 607
tri 8587 591 8603 607 sw
tri 8334 581 8344 591 ne
rect 8344 581 8603 591
tri 8603 581 8613 591 sw
rect 4021 575 4073 581
tri 8344 577 8348 581 ne
rect 8348 577 8613 581
tri 8613 577 8617 581 sw
rect 3858 523 4021 553
rect 3858 511 4073 523
rect 3858 501 4021 511
rect 8186 571 8238 577
tri 8348 564 8361 577 ne
rect 8361 564 8617 577
rect 8186 507 8238 519
tri 8556 517 8603 564 ne
rect 8603 517 8617 564
tri 8617 517 8677 577 sw
rect 4021 453 4073 459
rect 4752 451 4758 503
rect 4810 451 4822 503
rect 4874 451 4880 503
tri 8603 495 8625 517 ne
tri 8118 371 8186 439 se
rect 8186 417 8238 455
rect 8186 371 8192 417
tri 8192 371 8238 417 nw
rect 4128 308 4184 317
tri 1632 247 1641 256 sw
tri -341 211 -317 235 sw
rect -369 205 -317 211
rect 1580 213 1641 247
tri 1641 213 1675 247 sw
tri 4094 213 4128 247 se
rect 4128 228 4184 252
rect 1580 202 4128 213
tri 1580 161 1621 202 ne
rect 1621 172 4128 202
rect 1621 161 4184 172
rect -369 141 -317 153
rect -369 83 -317 89
tri -341 59 -317 83 nw
rect 872 83 878 135
rect 930 83 942 135
rect 994 83 1000 135
tri 872 59 896 83 ne
rect 896 59 970 83
tri 896 53 902 59 ne
rect 902 53 970 59
tri 970 53 1000 83 nw
tri 8108 53 8118 63 se
rect 8118 53 8170 371
tri 8170 349 8192 371 nw
tri 902 17 938 53 ne
rect 938 -80 970 53
tri 8104 49 8108 53 se
rect 8108 49 8170 53
rect 3157 40 3213 49
tri 3213 16 3246 49 sw
tri 8077 22 8104 49 se
rect 8104 41 8170 49
rect 8104 22 8118 41
rect 6433 16 6485 22
tri 8073 18 8077 22 se
rect 8077 18 8118 22
rect 3213 -16 3246 16
rect 3157 -34 3246 -16
tri 3246 -34 3296 16 sw
rect 3157 -36 5865 -34
tri 5865 -36 5867 -34 sw
tri 6485 -11 6514 18 sw
tri 8044 -11 8073 18 se
rect 8073 -11 8118 18
tri 8118 -11 8170 41 nw
tri 8571 -11 8625 43 se
rect 8625 21 8677 517
rect 6485 -16 6514 -11
tri 6514 -16 6519 -11 sw
tri 8039 -16 8044 -11 se
rect 8044 -16 8113 -11
tri 8113 -16 8118 -11 nw
tri 8566 -16 8571 -11 se
rect 8571 -16 8625 -11
rect 6485 -34 8095 -16
tri 8095 -34 8113 -16 nw
tri 8551 -31 8566 -16 se
rect 8566 -31 8625 -16
tri 8625 -31 8677 21 nw
tri 8548 -34 8551 -31 se
rect 6485 -36 8063 -34
rect 3157 -40 5867 -36
tri 938 -100 958 -80 ne
rect 958 -100 970 -80
tri 970 -100 1004 -66 sw
rect 3213 -48 5867 -40
tri 5867 -48 5879 -36 sw
rect 6433 -48 8063 -36
rect 3213 -66 5879 -48
tri 5879 -66 5897 -48 sw
rect 3213 -86 5897 -66
rect 3213 -96 3219 -86
rect 3157 -99 3219 -96
tri 3219 -99 3232 -86 nw
tri 5843 -99 5856 -86 ne
rect 5856 -99 5897 -86
tri 5897 -99 5930 -66 sw
rect 3157 -100 3218 -99
tri 3218 -100 3219 -99 nw
tri 5856 -100 5857 -99 ne
rect 5857 -100 5930 -99
tri 5930 -100 5931 -99 sw
rect 6485 -66 8063 -48
tri 8063 -66 8095 -34 nw
tri 8516 -66 8548 -34 se
rect 8548 -66 8551 -34
rect 6485 -68 8061 -66
tri 8061 -68 8063 -66 nw
tri 8514 -68 8516 -66 se
rect 8516 -68 8551 -66
rect 6485 -99 6488 -68
tri 6488 -99 6519 -68 nw
tri 8483 -99 8514 -68 se
rect 8514 -99 8551 -68
tri 958 -102 960 -100 ne
rect 960 -102 1004 -100
tri 1004 -102 1006 -100 sw
rect 3157 -102 3216 -100
tri 3216 -102 3218 -100 nw
tri 5857 -102 5859 -100 ne
rect 5859 -102 5931 -100
tri 5931 -102 5933 -100 sw
tri 960 -112 970 -102 ne
rect 970 -112 1006 -102
tri 970 -148 1006 -112 ne
tri 1006 -148 1052 -102 sw
rect 3157 -105 3213 -102
tri 3213 -105 3216 -102 nw
tri 5859 -105 5862 -102 ne
rect 5862 -105 5933 -102
tri 5862 -108 5865 -105 ne
rect 5865 -108 5933 -105
tri 5865 -148 5905 -108 ne
rect 5905 -148 5933 -108
tri 5933 -148 5979 -102 sw
rect 6433 -106 6485 -100
tri 6485 -102 6488 -99 nw
tri 8480 -102 8483 -99 se
rect 8483 -102 8551 -99
tri 8477 -105 8480 -102 se
rect 8480 -105 8551 -102
tri 8551 -105 8625 -31 nw
tri 8476 -106 8477 -105 se
rect 8477 -106 8504 -105
tri 8434 -148 8476 -106 se
rect 8476 -148 8504 -106
tri 1006 -158 1016 -148 ne
rect 1016 -158 1052 -148
tri 1052 -158 1062 -148 sw
tri 5905 -158 5915 -148 ne
rect 5915 -158 5979 -148
tri 5979 -158 5989 -148 sw
tri 8430 -152 8434 -148 se
rect 8434 -152 8504 -148
tri 8504 -152 8551 -105 nw
rect 6433 -158 8483 -152
tri 1016 -194 1052 -158 ne
rect 1052 -194 1062 -158
tri 1062 -194 1098 -158 sw
tri 5915 -173 5930 -158 ne
rect 5930 -173 5989 -158
tri 5989 -173 6004 -158 sw
tri 5930 -194 5951 -173 ne
rect 5951 -194 6004 -173
tri 6004 -194 6025 -173 sw
tri 1052 -210 1068 -194 ne
rect 1068 -210 1098 -194
tri 1098 -210 1114 -194 sw
tri 5951 -210 5967 -194 ne
rect 5967 -210 6025 -194
tri 6025 -210 6041 -194 sw
rect 6485 -173 8483 -158
tri 8483 -173 8504 -152 nw
rect 6485 -194 8462 -173
tri 8462 -194 8483 -173 nw
rect 6485 -204 8452 -194
tri 8452 -204 8462 -194 nw
tri 1068 -222 1080 -210 ne
rect 1080 -222 1114 -210
tri 1114 -222 1126 -210 sw
tri 5967 -222 5979 -210 ne
rect 5979 -222 6041 -210
tri 6041 -222 6053 -210 sw
rect 6433 -222 6485 -210
tri 1080 -240 1098 -222 ne
rect 1098 -240 1126 -222
tri 1126 -240 1144 -222 sw
tri 5979 -240 5997 -222 ne
rect 5997 -240 6053 -222
tri 6053 -240 6071 -222 sw
tri 1098 -274 1132 -240 ne
rect 1132 -274 1144 -240
tri 1144 -274 1178 -240 sw
tri 5997 -247 6004 -240 ne
rect 6004 -247 6071 -240
tri 6071 -247 6078 -240 sw
tri 6004 -274 6031 -247 ne
rect 6031 -274 6078 -247
tri 6078 -274 6105 -247 sw
tri 6485 -238 6519 -204 nw
tri 1132 -286 1144 -274 ne
rect 1144 -286 1178 -274
tri 1178 -286 1190 -274 sw
tri 6031 -286 6043 -274 ne
rect 6043 -286 6105 -274
tri 6105 -286 6117 -274 sw
tri 1144 -300 1158 -286 ne
rect 1158 -300 1324 -286
tri 1324 -300 1338 -286 sw
tri 6043 -300 6057 -286 ne
rect 6057 -288 6117 -286
tri 6117 -288 6119 -286 sw
rect 6057 -300 6119 -288
tri 6119 -300 6131 -288 sw
tri 6421 -300 6433 -288 se
rect 6433 -300 6485 -274
tri 1158 -318 1176 -300 ne
rect 1176 -318 1338 -300
tri 1310 -346 1338 -318 ne
tri 1338 -346 1384 -300 sw
tri 6057 -321 6078 -300 ne
rect 6078 -321 6131 -300
tri 6131 -321 6152 -300 sw
tri 6400 -321 6421 -300 se
rect 6421 -310 6485 -300
rect 6421 -321 6474 -310
tri 6474 -321 6485 -310 nw
tri 6078 -346 6103 -321 ne
rect 6103 -346 6422 -321
tri 1338 -392 1384 -346 ne
tri 1384 -392 1430 -346 sw
tri 6103 -373 6130 -346 ne
rect 6130 -373 6422 -346
tri 6422 -373 6474 -321 nw
tri 1384 -438 1430 -392 ne
tri 1430 -438 1476 -392 sw
tri 1430 -484 1476 -438 ne
tri 1476 -484 1522 -438 sw
tri 1476 -530 1522 -484 ne
tri 1522 -530 1568 -484 sw
tri 1522 -576 1568 -530 ne
tri 1568 -576 1614 -530 sw
tri 1568 -622 1614 -576 ne
tri 1614 -622 1660 -576 sw
tri 1614 -668 1660 -622 ne
tri 1660 -668 1706 -622 sw
rect 2250 -645 2306 -636
tri 1660 -714 1706 -668 ne
tri 1706 -696 1734 -668 sw
rect 1706 -714 1734 -696
tri 1734 -714 1752 -696 sw
tri 2232 -714 2250 -696 se
rect 2250 -714 2306 -701
tri 1706 -760 1752 -714 ne
tri 1752 -760 1798 -714 sw
tri 2186 -760 2232 -714 se
rect 2232 -725 2306 -714
rect 2232 -760 2250 -725
tri 1752 -792 1784 -760 ne
rect 1784 -781 2250 -760
rect 1784 -792 2306 -781
<< via2 >>
rect 2197 1801 2253 1809
rect 2197 1753 2201 1801
rect 2201 1753 2253 1801
rect 3007 2507 3063 2563
rect 3007 2444 3063 2483
rect 3007 2427 3059 2444
rect 3059 2427 3063 2444
rect 2197 1685 2201 1729
rect 2201 1685 2253 1729
rect 2197 1673 2253 1685
rect 2424 1723 2476 1772
rect 2476 1723 2480 1772
rect 2424 1716 2480 1723
rect 2424 1658 2476 1692
rect 2476 1658 2480 1692
rect 2424 1636 2480 1658
rect 3538 2507 3594 2563
rect 3618 2507 3674 2563
rect 3827 2332 3883 2388
rect 3503 2241 3559 2297
rect 3583 2291 3639 2297
rect 3583 2241 3596 2291
rect 3596 2241 3639 2291
rect 3827 2252 3883 2308
rect 3417 2113 3473 2169
rect 3497 2113 3553 2169
rect 2427 1329 2483 1385
rect 2427 1249 2483 1305
rect 3157 1041 3213 1097
rect 3157 961 3213 1017
rect 4128 252 4184 308
rect 4128 172 4184 228
rect 3157 -16 3213 40
rect 3157 -96 3213 -40
rect 2250 -701 2306 -645
rect 2250 -781 2306 -725
<< metal3 >>
rect 3002 2563 3679 2568
rect 3002 2507 3007 2563
rect 3063 2507 3538 2563
rect 3594 2507 3618 2563
rect 3674 2507 3679 2563
rect 3002 2502 3679 2507
rect 3002 2483 3068 2502
rect 3002 2427 3007 2483
rect 3063 2427 3068 2483
tri 3068 2468 3102 2502 nw
rect 3002 2422 3068 2427
tri 3266 2422 3274 2430 se
rect 3274 2422 3888 2430
tri 3237 2393 3266 2422 se
rect 3266 2393 3888 2422
tri 3232 2388 3237 2393 se
rect 3237 2388 3888 2393
tri 3180 2336 3232 2388 se
rect 3232 2364 3827 2388
rect 3232 2336 3274 2364
tri 3274 2336 3302 2364 nw
tri 3778 2336 3806 2364 ne
rect 3806 2336 3827 2364
tri 3176 2332 3180 2336 se
rect 3180 2332 3270 2336
tri 3270 2332 3274 2336 nw
tri 3806 2332 3810 2336 ne
rect 3810 2332 3827 2336
rect 3883 2332 3888 2388
tri 3161 2317 3176 2332 se
rect 3176 2317 3255 2332
tri 3255 2317 3270 2332 nw
tri 3810 2320 3822 2332 ne
tri 2694 2308 2703 2317 se
rect 2703 2308 3246 2317
tri 3246 2308 3255 2317 nw
rect 3822 2308 3888 2332
tri 2688 2302 2694 2308 se
rect 2694 2302 3240 2308
tri 3240 2302 3246 2308 nw
tri 2683 2297 2688 2302 se
rect 2688 2297 3235 2302
tri 3235 2297 3240 2302 nw
rect 3498 2297 3648 2302
tri 2627 2241 2683 2297 se
rect 2683 2251 3189 2297
tri 3189 2251 3235 2297 nw
rect 2683 2241 2721 2251
tri 2721 2241 2731 2251 nw
rect 3498 2241 3503 2297
rect 3559 2241 3583 2297
rect 3639 2252 3648 2297
tri 3648 2252 3698 2302 sw
rect 3822 2252 3827 2308
rect 3883 2252 3888 2308
rect 3639 2241 3698 2252
tri 2622 2236 2627 2241 se
rect 2627 2236 2716 2241
tri 2716 2236 2721 2241 nw
rect 3498 2236 3698 2241
tri 2609 2223 2622 2236 se
rect 2622 2223 2703 2236
tri 2703 2223 2716 2236 nw
tri 3620 2223 3633 2236 ne
rect 3633 2223 3698 2236
tri 2560 2174 2609 2223 se
rect 2609 2174 2654 2223
tri 2654 2174 2703 2223 nw
tri 3633 2174 3682 2223 ne
rect 3682 2174 3698 2223
tri 3698 2174 3776 2252 sw
rect 3822 2247 3888 2252
tri 2555 2169 2560 2174 se
rect 2560 2169 2649 2174
tri 2649 2169 2654 2174 nw
tri 2928 2169 2933 2174 se
rect 2933 2169 3558 2174
tri 2515 2129 2555 2169 se
rect 2555 2129 2609 2169
tri 2609 2129 2649 2169 nw
tri 2888 2129 2928 2169 se
rect 2928 2129 3417 2169
tri 2499 2113 2515 2129 se
rect 2515 2113 2593 2129
tri 2593 2113 2609 2129 nw
tri 2872 2113 2888 2129 se
rect 2888 2113 3417 2129
rect 3473 2113 3497 2169
rect 3553 2113 3558 2169
tri 3682 2158 3698 2174 ne
rect 3698 2158 3776 2174
tri 3776 2158 3792 2174 sw
tri 2466 2080 2499 2113 se
rect 2499 2080 2560 2113
tri 2560 2080 2593 2113 nw
tri 2839 2080 2872 2113 se
rect 2872 2108 3558 2113
tri 3698 2108 3748 2158 ne
rect 3748 2108 3792 2158
tri 3792 2108 3842 2158 sw
rect 2872 2080 2933 2108
tri 2933 2080 2961 2108 nw
tri 3748 2080 3776 2108 ne
rect 3776 2080 3842 2108
tri 3842 2080 3870 2108 sw
tri 2421 2035 2466 2080 se
rect 2466 2035 2515 2080
tri 2515 2035 2560 2080 nw
tri 2794 2035 2839 2080 se
tri 2419 2033 2421 2035 se
rect 2421 2033 2513 2035
tri 2513 2033 2515 2035 nw
tri 2792 2033 2794 2035 se
rect 2794 2033 2839 2035
rect 2192 1809 2258 1814
rect 2192 1753 2197 1809
rect 2253 1753 2258 1809
rect 2192 1729 2258 1753
rect 2192 1673 2197 1729
rect 2253 1673 2258 1729
rect 2192 1636 2258 1673
rect 2419 1772 2485 2033
tri 2485 2005 2513 2033 nw
tri 2764 2005 2792 2033 se
rect 2792 2005 2839 2033
tri 2745 1986 2764 2005 se
rect 2764 1986 2839 2005
tri 2839 1986 2933 2080 nw
tri 3776 2064 3792 2080 ne
rect 3792 2064 3870 2080
tri 3870 2064 3886 2080 sw
tri 3792 2036 3820 2064 ne
tri 2651 1892 2745 1986 se
tri 2745 1892 2839 1986 nw
rect 2419 1716 2424 1772
rect 2480 1716 2485 1772
rect 2419 1692 2485 1716
tri 2258 1636 2272 1650 sw
rect 2419 1636 2424 1692
rect 2480 1636 2485 1692
rect 2192 1631 2272 1636
tri 2272 1631 2277 1636 sw
rect 2419 1631 2485 1636
tri 2560 1801 2651 1892 se
rect 2651 1801 2654 1892
tri 2654 1801 2745 1892 nw
rect 2192 1622 2277 1631
tri 2277 1622 2286 1631 sw
tri 2192 1528 2286 1622 ne
tri 2286 1528 2380 1622 sw
tri 2286 1434 2380 1528 ne
tri 2380 1486 2422 1528 sw
rect 2380 1434 2422 1486
tri 2422 1434 2474 1486 sw
tri 2380 1392 2422 1434 ne
rect 2422 1420 2474 1434
tri 2474 1420 2488 1434 sw
rect 2422 1385 2488 1420
rect 2422 1329 2427 1385
rect 2483 1329 2488 1385
rect 2422 1305 2488 1329
rect 2422 1249 2427 1305
rect 2483 1249 2488 1305
rect 2422 1244 2488 1249
tri 2466 534 2560 628 se
rect 2560 600 2626 1801
tri 2626 1773 2654 1801 nw
tri 2560 534 2626 600 nw
rect 3152 1097 3218 1102
rect 3152 1041 3157 1097
rect 3213 1041 3218 1097
rect 3152 1017 3218 1041
rect 3152 961 3157 1017
rect 3213 961 3218 1017
tri 2372 440 2466 534 se
tri 2466 440 2560 534 nw
tri 2278 346 2372 440 se
tri 2372 346 2466 440 nw
tri 2245 313 2278 346 se
rect 2278 313 2339 346
tri 2339 313 2372 346 nw
rect 2245 308 2334 313
tri 2334 308 2339 313 nw
rect 2245 -645 2311 308
tri 2311 285 2334 308 nw
rect 3152 40 3218 961
rect 3820 660 3886 2064
tri 3886 660 3907 681 sw
rect 3820 653 3907 660
tri 3820 566 3907 653 ne
tri 3907 566 4001 660 sw
tri 3907 472 4001 566 ne
tri 4001 472 4095 566 sw
tri 4001 378 4095 472 ne
tri 4095 378 4189 472 sw
tri 4095 350 4123 378 ne
rect 4123 308 4189 378
rect 4123 252 4128 308
rect 4184 252 4189 308
rect 4123 228 4189 252
rect 4123 172 4128 228
rect 4184 172 4189 228
rect 4123 167 4189 172
rect 3152 -16 3157 40
rect 3213 -16 3218 40
rect 3152 -40 3218 -16
rect 3152 -96 3157 -40
rect 3213 -96 3218 -40
rect 3152 -101 3218 -96
rect 2245 -701 2250 -645
rect 2306 -701 2311 -645
rect 2245 -725 2311 -701
rect 2245 -781 2250 -725
rect 2306 -781 2311 -725
rect 2245 -786 2311 -781
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_0
timestamp 1624884095
transform -1 0 2178 0 1 139
box -42 24 569 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_1
timestamp 1624884095
transform 1 0 1996 0 1 139
box -42 24 569 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_2
timestamp 1624884095
transform -1 0 3457 0 1 139
box -42 24 569 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_3
timestamp 1624884095
transform -1 0 2992 0 1 139
box -42 24 569 1116
use sky130_fd_io__gpiov2_amux_nand4  sky130_fd_io__gpiov2_amux_nand4_0
timestamp 1624884095
transform 1 0 5688 0 -1 3114
box -62 33 1000 1842
use sky130_fd_io__gpiov2_amux_nand4  sky130_fd_io__gpiov2_amux_nand4_1
timestamp 1624884095
transform -1 0 5746 0 -1 3114
box -62 33 1000 1842
use sky130_fd_io__gpiov2_amux_nand5  sky130_fd_io__gpiov2_amux_nand5_0
timestamp 1624884095
transform 0 1 4701 1 0 140
box -47 33 1089 1846
use sky130_fd_io__gpiov2_amux_nand5  sky130_fd_io__gpiov2_amux_nand5_1
timestamp 1624884095
transform 0 -1 8349 1 0 140
box -47 33 1089 1846
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_0
timestamp 1624884095
transform 1 0 3391 0 1 139
box 0 24 534 1116
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_1
timestamp 1624884095
transform -1 0 4396 0 1 139
box 0 24 534 1116
use sky130_fd_io__nor2_1  sky130_fd_io__nor2_1_0
timestamp 1624884095
transform 1 0 688 0 1 1356
box -38 -49 326 715
use sky130_fd_io__nor2_1  sky130_fd_io__nor2_1_1
timestamp 1624884095
transform 1 0 1360 0 1 1356
box -38 -49 326 715
use sky130_fd_io__nor2_1  sky130_fd_io__nor2_1_2
timestamp 1624884095
transform 1 0 2800 0 1 1356
box -38 -49 326 715
use sky130_fd_io__nor2_1  sky130_fd_io__nor2_1_3
timestamp 1624884095
transform 1 0 2224 0 1 1356
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_0
timestamp 1624884095
transform 1 0 2512 0 1 1356
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_1
timestamp 1624884095
transform -1 0 1936 0 1 1356
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_2
timestamp 1624884095
transform 1 0 976 0 1 1356
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_3
timestamp 1624884095
transform -1 0 3760 0 1 1356
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_4
timestamp 1624884095
transform -1 0 4048 0 1 1356
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_5
timestamp 1624884095
transform -1 0 3088 0 -1 2688
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_6
timestamp 1624884095
transform 1 0 1936 0 1 1356
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_7
timestamp 1624884095
transform 1 0 4336 0 -1 2688
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_8
timestamp 1624884095
transform 1 0 1264 0 -1 2688
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_9
timestamp 1624884095
transform 1 0 2512 0 -1 2688
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_10
timestamp 1624884095
transform -1 0 4048 0 -1 2688
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_11
timestamp 1624884095
transform -1 0 3760 0 -1 2688
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_12
timestamp 1624884095
transform 1 0 688 0 -1 2688
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_13
timestamp 1624884095
transform 1 0 400 0 -1 2688
box -38 -49 326 715
use sky130_fd_io__inv_1  sky130_fd_io__inv_1_14
timestamp 1624884095
transform 1 0 3088 0 1 1356
box -38 -49 326 715
use sky130_fd_io__nand2_1  sky130_fd_io__nand2_1_0
timestamp 1624884095
transform 1 0 2224 0 -1 2688
box -38 -49 326 715
use sky130_fd_io__nand2_1  sky130_fd_io__nand2_1_1
timestamp 1624884095
transform 1 0 976 0 -1 2688
box -38 -49 326 715
use sky130_fd_io__nand2_1  sky130_fd_io__nand2_1_2
timestamp 1624884095
transform 1 0 4048 0 -1 2688
box -38 -49 326 715
use sky130_fd_io__nand2_1  sky130_fd_io__nand2_1_3
timestamp 1624884095
transform 1 0 3088 0 -1 2688
box -38 -49 326 715
use sky130_fd_io__xor2_1  sky130_fd_io__xor2_1_0
timestamp 1624884095
transform 1 0 1552 0 -1 2688
box -38 -49 710 715
use sky130_fd_io__tap_1  sky130_fd_io__tap_1_0
timestamp 1624884095
transform 1 0 1264 0 1 1356
box -38 -49 134 715
use sky130_fd_io__tap_1  sky130_fd_io__tap_1_1
timestamp 1624884095
transform 1 0 3376 0 1 1356
box -38 -49 134 715
use sky130_fd_io__tap_1  sky130_fd_io__tap_1_2
timestamp 1624884095
transform 1 0 3376 0 -1 2688
box -38 -49 134 715
<< labels >>
flabel comment s 3093 2901 3093 2901 0 FreeSans 440 0 0 0 AMUXBUSB_ON_N
flabel metal1 s 1858 808 1886 836 3 FreeSans 280 90 0 0 NMIDA_ON_N
port 1 nsew
flabel metal1 s 2251 730 2279 758 3 FreeSans 280 0 0 0 D_B
port 2 nsew
flabel metal1 s 3075 495 3103 523 3 FreeSans 280 90 0 0 PGB_AMX_VDDA_H_N
port 3 nsew
flabel metal1 s 3270 712 3298 740 3 FreeSans 280 90 0 0 PGB_PAD_VDDIOQ_H_N
port 4 nsew
flabel metal1 s 2628 718 2656 746 3 FreeSans 280 90 0 0 PGA_AMX_VDDA_H_N
port 5 nsew
flabel metal1 s 2793 817 2821 845 3 FreeSans 280 90 0 0 PGA_PAD_VDDIOQ_H_N
port 6 nsew
flabel metal1 s 2601 2851 2629 2879 3 FreeSans 280 0 0 0 PD_ON
port 7 nsew
flabel metal1 s 2738 1771 2766 1799 3 FreeSans 280 0 0 0 PD_ON_N
port 8 nsew
flabel metal1 s 6448 -205 6476 -177 3 FreeSans 280 0 0 0 PU_ON
port 9 nsew
flabel metal1 s 1693 1453 1721 1481 3 FreeSans 280 90 0 0 PU_ON_N
port 10 nsew
flabel metal1 s 2729 2507 2757 2535 3 FreeSans 280 0 0 0 AMUXBUSB_ON
port 11 nsew
flabel metal1 s 2576 2369 2604 2397 3 FreeSans 280 0 0 0 AMUXBUSB_ON_N
port 12 nsew
flabel metal1 s 3986 1654 4014 1682 3 FreeSans 280 0 0 0 OUT
port 13 nsew
flabel metal1 s 1970 1675 1998 1703 3 FreeSans 280 0 0 0 ANALOG_EN
port 14 nsew
flabel metal1 s 3986 2341 4014 2369 3 FreeSans 280 0 0 0 ANALOG_POL
port 15 nsew
flabel metal1 s 434 2341 462 2369 3 FreeSans 280 0 0 0 ANALOG_SEL
port 16 nsew
flabel metal1 s 1476 2382 1504 2410 3 FreeSans 280 0 0 0 AMUXBUSA_ON
port 17 nsew
flabel metal1 s 218 2765 246 2793 3 FreeSans 280 0 0 0 AMUXBUSA_ON_N
port 18 nsew
flabel metal1 s 3602 2649 3630 2677 3 FreeSans 280 0 0 0 VSSD
port 19 nsew
flabel metal1 s 3602 2033 3630 2061 3 FreeSans 280 0 0 0 VCCD
port 20 nsew
flabel metal1 s 3602 1370 3630 1398 3 FreeSans 280 0 0 0 VSSD
port 19 nsew
flabel metal1 s 3495 275 3523 303 3 FreeSans 280 0 0 0 VSSD
port 19 nsew
flabel metal1 s 5233 1323 5261 1351 3 FreeSans 280 0 0 0 VCCD
port 20 nsew
flabel metal1 s 5606 2567 5634 2595 3 FreeSans 280 0 0 0 VSSD
port 19 nsew
flabel metal1 s 3464 1098 3492 1126 3 FreeSans 280 0 0 0 VCCD
port 20 nsew
flabel metal1 s 4208 501 4236 529 3 FreeSans 280 0 0 0 NGB_PAD_VSWITCH_H
port 21 nsew
flabel metal1 s 3552 501 3580 529 3 FreeSans 280 0 0 0 NGA_PAD_VSWITCH_H
port 22 nsew
flabel metal1 s 7861 774 7889 802 3 FreeSans 280 0 0 0 NGA_PAD_VSWITCH_H_N
port 23 nsew
flabel metal1 s 7851 618 7879 646 3 FreeSans 280 0 0 0 NGB_PAD_VSWITCH_H_N
port 24 nsew
flabel metal1 s 6136 2977 6164 3005 3 FreeSans 280 0 0 0 NMIDA_VCCD_N
port 25 nsew
flabel metal1 s 4928 2977 4956 3005 3 FreeSans 280 0 0 0 PU_VDDIOQ_H_N
port 26 nsew
flabel metal1 s 5084 2977 5112 3005 3 FreeSans 280 0 0 0 PD_VSWITCH_H_N
port 27 nsew
flabel metal1 s 5240 2977 5268 3005 3 FreeSans 280 0 0 0 D_B
port 2 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 13317602
string GDS_START 13249762
<< end >>
