* NGSPICE file created from ota.ext - technology: sky130A


* Top level circuit ota

X0 Vout D2 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u M=20
X1 D2 Vout sky130_fd_pr__cap_mim_m3_2 l=2.5e+07u w=2.5e+07u
X2 Ibias Ibias GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+06u l=1e+06u M=8
X3 D2 Vp D5 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+07u l=500000u M=8
X4 Vout Ibias GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+06u l=1e+06u M=16
X5 VDD D1 D2 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u M=4
X6 D5 Ibias GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=3e+06u l=1e+06u M=8
X7 D1 D1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u M=4
X8 D1 Vn D5 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+07u l=500000u M=8
C0 Vp D2 0.90fF
C1 D5 D1 12.93fF
C2 Vp Vn 0.76fF
C3 D5 Ibias 5.39fF
C4 D5 D2 13.43fF
C5 D2 D1 6.82fF
C6 D5 Vn 0.86fF
C7 Vn D1 0.95fF
C8 D5 VDD 0.02fF
C9 VDD D1 8.11fF
C10 Vout D5 6.66fF
C11 Vout D1 2.21fF
C12 VDD Ibias 0.04fF
C13 Vn D2 0.40fF
C14 VDD D2 13.04fF
C15 Vout Ibias 5.46fF
C16 Vout D2 60.06fF
C17 Vout VDD 26.82fF
C18 Vp D5 1.55fF
C19 Vp D1 0.46fF
C20 Ibias GND 24.85fF
C21 Vout GND 32.21fF
C22 D1 GND 1.22fF
C23 D2 GND 12.13fF
C24 D5 GND 9.87fF
C25 Vn GND 3.02fF
C26 Vp GND 3.97fF
C27 VDD GND 74.72fF
.end

