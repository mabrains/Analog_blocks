magic
tech sky130A
magscale 1 2
timestamp 1624883981
<< checkpaint >>
rect -1260 -1260 1924 2474
<< nwell >>
rect 0 0 664 1214
<< pmoslvt >>
rect 204 102 304 1112
rect 360 102 460 1112
<< pdiff >>
rect 148 1100 204 1112
rect 148 1066 159 1100
rect 193 1066 204 1100
rect 148 1032 204 1066
rect 148 998 159 1032
rect 193 998 204 1032
rect 148 964 204 998
rect 148 930 159 964
rect 193 930 204 964
rect 148 896 204 930
rect 148 862 159 896
rect 193 862 204 896
rect 148 828 204 862
rect 148 794 159 828
rect 193 794 204 828
rect 148 760 204 794
rect 148 726 159 760
rect 193 726 204 760
rect 148 692 204 726
rect 148 658 159 692
rect 193 658 204 692
rect 148 624 204 658
rect 148 590 159 624
rect 193 590 204 624
rect 148 556 204 590
rect 148 522 159 556
rect 193 522 204 556
rect 148 488 204 522
rect 148 454 159 488
rect 193 454 204 488
rect 148 420 204 454
rect 148 386 159 420
rect 193 386 204 420
rect 148 352 204 386
rect 148 318 159 352
rect 193 318 204 352
rect 148 284 204 318
rect 148 250 159 284
rect 193 250 204 284
rect 148 216 204 250
rect 148 182 159 216
rect 193 182 204 216
rect 148 148 204 182
rect 148 114 159 148
rect 193 114 204 148
rect 148 102 204 114
rect 304 1100 360 1112
rect 304 1066 315 1100
rect 349 1066 360 1100
rect 304 1032 360 1066
rect 304 998 315 1032
rect 349 998 360 1032
rect 304 964 360 998
rect 304 930 315 964
rect 349 930 360 964
rect 304 896 360 930
rect 304 862 315 896
rect 349 862 360 896
rect 304 828 360 862
rect 304 794 315 828
rect 349 794 360 828
rect 304 760 360 794
rect 304 726 315 760
rect 349 726 360 760
rect 304 692 360 726
rect 304 658 315 692
rect 349 658 360 692
rect 304 624 360 658
rect 304 590 315 624
rect 349 590 360 624
rect 304 556 360 590
rect 304 522 315 556
rect 349 522 360 556
rect 304 488 360 522
rect 304 454 315 488
rect 349 454 360 488
rect 304 420 360 454
rect 304 386 315 420
rect 349 386 360 420
rect 304 352 360 386
rect 304 318 315 352
rect 349 318 360 352
rect 304 284 360 318
rect 304 250 315 284
rect 349 250 360 284
rect 304 216 360 250
rect 304 182 315 216
rect 349 182 360 216
rect 304 148 360 182
rect 304 114 315 148
rect 349 114 360 148
rect 304 102 360 114
rect 460 1100 516 1112
rect 460 1066 471 1100
rect 505 1066 516 1100
rect 460 1032 516 1066
rect 460 998 471 1032
rect 505 998 516 1032
rect 460 964 516 998
rect 460 930 471 964
rect 505 930 516 964
rect 460 896 516 930
rect 460 862 471 896
rect 505 862 516 896
rect 460 828 516 862
rect 460 794 471 828
rect 505 794 516 828
rect 460 760 516 794
rect 460 726 471 760
rect 505 726 516 760
rect 460 692 516 726
rect 460 658 471 692
rect 505 658 516 692
rect 460 624 516 658
rect 460 590 471 624
rect 505 590 516 624
rect 460 556 516 590
rect 460 522 471 556
rect 505 522 516 556
rect 460 488 516 522
rect 460 454 471 488
rect 505 454 516 488
rect 460 420 516 454
rect 460 386 471 420
rect 505 386 516 420
rect 460 352 516 386
rect 460 318 471 352
rect 505 318 516 352
rect 460 284 516 318
rect 460 250 471 284
rect 505 250 516 284
rect 460 216 516 250
rect 460 182 471 216
rect 505 182 516 216
rect 460 148 516 182
rect 460 114 471 148
rect 505 114 516 148
rect 460 102 516 114
<< pdiffc >>
rect 159 1066 193 1100
rect 159 998 193 1032
rect 159 930 193 964
rect 159 862 193 896
rect 159 794 193 828
rect 159 726 193 760
rect 159 658 193 692
rect 159 590 193 624
rect 159 522 193 556
rect 159 454 193 488
rect 159 386 193 420
rect 159 318 193 352
rect 159 250 193 284
rect 159 182 193 216
rect 159 114 193 148
rect 315 1066 349 1100
rect 315 998 349 1032
rect 315 930 349 964
rect 315 862 349 896
rect 315 794 349 828
rect 315 726 349 760
rect 315 658 349 692
rect 315 590 349 624
rect 315 522 349 556
rect 315 454 349 488
rect 315 386 349 420
rect 315 318 349 352
rect 315 250 349 284
rect 315 182 349 216
rect 315 114 349 148
rect 471 1066 505 1100
rect 471 998 505 1032
rect 471 930 505 964
rect 471 862 505 896
rect 471 794 505 828
rect 471 726 505 760
rect 471 658 505 692
rect 471 590 505 624
rect 471 522 505 556
rect 471 454 505 488
rect 471 386 505 420
rect 471 318 505 352
rect 471 250 505 284
rect 471 182 505 216
rect 471 114 505 148
<< nsubdiff >>
rect 36 1066 94 1112
rect 36 1032 48 1066
rect 82 1032 94 1066
rect 36 998 94 1032
rect 36 964 48 998
rect 82 964 94 998
rect 36 930 94 964
rect 36 896 48 930
rect 82 896 94 930
rect 36 862 94 896
rect 36 828 48 862
rect 82 828 94 862
rect 36 794 94 828
rect 36 760 48 794
rect 82 760 94 794
rect 36 726 94 760
rect 36 692 48 726
rect 82 692 94 726
rect 36 658 94 692
rect 36 624 48 658
rect 82 624 94 658
rect 36 590 94 624
rect 36 556 48 590
rect 82 556 94 590
rect 36 522 94 556
rect 36 488 48 522
rect 82 488 94 522
rect 36 454 94 488
rect 36 420 48 454
rect 82 420 94 454
rect 36 386 94 420
rect 36 352 48 386
rect 82 352 94 386
rect 36 318 94 352
rect 36 284 48 318
rect 82 284 94 318
rect 36 250 94 284
rect 36 216 48 250
rect 82 216 94 250
rect 36 182 94 216
rect 36 148 48 182
rect 82 148 94 182
rect 36 102 94 148
rect 570 1066 628 1112
rect 570 1032 582 1066
rect 616 1032 628 1066
rect 570 998 628 1032
rect 570 964 582 998
rect 616 964 628 998
rect 570 930 628 964
rect 570 896 582 930
rect 616 896 628 930
rect 570 862 628 896
rect 570 828 582 862
rect 616 828 628 862
rect 570 794 628 828
rect 570 760 582 794
rect 616 760 628 794
rect 570 726 628 760
rect 570 692 582 726
rect 616 692 628 726
rect 570 658 628 692
rect 570 624 582 658
rect 616 624 628 658
rect 570 590 628 624
rect 570 556 582 590
rect 616 556 628 590
rect 570 522 628 556
rect 570 488 582 522
rect 616 488 628 522
rect 570 454 628 488
rect 570 420 582 454
rect 616 420 628 454
rect 570 386 628 420
rect 570 352 582 386
rect 616 352 628 386
rect 570 318 628 352
rect 570 284 582 318
rect 616 284 628 318
rect 570 250 628 284
rect 570 216 582 250
rect 616 216 628 250
rect 570 182 628 216
rect 570 148 582 182
rect 616 148 628 182
rect 570 102 628 148
<< nsubdiffcont >>
rect 48 1032 82 1066
rect 48 964 82 998
rect 48 896 82 930
rect 48 828 82 862
rect 48 760 82 794
rect 48 692 82 726
rect 48 624 82 658
rect 48 556 82 590
rect 48 488 82 522
rect 48 420 82 454
rect 48 352 82 386
rect 48 284 82 318
rect 48 216 82 250
rect 48 148 82 182
rect 582 1032 616 1066
rect 582 964 616 998
rect 582 896 616 930
rect 582 828 616 862
rect 582 760 616 794
rect 582 692 616 726
rect 582 624 616 658
rect 582 556 616 590
rect 582 488 616 522
rect 582 420 616 454
rect 582 352 616 386
rect 582 284 616 318
rect 582 216 616 250
rect 582 148 616 182
<< poly >>
rect 159 1194 505 1214
rect 159 1160 179 1194
rect 213 1160 247 1194
rect 281 1160 315 1194
rect 349 1160 383 1194
rect 417 1160 451 1194
rect 485 1160 505 1194
rect 159 1144 505 1160
rect 204 1112 304 1144
rect 360 1112 460 1144
rect 204 70 304 102
rect 360 70 460 102
rect 159 54 505 70
rect 159 20 179 54
rect 213 20 247 54
rect 281 20 315 54
rect 349 20 383 54
rect 417 20 451 54
rect 485 20 505 54
rect 159 0 505 20
<< polycont >>
rect 179 1160 213 1194
rect 247 1160 281 1194
rect 315 1160 349 1194
rect 383 1160 417 1194
rect 451 1160 485 1194
rect 179 20 213 54
rect 247 20 281 54
rect 315 20 349 54
rect 383 20 417 54
rect 451 20 485 54
<< locali >>
rect 159 1160 171 1194
rect 213 1160 243 1194
rect 281 1160 315 1194
rect 349 1160 383 1194
rect 421 1160 451 1194
rect 493 1160 505 1194
rect 159 1100 193 1116
rect 48 1020 82 1032
rect 48 948 82 964
rect 48 876 82 896
rect 48 804 82 828
rect 48 732 82 760
rect 48 660 82 692
rect 48 590 82 624
rect 48 522 82 554
rect 48 454 82 482
rect 48 386 82 410
rect 48 318 82 338
rect 48 250 82 266
rect 48 182 82 194
rect 159 1032 193 1058
rect 159 964 193 986
rect 159 896 193 914
rect 159 828 193 842
rect 159 760 193 770
rect 159 692 193 698
rect 159 624 193 626
rect 159 588 193 590
rect 159 516 193 522
rect 159 444 193 454
rect 159 372 193 386
rect 159 300 193 318
rect 159 228 193 250
rect 159 156 193 182
rect 159 98 193 114
rect 315 1100 349 1116
rect 315 1032 349 1058
rect 315 964 349 986
rect 315 896 349 914
rect 315 828 349 842
rect 315 760 349 770
rect 315 692 349 698
rect 315 624 349 626
rect 315 588 349 590
rect 315 516 349 522
rect 315 444 349 454
rect 315 372 349 386
rect 315 300 349 318
rect 315 228 349 250
rect 315 156 349 182
rect 315 98 349 114
rect 471 1100 505 1116
rect 471 1032 505 1058
rect 471 964 505 986
rect 471 896 505 914
rect 471 828 505 842
rect 471 760 505 770
rect 471 692 505 698
rect 471 624 505 626
rect 471 588 505 590
rect 471 516 505 522
rect 471 444 505 454
rect 471 372 505 386
rect 471 300 505 318
rect 471 228 505 250
rect 471 156 505 182
rect 582 1020 616 1032
rect 582 948 616 964
rect 582 876 616 896
rect 582 804 616 828
rect 582 732 616 760
rect 582 660 616 692
rect 582 590 616 624
rect 582 522 616 554
rect 582 454 616 482
rect 582 386 616 410
rect 582 318 616 338
rect 582 250 616 266
rect 582 182 616 194
rect 471 98 505 114
rect 159 20 171 54
rect 213 20 243 54
rect 281 20 315 54
rect 349 20 383 54
rect 421 20 451 54
rect 493 20 505 54
<< viali >>
rect 171 1160 179 1194
rect 179 1160 205 1194
rect 243 1160 247 1194
rect 247 1160 277 1194
rect 315 1160 349 1194
rect 387 1160 417 1194
rect 417 1160 421 1194
rect 459 1160 485 1194
rect 485 1160 493 1194
rect 48 1066 82 1092
rect 48 1058 82 1066
rect 48 998 82 1020
rect 48 986 82 998
rect 48 930 82 948
rect 48 914 82 930
rect 48 862 82 876
rect 48 842 82 862
rect 48 794 82 804
rect 48 770 82 794
rect 48 726 82 732
rect 48 698 82 726
rect 48 658 82 660
rect 48 626 82 658
rect 48 556 82 588
rect 48 554 82 556
rect 48 488 82 516
rect 48 482 82 488
rect 48 420 82 444
rect 48 410 82 420
rect 48 352 82 372
rect 48 338 82 352
rect 48 284 82 300
rect 48 266 82 284
rect 48 216 82 228
rect 48 194 82 216
rect 48 148 82 156
rect 48 122 82 148
rect 159 1066 193 1092
rect 159 1058 193 1066
rect 159 998 193 1020
rect 159 986 193 998
rect 159 930 193 948
rect 159 914 193 930
rect 159 862 193 876
rect 159 842 193 862
rect 159 794 193 804
rect 159 770 193 794
rect 159 726 193 732
rect 159 698 193 726
rect 159 658 193 660
rect 159 626 193 658
rect 159 556 193 588
rect 159 554 193 556
rect 159 488 193 516
rect 159 482 193 488
rect 159 420 193 444
rect 159 410 193 420
rect 159 352 193 372
rect 159 338 193 352
rect 159 284 193 300
rect 159 266 193 284
rect 159 216 193 228
rect 159 194 193 216
rect 159 148 193 156
rect 159 122 193 148
rect 315 1066 349 1092
rect 315 1058 349 1066
rect 315 998 349 1020
rect 315 986 349 998
rect 315 930 349 948
rect 315 914 349 930
rect 315 862 349 876
rect 315 842 349 862
rect 315 794 349 804
rect 315 770 349 794
rect 315 726 349 732
rect 315 698 349 726
rect 315 658 349 660
rect 315 626 349 658
rect 315 556 349 588
rect 315 554 349 556
rect 315 488 349 516
rect 315 482 349 488
rect 315 420 349 444
rect 315 410 349 420
rect 315 352 349 372
rect 315 338 349 352
rect 315 284 349 300
rect 315 266 349 284
rect 315 216 349 228
rect 315 194 349 216
rect 315 148 349 156
rect 315 122 349 148
rect 471 1066 505 1092
rect 471 1058 505 1066
rect 471 998 505 1020
rect 471 986 505 998
rect 471 930 505 948
rect 471 914 505 930
rect 471 862 505 876
rect 471 842 505 862
rect 471 794 505 804
rect 471 770 505 794
rect 471 726 505 732
rect 471 698 505 726
rect 471 658 505 660
rect 471 626 505 658
rect 471 556 505 588
rect 471 554 505 556
rect 471 488 505 516
rect 471 482 505 488
rect 471 420 505 444
rect 471 410 505 420
rect 471 352 505 372
rect 471 338 505 352
rect 471 284 505 300
rect 471 266 505 284
rect 471 216 505 228
rect 471 194 505 216
rect 471 148 505 156
rect 471 122 505 148
rect 582 1066 616 1092
rect 582 1058 616 1066
rect 582 998 616 1020
rect 582 986 616 998
rect 582 930 616 948
rect 582 914 616 930
rect 582 862 616 876
rect 582 842 616 862
rect 582 794 616 804
rect 582 770 616 794
rect 582 726 616 732
rect 582 698 616 726
rect 582 658 616 660
rect 582 626 616 658
rect 582 556 616 588
rect 582 554 616 556
rect 582 488 616 516
rect 582 482 616 488
rect 582 420 616 444
rect 582 410 616 420
rect 582 352 616 372
rect 582 338 616 352
rect 582 284 616 300
rect 582 266 616 284
rect 582 216 616 228
rect 582 194 616 216
rect 582 148 616 156
rect 582 122 616 148
rect 171 20 179 54
rect 179 20 205 54
rect 243 20 247 54
rect 247 20 277 54
rect 315 20 349 54
rect 387 20 417 54
rect 417 20 421 54
rect 459 20 485 54
rect 485 20 493 54
<< metal1 >>
rect 159 1194 505 1214
rect 159 1160 171 1194
rect 205 1160 243 1194
rect 277 1160 315 1194
rect 349 1160 387 1194
rect 421 1160 459 1194
rect 493 1160 505 1194
rect 159 1148 505 1160
rect 36 1092 94 1104
rect 36 1058 48 1092
rect 82 1058 94 1092
rect 36 1020 94 1058
rect 36 986 48 1020
rect 82 986 94 1020
rect 36 948 94 986
rect 36 914 48 948
rect 82 914 94 948
rect 36 876 94 914
rect 36 842 48 876
rect 82 842 94 876
rect 36 804 94 842
rect 36 770 48 804
rect 82 770 94 804
rect 36 732 94 770
rect 36 698 48 732
rect 82 698 94 732
rect 36 660 94 698
rect 36 626 48 660
rect 82 626 94 660
rect 36 588 94 626
rect 36 554 48 588
rect 82 554 94 588
rect 36 516 94 554
rect 36 482 48 516
rect 82 482 94 516
rect 36 444 94 482
rect 36 410 48 444
rect 82 410 94 444
rect 36 372 94 410
rect 36 338 48 372
rect 82 338 94 372
rect 36 300 94 338
rect 36 266 48 300
rect 82 266 94 300
rect 36 228 94 266
rect 36 194 48 228
rect 82 194 94 228
rect 36 156 94 194
rect 36 122 48 156
rect 82 122 94 156
rect 36 110 94 122
rect 150 1092 202 1104
rect 150 1058 159 1092
rect 193 1058 202 1092
rect 150 1020 202 1058
rect 150 986 159 1020
rect 193 986 202 1020
rect 150 948 202 986
rect 150 914 159 948
rect 193 914 202 948
rect 150 876 202 914
rect 150 842 159 876
rect 193 842 202 876
rect 150 804 202 842
rect 150 770 159 804
rect 193 770 202 804
rect 150 732 202 770
rect 150 698 159 732
rect 193 698 202 732
rect 150 660 202 698
rect 150 626 159 660
rect 193 626 202 660
rect 150 588 202 626
rect 150 554 159 588
rect 193 554 202 588
rect 150 552 202 554
rect 150 488 159 500
rect 193 488 202 500
rect 150 424 159 436
rect 193 424 202 436
rect 150 360 159 372
rect 193 360 202 372
rect 150 300 202 308
rect 150 296 159 300
rect 193 296 202 300
rect 150 232 202 244
rect 150 168 202 180
rect 150 110 202 116
rect 306 1098 358 1104
rect 306 1034 358 1046
rect 306 970 358 982
rect 306 914 315 918
rect 349 914 358 918
rect 306 906 358 914
rect 306 842 315 854
rect 349 842 358 854
rect 306 778 315 790
rect 349 778 358 790
rect 306 714 315 726
rect 349 714 358 726
rect 306 660 358 662
rect 306 626 315 660
rect 349 626 358 660
rect 306 588 358 626
rect 306 554 315 588
rect 349 554 358 588
rect 306 516 358 554
rect 306 482 315 516
rect 349 482 358 516
rect 306 444 358 482
rect 306 410 315 444
rect 349 410 358 444
rect 306 372 358 410
rect 306 338 315 372
rect 349 338 358 372
rect 306 300 358 338
rect 306 266 315 300
rect 349 266 358 300
rect 306 228 358 266
rect 306 194 315 228
rect 349 194 358 228
rect 306 156 358 194
rect 306 122 315 156
rect 349 122 358 156
rect 306 110 358 122
rect 462 1092 514 1104
rect 462 1058 471 1092
rect 505 1058 514 1092
rect 462 1020 514 1058
rect 462 986 471 1020
rect 505 986 514 1020
rect 462 948 514 986
rect 462 914 471 948
rect 505 914 514 948
rect 462 876 514 914
rect 462 842 471 876
rect 505 842 514 876
rect 462 804 514 842
rect 462 770 471 804
rect 505 770 514 804
rect 462 732 514 770
rect 462 698 471 732
rect 505 698 514 732
rect 462 660 514 698
rect 462 626 471 660
rect 505 626 514 660
rect 462 588 514 626
rect 462 554 471 588
rect 505 554 514 588
rect 462 552 514 554
rect 462 488 471 500
rect 505 488 514 500
rect 462 424 471 436
rect 505 424 514 436
rect 462 360 471 372
rect 505 360 514 372
rect 462 300 514 308
rect 462 296 471 300
rect 505 296 514 300
rect 462 232 514 244
rect 462 168 514 180
rect 462 110 514 116
rect 570 1092 628 1104
rect 570 1058 582 1092
rect 616 1058 628 1092
rect 570 1020 628 1058
rect 570 986 582 1020
rect 616 986 628 1020
rect 570 948 628 986
rect 570 914 582 948
rect 616 914 628 948
rect 570 876 628 914
rect 570 842 582 876
rect 616 842 628 876
rect 570 804 628 842
rect 570 770 582 804
rect 616 770 628 804
rect 570 732 628 770
rect 570 698 582 732
rect 616 698 628 732
rect 570 660 628 698
rect 570 626 582 660
rect 616 626 628 660
rect 570 588 628 626
rect 570 554 582 588
rect 616 554 628 588
rect 570 516 628 554
rect 570 482 582 516
rect 616 482 628 516
rect 570 444 628 482
rect 570 410 582 444
rect 616 410 628 444
rect 570 372 628 410
rect 570 338 582 372
rect 616 338 628 372
rect 570 300 628 338
rect 570 266 582 300
rect 616 266 628 300
rect 570 228 628 266
rect 570 194 582 228
rect 616 194 628 228
rect 570 156 628 194
rect 570 122 582 156
rect 616 122 628 156
rect 570 110 628 122
rect 159 54 505 66
rect 159 20 171 54
rect 205 20 243 54
rect 277 20 315 54
rect 349 20 387 54
rect 421 20 459 54
rect 493 20 505 54
rect 159 0 505 20
<< via1 >>
rect 150 516 202 552
rect 150 500 159 516
rect 159 500 193 516
rect 193 500 202 516
rect 150 482 159 488
rect 159 482 193 488
rect 193 482 202 488
rect 150 444 202 482
rect 150 436 159 444
rect 159 436 193 444
rect 193 436 202 444
rect 150 410 159 424
rect 159 410 193 424
rect 193 410 202 424
rect 150 372 202 410
rect 150 338 159 360
rect 159 338 193 360
rect 193 338 202 360
rect 150 308 202 338
rect 150 266 159 296
rect 159 266 193 296
rect 193 266 202 296
rect 150 244 202 266
rect 150 228 202 232
rect 150 194 159 228
rect 159 194 193 228
rect 193 194 202 228
rect 150 180 202 194
rect 150 156 202 168
rect 150 122 159 156
rect 159 122 193 156
rect 193 122 202 156
rect 150 116 202 122
rect 306 1092 358 1098
rect 306 1058 315 1092
rect 315 1058 349 1092
rect 349 1058 358 1092
rect 306 1046 358 1058
rect 306 1020 358 1034
rect 306 986 315 1020
rect 315 986 349 1020
rect 349 986 358 1020
rect 306 982 358 986
rect 306 948 358 970
rect 306 918 315 948
rect 315 918 349 948
rect 349 918 358 948
rect 306 876 358 906
rect 306 854 315 876
rect 315 854 349 876
rect 349 854 358 876
rect 306 804 358 842
rect 306 790 315 804
rect 315 790 349 804
rect 349 790 358 804
rect 306 770 315 778
rect 315 770 349 778
rect 349 770 358 778
rect 306 732 358 770
rect 306 726 315 732
rect 315 726 349 732
rect 349 726 358 732
rect 306 698 315 714
rect 315 698 349 714
rect 349 698 358 714
rect 306 662 358 698
rect 462 516 514 552
rect 462 500 471 516
rect 471 500 505 516
rect 505 500 514 516
rect 462 482 471 488
rect 471 482 505 488
rect 505 482 514 488
rect 462 444 514 482
rect 462 436 471 444
rect 471 436 505 444
rect 505 436 514 444
rect 462 410 471 424
rect 471 410 505 424
rect 505 410 514 424
rect 462 372 514 410
rect 462 338 471 360
rect 471 338 505 360
rect 505 338 514 360
rect 462 308 514 338
rect 462 266 471 296
rect 471 266 505 296
rect 505 266 514 296
rect 462 244 514 266
rect 462 228 514 232
rect 462 194 471 228
rect 471 194 505 228
rect 505 194 514 228
rect 462 180 514 194
rect 462 156 514 168
rect 462 122 471 156
rect 471 122 505 156
rect 505 122 514 156
rect 462 116 514 122
<< metal2 >>
rect 10 1098 654 1104
rect 10 1046 306 1098
rect 358 1046 654 1098
rect 10 1034 654 1046
rect 10 982 306 1034
rect 358 982 654 1034
rect 10 970 654 982
rect 10 918 306 970
rect 358 918 654 970
rect 10 906 654 918
rect 10 854 306 906
rect 358 854 654 906
rect 10 842 654 854
rect 10 790 306 842
rect 358 790 654 842
rect 10 778 654 790
rect 10 726 306 778
rect 358 726 654 778
rect 10 714 654 726
rect 10 662 306 714
rect 358 662 654 714
rect 10 632 654 662
rect 10 552 654 582
rect 10 500 150 552
rect 202 500 462 552
rect 514 500 654 552
rect 10 488 654 500
rect 10 436 150 488
rect 202 436 462 488
rect 514 436 654 488
rect 10 424 654 436
rect 10 372 150 424
rect 202 372 462 424
rect 514 372 654 424
rect 10 360 654 372
rect 10 308 150 360
rect 202 308 462 360
rect 514 308 654 360
rect 10 296 654 308
rect 10 244 150 296
rect 202 244 462 296
rect 514 244 654 296
rect 10 232 654 244
rect 10 180 150 232
rect 202 180 462 232
rect 514 180 654 232
rect 10 168 654 180
rect 10 116 150 168
rect 202 116 462 168
rect 514 116 654 168
rect 10 110 654 116
<< labels >>
flabel metal2 s 16 757 35 827 0 FreeSans 400 90 0 0 DRAIN
port 2 nsew
flabel metal2 s 14 320 35 384 0 FreeSans 400 90 0 0 SOURCE
port 4 nsew
flabel metal1 s 159 1148 505 1214 0 FreeSans 300 0 0 0 GATE
port 3 nsew
flabel metal1 s 159 0 505 66 0 FreeSans 300 0 0 0 GATE
port 3 nsew
flabel metal1 s 56 732 56 732 7 FreeSans 400 90 0 0 BULK
port 1 nsew
flabel metal1 s 598 732 598 732 7 FreeSans 400 90 0 0 BULK
port 1 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 9989442
string GDS_START 9973406
<< end >>
