
.include ~/mabrains/Analog_blocks/Analog_Blocks/Bandgap/Netlists/Design/BGR_5v/Bandgap_self_3.3v.spice
*Supply Variation
.control
dc Vs 0 6 0.3
plot vdd bg_out
meas DC Vref_Sup_pos10per FIND bg_out AT=3
meas DC Vref_Sup_neg10per FIND bg_out AT=3.6
.endc
*Temprature Variation
.control
alter Vs DC = 3.3
dc temp -40 125 1
plot v(bg_out)
.endc

*PSRR Analysis
.control
alter Vs DC =3.3
alter Vs AC = 1
ac dec 10 1 1G
plot db(bg_out)
meas ac PSRR_1k FIND vdb(bg_out) AT=1k
meas ac PSRR_1M FIND vdb(bg_out) AT=1Meg
.endc
.op
**Transient
.control
alter @Vs[pwl] = [ 0 0 5u 0 15u 3.6 25u 3.6 ]
tran 1u 20u
plot vdd bg_out
.endc

