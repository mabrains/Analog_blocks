**** begin user architecture code
.nodeset v(inn)=1.1
.nodeset v(inp)=1.1
.nodeset v(mir)=0.9
.nodeset v(bg_out)=1.2
.nodeset v(ldo_out)=1.8
.nodeset v(pos)=1.2

*OP_Simulation
.control
op
print all
.endc

.control
dc Vs 2.5 0 -0.02
plot vdd ldo_out
meas DC Vref_Sup_pos10per FIND bg_out AT=2
meas DC Vref_Sup_neg10per FIND bg_out AT=2.4
.endc

*Temprature Variation
.control
let i=16
dc temp 85 0 -1
set appendwrite
write temp_var_ldo.raw
load temp_var_ldo.raw
plot v (ldo_out)
.endc



*Psrr_Simulation
.control
alter Vs AC =1
ac dec 10 1 1G
plot vdb (ldo_out)
let psrr = vdb(ldo_out)
meas ac PSRR_1k FIND vdb(ldo_out) AT=1k
meas ac PSRR_1M FIND vdb(ldo_out) AT=100k
set appendwrite
write psrr_ldo.raw
load psrr_ldo.raw
quit
.endc

*Transient
.control
alter @Vs[pulse] = [ 0 2 15u 1u 5u 100u 200u ]
tran 0.1u 100u
plot vdd ldo_out
.endc
.control
alter @Vs[pulse] = [ 0 2.2 15u 1u 5u 100u 200u ]
tran 0.1u 100u
plot vdd ldo_out
.endc
.control
alter @Vs[pulse] = [ 0 2.4 15u 1u 5u 100u 200u ]
tran 0.1u 100u
plot vdd ldo_out
.endc


**** end user architecture code
**.ends
.GLOBAL VDD
.GLOBAL GND
** flattened .save nodes
.end
