magic
tech sky130A
magscale 1 2
timestamp 1624884095
<< checkpaint >>
rect -524 2324 11010 40722
<< metal3 >>
rect 736 39434 2728 39446
rect 736 36730 780 39434
rect 2684 36730 2728 39434
rect 736 36718 2728 36730
rect 2908 39431 4894 39452
rect 2908 34887 2949 39431
rect 4853 34887 4894 39431
rect 2908 34866 4894 34887
rect 5280 39441 7266 39462
rect 5280 34897 5321 39441
rect 7225 34897 7266 39441
rect 5280 34876 7266 34897
rect 7624 18529 9746 18550
rect 7624 13665 7653 18529
rect 9717 13665 9746 18529
rect 7624 13644 9746 13665
rect 5216 5618 7336 5660
rect 5216 4834 5244 5618
rect 7308 4834 7336 5618
rect 5216 4792 7336 4834
rect 7604 4409 9750 4450
rect 7604 3625 7645 4409
rect 9709 3625 9750 4409
rect 7604 3584 9750 3625
<< via3 >>
rect 780 36730 2684 39434
rect 2949 34887 4853 39431
rect 5321 34897 7225 39441
rect 7653 13665 9717 18529
rect 5244 4834 7308 5618
rect 7645 3625 9709 4409
<< metal4 >>
rect 736 39434 2728 39446
rect 736 36730 780 39434
rect 2684 36730 2728 39434
rect 736 36718 2728 36730
rect 2908 39431 4894 39452
rect 2908 34887 2949 39431
rect 4853 34887 4894 39431
rect 2908 34866 4894 34887
rect 5280 39441 7266 39462
rect 5280 34897 5321 39441
rect 7225 34897 7266 39441
rect 5280 34876 7266 34897
rect 7624 18529 9746 18550
rect 7624 13665 7653 18529
rect 9717 13665 9746 18529
rect 7624 13644 9746 13665
rect 5216 5618 7336 5660
rect 5216 4834 5244 5618
rect 7308 4834 7336 5618
rect 5216 4792 7336 4834
rect 7604 4409 9750 4450
rect 7604 3625 7645 4409
rect 9709 3625 9750 4409
rect 7604 3584 9750 3625
<< properties >>
string FIXED_BBOX 0 -406 15000 39592
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io.gds
string GDS_END 363082
string GDS_START 134
<< end >>
