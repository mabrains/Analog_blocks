**.subckt Ideal_opamp Vp Vn Out
*.ipin Vp
*.ipin Vn
*.opin Out
V1 Vp PLUS_I 0
V2 Vn MINUS_I 0
B1 Out 0 V = 'VDD/2*(1+tanh(GAIN*(V(PLUS_I)-V(MINUS_I))))' 
**.ends
** flattened .save nodes
.save I(V1)
.save I(V2)
.end
