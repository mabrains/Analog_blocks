magic
tech sky130A
magscale 1 2
timestamp 1624883982
<< pwell >>
rect 894 821 918 872
<< obsli1 >>
rect 0 1502 1716 1568
rect 0 1361 66 1502
rect 100 1397 1616 1431
rect 0 1327 797 1361
rect 0 1221 66 1327
rect 831 1291 885 1397
rect 1650 1361 1716 1502
rect 919 1327 1716 1361
rect 100 1257 1616 1291
rect 0 1187 797 1221
rect 0 1081 66 1187
rect 831 1151 885 1257
rect 1650 1221 1716 1327
rect 919 1187 1716 1221
rect 100 1117 1616 1151
rect 0 1047 797 1081
rect 0 941 66 1047
rect 831 1011 885 1117
rect 1650 1081 1716 1187
rect 919 1047 1716 1081
rect 100 977 1616 1011
rect 0 907 797 941
rect 0 801 66 907
rect 831 871 885 977
rect 1650 941 1716 1047
rect 919 907 1716 941
rect 100 837 1616 871
rect 0 767 797 801
rect 0 661 66 767
rect 831 731 885 837
rect 1650 801 1716 907
rect 919 767 1716 801
rect 100 697 1616 731
rect 0 627 797 661
rect 0 521 66 627
rect 831 591 885 697
rect 1650 661 1716 767
rect 919 627 1716 661
rect 100 557 1616 591
rect 0 487 797 521
rect 0 381 66 487
rect 831 451 885 557
rect 1650 521 1716 627
rect 919 487 1716 521
rect 100 417 1616 451
rect 0 347 797 381
rect 0 241 66 347
rect 831 311 885 417
rect 1650 381 1716 487
rect 919 347 1716 381
rect 100 277 1616 311
rect 0 207 797 241
rect 0 66 66 207
rect 831 171 885 277
rect 1650 241 1716 347
rect 919 207 1716 241
rect 100 137 1616 171
rect 1650 66 1716 207
rect 0 0 1716 66
<< obsm1 >>
rect 0 1502 1716 1568
rect 0 66 66 1502
rect 99 816 127 1474
rect 155 844 183 1502
rect 211 816 239 1474
rect 267 844 295 1502
rect 323 816 351 1474
rect 379 844 407 1502
rect 435 816 463 1474
rect 491 844 519 1502
rect 547 816 575 1474
rect 603 844 631 1502
rect 659 816 687 1474
rect 715 844 743 1502
rect 771 816 799 1474
rect 831 816 885 1474
rect 917 816 945 1474
rect 973 844 1001 1502
rect 1029 816 1057 1474
rect 1085 844 1113 1502
rect 1141 816 1169 1474
rect 1197 844 1225 1502
rect 1253 816 1281 1474
rect 1309 844 1337 1502
rect 1365 816 1393 1474
rect 1421 844 1449 1502
rect 1477 816 1505 1474
rect 1533 844 1561 1502
rect 1589 816 1617 1474
rect 99 752 1617 816
rect 99 94 127 752
rect 155 66 183 724
rect 211 94 239 752
rect 267 66 295 724
rect 323 94 351 752
rect 379 66 407 724
rect 435 94 463 752
rect 491 66 519 724
rect 547 94 575 752
rect 603 66 631 724
rect 659 94 687 752
rect 715 66 743 724
rect 771 94 799 752
rect 831 94 885 752
rect 917 94 945 752
rect 973 66 1001 724
rect 1029 94 1057 752
rect 1085 66 1113 724
rect 1141 94 1169 752
rect 1197 66 1225 724
rect 1253 94 1281 752
rect 1309 66 1337 724
rect 1365 94 1393 752
rect 1421 66 1449 724
rect 1477 94 1505 752
rect 1533 66 1561 724
rect 1589 94 1617 752
rect 1650 66 1716 1502
rect 0 0 1716 66
<< metal2 >>
rect 0 1502 803 1568
rect 0 1418 66 1502
rect 831 1474 885 1568
rect 913 1502 1716 1568
rect 94 1446 1622 1474
rect 0 1390 803 1418
rect 0 1306 66 1390
rect 831 1362 885 1446
rect 1650 1418 1716 1502
rect 913 1390 1716 1418
rect 94 1334 1622 1362
rect 0 1278 803 1306
rect 0 1194 66 1278
rect 831 1250 885 1334
rect 1650 1306 1716 1390
rect 913 1278 1716 1306
rect 94 1222 1622 1250
rect 0 1166 803 1194
rect 0 1082 66 1166
rect 831 1138 885 1222
rect 1650 1194 1716 1278
rect 913 1166 1716 1194
rect 94 1110 1622 1138
rect 0 1054 803 1082
rect 0 970 66 1054
rect 831 1026 885 1110
rect 1650 1082 1716 1166
rect 913 1054 1716 1082
rect 94 998 1622 1026
rect 0 942 803 970
rect 0 839 66 942
rect 831 914 885 998
rect 1650 970 1716 1054
rect 913 942 1716 970
rect 94 886 1622 914
rect 831 811 885 886
rect 1650 839 1716 942
rect 0 757 1716 811
rect 0 626 66 729
rect 831 682 885 757
rect 94 654 1622 682
rect 0 598 803 626
rect 0 514 66 598
rect 831 570 885 654
rect 1650 626 1716 729
rect 913 598 1716 626
rect 94 542 1622 570
rect 0 486 803 514
rect 0 402 66 486
rect 831 458 885 542
rect 1650 514 1716 598
rect 913 486 1716 514
rect 94 430 1622 458
rect 0 374 803 402
rect 0 290 66 374
rect 831 346 885 430
rect 1650 402 1716 486
rect 913 374 1716 402
rect 94 318 1622 346
rect 0 262 803 290
rect 0 178 66 262
rect 831 234 885 318
rect 1650 290 1716 374
rect 913 262 1716 290
rect 94 206 1622 234
rect 0 150 803 178
rect 0 66 66 150
rect 831 122 885 206
rect 1650 178 1716 262
rect 913 150 1716 178
rect 94 94 1622 122
rect 0 0 803 66
rect 831 0 885 94
rect 1650 66 1716 150
rect 913 0 1716 66
<< metal3 >>
rect 0 0 1716 1568
<< labels >>
rlabel metal2 s 1650 1418 1716 1502 6 C0
port 1 nsew
rlabel metal2 s 1650 1306 1716 1390 6 C0
port 1 nsew
rlabel metal2 s 1650 1194 1716 1278 6 C0
port 1 nsew
rlabel metal2 s 1650 1082 1716 1166 6 C0
port 1 nsew
rlabel metal2 s 1650 970 1716 1054 6 C0
port 1 nsew
rlabel metal2 s 1650 839 1716 942 6 C0
port 1 nsew
rlabel metal2 s 1650 626 1716 729 6 C0
port 1 nsew
rlabel metal2 s 1650 514 1716 598 6 C0
port 1 nsew
rlabel metal2 s 1650 402 1716 486 6 C0
port 1 nsew
rlabel metal2 s 1650 290 1716 374 6 C0
port 1 nsew
rlabel metal2 s 1650 178 1716 262 6 C0
port 1 nsew
rlabel metal2 s 1650 66 1716 150 6 C0
port 1 nsew
rlabel metal2 s 913 1502 1716 1568 6 C0
port 1 nsew
rlabel metal2 s 913 1390 1716 1418 6 C0
port 1 nsew
rlabel metal2 s 913 1278 1716 1306 6 C0
port 1 nsew
rlabel metal2 s 913 1166 1716 1194 6 C0
port 1 nsew
rlabel metal2 s 913 1054 1716 1082 6 C0
port 1 nsew
rlabel metal2 s 913 942 1716 970 6 C0
port 1 nsew
rlabel metal2 s 913 598 1716 626 6 C0
port 1 nsew
rlabel metal2 s 913 486 1716 514 6 C0
port 1 nsew
rlabel metal2 s 913 374 1716 402 6 C0
port 1 nsew
rlabel metal2 s 913 262 1716 290 6 C0
port 1 nsew
rlabel metal2 s 913 150 1716 178 6 C0
port 1 nsew
rlabel metal2 s 913 0 1716 66 6 C0
port 1 nsew
rlabel metal2 s 0 1502 803 1568 6 C0
port 1 nsew
rlabel metal2 s 0 1418 66 1502 6 C0
port 1 nsew
rlabel metal2 s 0 1390 803 1418 6 C0
port 1 nsew
rlabel metal2 s 0 1306 66 1390 6 C0
port 1 nsew
rlabel metal2 s 0 1278 803 1306 6 C0
port 1 nsew
rlabel metal2 s 0 1194 66 1278 6 C0
port 1 nsew
rlabel metal2 s 0 1166 803 1194 6 C0
port 1 nsew
rlabel metal2 s 0 1082 66 1166 6 C0
port 1 nsew
rlabel metal2 s 0 1054 803 1082 6 C0
port 1 nsew
rlabel metal2 s 0 970 66 1054 6 C0
port 1 nsew
rlabel metal2 s 0 942 803 970 6 C0
port 1 nsew
rlabel metal2 s 0 839 66 942 6 C0
port 1 nsew
rlabel metal2 s 0 626 66 729 6 C0
port 1 nsew
rlabel metal2 s 0 598 803 626 6 C0
port 1 nsew
rlabel metal2 s 0 514 66 598 6 C0
port 1 nsew
rlabel metal2 s 0 486 803 514 6 C0
port 1 nsew
rlabel metal2 s 0 402 66 486 6 C0
port 1 nsew
rlabel metal2 s 0 374 803 402 6 C0
port 1 nsew
rlabel metal2 s 0 290 66 374 6 C0
port 1 nsew
rlabel metal2 s 0 262 803 290 6 C0
port 1 nsew
rlabel metal2 s 0 178 66 262 6 C0
port 1 nsew
rlabel metal2 s 0 150 803 178 6 C0
port 1 nsew
rlabel metal2 s 0 66 66 150 6 C0
port 1 nsew
rlabel metal2 s 0 0 803 66 6 C0
port 1 nsew
rlabel metal2 s 831 1474 885 1568 6 C1
port 2 nsew
rlabel metal2 s 831 1362 885 1446 6 C1
port 2 nsew
rlabel metal2 s 831 1250 885 1334 6 C1
port 2 nsew
rlabel metal2 s 831 1138 885 1222 6 C1
port 2 nsew
rlabel metal2 s 831 1026 885 1110 6 C1
port 2 nsew
rlabel metal2 s 831 914 885 998 6 C1
port 2 nsew
rlabel metal2 s 831 811 885 886 6 C1
port 2 nsew
rlabel metal2 s 831 682 885 757 6 C1
port 2 nsew
rlabel metal2 s 831 570 885 654 6 C1
port 2 nsew
rlabel metal2 s 831 458 885 542 6 C1
port 2 nsew
rlabel metal2 s 831 346 885 430 6 C1
port 2 nsew
rlabel metal2 s 831 234 885 318 6 C1
port 2 nsew
rlabel metal2 s 831 122 885 206 6 C1
port 2 nsew
rlabel metal2 s 831 0 885 94 6 C1
port 2 nsew
rlabel metal2 s 94 1446 1622 1474 6 C1
port 2 nsew
rlabel metal2 s 94 1334 1622 1362 6 C1
port 2 nsew
rlabel metal2 s 94 1222 1622 1250 6 C1
port 2 nsew
rlabel metal2 s 94 1110 1622 1138 6 C1
port 2 nsew
rlabel metal2 s 94 998 1622 1026 6 C1
port 2 nsew
rlabel metal2 s 94 886 1622 914 6 C1
port 2 nsew
rlabel metal2 s 94 654 1622 682 6 C1
port 2 nsew
rlabel metal2 s 94 542 1622 570 6 C1
port 2 nsew
rlabel metal2 s 94 430 1622 458 6 C1
port 2 nsew
rlabel metal2 s 94 318 1622 346 6 C1
port 2 nsew
rlabel metal2 s 94 206 1622 234 6 C1
port 2 nsew
rlabel metal2 s 94 94 1622 122 6 C1
port 2 nsew
rlabel metal2 s 0 757 1716 811 6 C1
port 2 nsew
rlabel metal3 s 0 0 1716 1568 6 MET3
port 4 nsew
rlabel pwell s 894 821 918 872 6 SUB
port 3 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 1716 1568
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 312234
string GDS_START 277482
<< end >>
