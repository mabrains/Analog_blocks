magic
tech sky130A
magscale 1 2
timestamp 1624884095
<< checkpaint >>
rect -1288 -1260 1488 1273
use sky130_fd_pr__hvdfm1sd2__example_5595914180890  sky130_fd_pr__hvdfm1sd2__example_5595914180890_0
timestamp 1624884095
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_5595914180890  sky130_fd_pr__hvdfm1sd2__example_5595914180890_1
timestamp 1624884095
transform 1 0 200 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 228 13 228 13 0 FreeSans 300 0 0 0 D
flabel comment s -28 13 -28 13 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 16026
string GDS_START 15100
<< end >>
