magic
tech sky130A
magscale 1 2
timestamp 1624884095
<< checkpaint >>
rect -1288 -1260 1544 1527
use sky130_fd_pr__dfl1sd2__example_5595914180884  sky130_fd_pr__dfl1sd2__example_5595914180884_0
timestamp 1624884095
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808115  sky130_fd_pr__hvdfl1sd__example_55959141808115_0
timestamp 1624884095
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808115  sky130_fd_pr__hvdfl1sd__example_55959141808115_1
timestamp 1624884095
transform 1 0 256 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 284 267 284 267 0 FreeSans 300 0 0 0 S
flabel comment s 128 267 128 267 0 FreeSans 300 0 0 0 D
flabel comment s -28 267 -28 267 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 40040616
string GDS_START 40039176
<< end >>
