* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre = 0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre = 0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre = 0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre = 0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt  sky130_fd_pr__nfet_01v8_lvt d g s b
+ 
.param  l = 1 w = 1 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1 
msky130_fd_pr__nfet_01v8_lvt d g s b sky130_fd_pr__nfet_01v8_lvt__model l = {l} w = {w} nf = {nf} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd} 
.model sky130_fd_pr__nfet_01v8_lvt__model.0 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.4181113+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.47213
+ k2 = -0.0321739
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 161140.0
+ ua = -1.3019497e-9
+ ub = 2.64393e-18
+ uc = 7.0152e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.03208538
+ a0 = 1.9632567
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.5148757
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11559919+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.1534679+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0047977
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 8.4345657e-5
+ alpha1 = 0.0
+ beta0 = 17.822982
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25364
+ kt2 = -0.034423
+ at = 333080.0
+ ute = -1.0777
+ ua1 = 2.6823e-9
+ ub1 = -2.4433e-18
+ uc1 = -1.9223e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.1 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.039508629e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope2/sqrt(l*w*mult))} lvth0 = 1.134335973e-07 wvth0 = 9.747549271e-08 pvth0 = -7.808371819e-13
+ k1 = 5.494703645e-01 lk1 = -6.195427239e-07 wk1 = -5.323840001e-07 pk1 = 4.264715271e-12
+ k2 = -5.912813589e-02 lk2 = 2.159196020e-07 wk2 = 1.855435259e-07 pk2 = -1.486314969e-12
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 7.304176524e+04 lvsat = 7.057197193e-01 wvsat = 6.064374137e-01 pvsat = -4.857927546e-6
+ ua = -1.340324789e-09 lua = 3.074074899e-16 wua = 2.641606831e-16 pua = -2.116085568e-21
+ ub = 2.675649026e-18 lub = -2.540884285e-25 wub = -2.183426723e-25 pub = 1.749055811e-30
+ uc = 6.984078634e-11 luc = 2.493008176e-18 wuc = 2.142285938e-18 puc = -1.716099573e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.162412689e-02 lu0 = 3.694914159e-09 wu0 = 3.175104968e-09 pu0 = -2.543449585e-14
+ a0 = 2.000299418e+00 la0 = -2.967343957e-07 wa0 = -2.549891048e-07 pa0 = 2.042615723e-12
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 5.008643009e-01 lags = 1.122397138e-07 wags = 9.644956754e-08 pags = -7.726189057e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.120409948e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.850327846e-08 wvoff = -2.449337038e-08 pvoff = 1.962065928e-13
+ nfactor = {1.261889959e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -8.685257477e-07 wnfactor = -7.463395080e-07 pnfactor = 5.978627263e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.416657520e-01 lpclm = -1.134827673e-06 wpclm = -9.751774541e-07 ppclm = 7.811756514e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 2.870867443e-03 lpdiblc2 = 1.543508488e-08 wpdiblc2 = 1.326364093e-08 ppdiblc2 = -1.062497220e-13
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.387872744e-04 lalpha0 = -4.361100204e-10 walpha0 = -3.747570396e-10 palpha0 = 3.002028742e-15
+ alpha1 = 0.0
+ beta0 = 1.812625487e+01 lbeta0 = -2.429397649e-06 wbeta0 = -2.087624289e-06 pbeta0 = 1.672312313e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.532200231e-01 lkt1 = -3.364267089e-09 wkt1 = -2.890974103e-09 pkt1 = 2.315843715e-14
+ kt2 = -3.413547734e-02 lkt2 = -2.303229007e-09 wkt2 = -1.979205347e-09 pkt2 = 1.585462235e-14
+ at = 6.184327776e+05 lat = -2.285846960e+00 wat = -1.964268648e+00 pat = 1.573497043e-5
+ ute = -9.493378244e-01 lute = -1.028258044e-06 wute = -8.836002898e-07 pute = 7.078168482e-12
+ ua1 = 2.420622075e-09 lua1 = 2.096197186e-15 wua1 = 1.801299249e-15 pua1 = -1.442948776e-20
+ ub1 = -1.549718345e-18 lub1 = -7.158125206e-24 wub1 = -6.151103360e-24 pub1 = 4.927402857e-29
+ uc1 = -1.087192054e-11 luc1 = -6.689715711e-17 wuc1 = -5.748590812e-17 puc1 = 4.604966156e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.2 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.321459564e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.543554001e-10 wvth0 = -1.949509854e-07 pvth0 = 3.919684513e-13
+ k1 = 3.594104930e-01 lk1 = 1.427113968e-07 wk1 = 1.064768000e-06 pk1 = -2.140822541e-12
+ k2 = 6.612547593e-03 lk2 = -4.773998315e-08 wk2 = -3.710870518e-07 pk2 = 7.461076263e-13
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 4.535984092e+05 lvsat = -8.205407570e-01 wvsat = -1.212874827e+00 pvsat = 2.438606128e-6
+ ua = -1.302525680e-09 lua = 1.558103804e-16 wua = -5.283213661e-16 pua = 1.062242939e-21
+ ub = 2.594422390e-18 lub = 7.167911566e-26 wub = 4.366853446e-25 pub = -8.779995538e-31
+ uc = 6.796662443e-11 luc = 1.000952193e-17 wuc = -4.284571875e-18 puc = 8.614560212e-24
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.076770586e-02 lu0 = 7.129676352e-09 wu0 = -6.350209935e-09 pu0 = 1.276773210e-14
+ a0 = 1.900878686e+00 la0 = 1.020023895e-07 wa0 = 5.099782096e-07 pa0 = -1.025362188e-12
+ keta = 1.855080090e-01 lketa = -7.439984209e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -3.747436646e-01 lags = 3.623953020e-06 wags = -1.928991351e-07 pags = 3.878430010e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.224166343e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.310926146e-08 wvoff = 4.898674077e-08 pvoff = -9.849274098e-14
+ nfactor = {7.073644128e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.355454409e-06 wnfactor = 1.492679016e-06 pnfactor = -3.001180430e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.599213500e-01 leta0 = -3.205325663e-7
+ etab = -1.398683500e-01 letab = 2.802140045e-7
+ dsub = 8.384947203e-01 ldsub = -1.116930925e-6
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.135910341e-01 lpclm = 6.910251931e-07 wpclm = 1.950354908e-06 ppclm = -3.921383578e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 4.736927973e-03 lpdiblc2 = 7.951062517e-09 wpdiblc2 = -2.652728186e-08 ppdiblc2 = 5.333575290e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.619115086e-05 lalpha0 = 3.859764520e-10 walpha0 = 7.495140793e-10 palpha0 = -1.506973008e-15
+ alpha1 = 0.0
+ beta0 = 1.372440306e+01 lbeta0 = 1.522466922e-05 wbeta0 = 4.175248578e-06 pbeta0 = -8.394754790e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.544900068e-01 lkt1 = 1.729129739e-09 wkt1 = 5.781948205e-09 pkt1 = -1.162518506e-14
+ kt2 = -3.979131572e-02 lkt2 = 2.038007638e-08 wkt2 = 3.958410694e-09 pkt2 = -7.958780542e-15
+ at = 4.556946537e+04 lat = 1.167863972e-02 wat = 3.928537295e+00 pat = -7.898717086e-6
+ ute = -1.242439401e+00 lute = 1.472551399e-07 wute = 1.767200580e-06 pute = -3.553133485e-12
+ ua1 = 2.632835910e-09 lua1 = 1.245092379e-15 wua1 = -3.602598497e-15 pua1 = 7.243384538e-21
+ ub1 = -2.899948760e-18 lub1 = -1.742891103e-24 wub1 = 1.230220672e-23 pub1 = -2.473481683e-29
+ uc1 = -2.031787642e-11 luc1 = -2.901320647e-17 wuc1 = 1.149718162e-16 puc1 = -2.311623337e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.3 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.296412904e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.390236789e-9
+ k1 = 4.289650540e-01 lk1 = 2.864996428e-9
+ k2 = -1.322128542e-02 lk2 = -7.862078495e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.825027700e+04 lvsat = 5.477019766e-2
+ ua = -9.408298839e-10 lua = -5.714151863e-16
+ ub = 2.567681588e-18 lub = 1.254441734e-25
+ uc = 5.919376580e-11 luc = 2.764823148e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.856590003e-02 lu0 = -8.549372850e-9
+ a0 = 2.194610781e+00 la0 = -4.885753589e-7
+ keta = -1.435097460e-01 lketa = -8.247532269e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 7.402628058e-01 lags = 1.382121011e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.171097954e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.439331107e-9
+ nfactor = {9.970702915e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.729717692e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.505300000e-05 lcit = -1.015956180e-11
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 5.944506760e-04 leta0 = -1.899025292e-10
+ etab = -5.430717720e-04 letab = 8.660010478e-11
+ dsub = -6.340633544e-02 ldsub = 6.964313374e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.292005660e-01 lpclm = 1.808402000e-9
+ pdiblc1 = 0.39
+ pdiblc2 = 6.955794500e-03 lpdiblc2 = 3.489809478e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.887537269e-04 lalpha0 = -1.266157192e-10
+ alpha1 = 0.0
+ beta0 = 2.119341263e+01 lbeta0 = 2.074785711e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.505779880e-01 lkt1 = -6.136375327e-9
+ kt2 = -4.652898820e-02 lkt2 = 3.392684067e-8
+ at = 3.027262960e+04 lat = 4.243445773e-2
+ ute = -1.329885400e+00 lute = 3.230740652e-7
+ ua1 = 3.274737440e-09 lua1 = -4.551483686e-17
+ ub1 = -3.913337000e-18 lub1 = 2.946272922e-25
+ uc1 = 1.290785360e-11 luc1 = -9.581685925e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.4 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.400250589e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -5.103599606e-9
+ k1 = 4.339445200e-01 lk1 = -2.167251912e-9
+ k2 = -1.418804385e-02 lk2 = -6.885072422e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.026880832e+04 lvsat = 6.283626991e-2
+ ua = -1.198824854e-09 lua = -3.106854690e-16
+ ub = 2.616425016e-18 lub = 7.618406483e-26
+ uc = 1.089428312e-10 luc = -2.262817401e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.375954300e-02 lu0 = -3.692068436e-9
+ a0 = 1.969380632e+00 la0 = -2.609577707e-7
+ keta = -4.454529355e-01 lketa = 2.226684646e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 2.902775804e+00 lags = -8.033146257e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.149895327e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.965935843e-10
+ nfactor = {1.194371862e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.735788021e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 8.114866480e-04 leta0 = -4.092390825e-10
+ etab = -8.606660737e-04 letab = 4.075609060e-10
+ dsub = 2.435057895e-01 ldsub = 3.862659439e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -6.109362400e-02 lpclm = 2.951797104e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 1.029564680e-02 lpdiblc2 = 1.145547439e-10
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.483090005e-05 lalpha0 = 9.933890479e-11
+ alpha1 = 0.0
+ beta0 = 1.835426046e+01 lbeta0 = 3.076725761e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.502470760e-01 lkt1 = -6.470794994e-9
+ kt2 = -4.901692000e-04 lkt2 = -1.259998981e-8
+ at = 7.237126840e+04 lat = -1.104266450e-4
+ ute = -1.004685520e+00 lute = -5.572933488e-9
+ ua1 = 4.088120720e-09 lua1 = -8.675199796e-16
+ ub1 = -4.763807960e-18 lub1 = 1.154113244e-24
+ uc1 = -1.743066693e-10 luc1 = 9.338213757e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.5 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {5.053773090e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.847245853e-8
+ k1 = 2.731315200e-01 lk1 = 7.994386589e-8
+ k2 = 2.685855531e-02 lk2 = -2.784346596e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 6.935343216e+04 lvsat = 3.266766098e-2
+ ua = -1.672033646e-09 lua = -6.906505991e-17
+ ub = 2.983232042e-18 lub = -1.111076028e-25
+ uc = 7.538546830e-11 luc = -5.493784512e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.311010088e-02 lu0 = -3.360463289e-9
+ a0 = 1.296832240e+00 la0 = 8.244543826e-8
+ keta = -1.428146283e-02 lketa = 2.512310660e-9
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 2.715370800e+00 lags = -7.076256305e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.192914701e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.493162827e-9
+ nfactor = {1.795148014e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.668224990e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -5.996306819e-03 leta0 = 3.066820262e-09 weta0 = -1.525114254e-24 peta0 = -4.252453317e-31
+ etab = 2.833070331e-02 letab = -1.449755230e-08 wetab = 5.169878828e-24 petab = 5.472722530e-30
+ dsub = 1.760787113e+00 ldsub = -3.884579000e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 6.596832880e-01 lpclm = -7.284898085e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 6.953949600e-03 lpdiblc2 = 1.820825334e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.658135538e-03 lalpha0 = 1.438798253e-09 walpha0 = -4.135903063e-25 palpha0 = 3.944304526e-31
+ alpha1 = 0.0
+ beta0 = 1.719950301e+01 lbeta0 = 3.666344913e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.525689680e-01 lkt1 = -5.285236939e-9
+ kt2 = -2.883937520e-02 lkt2 = 1.875114777e-9
+ at = 8.981221360e+04 lat = -9.015773264e-3
+ ute = -3.364764000e-01 lute = -3.467605102e-7
+ ua1 = 4.368482088e-09 lua1 = -1.010672494e-15
+ ub1 = -4.381560808e-18 lub1 = 9.589378486e-25
+ uc1 = 5.561182016e-11 luc1 = -2.401424313e-17 wuc1 = -2.465190329e-32 puc1 = 5.877471754e-39
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.6 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {6.162803797e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -6.737379875e-8
+ k1 = 2.569146857e-01 lk1 = 8.416997290e-8
+ k2 = 3.072747161e-02 lk2 = -2.885170554e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.954686771e+05 lvsat = -1.979718634e-4
+ ua = -6.981024429e-10 lua = -3.228715315e-16
+ ub = 1.429150534e-18 lub = 2.938860382e-25
+ uc = 8.960922466e-11 luc = -9.200495420e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.561932686e-02 lu0 = -1.408367579e-9
+ a0 = 6.005713143e+00 la0 = -1.144688925e-6
+ keta = 3.021383089e-01 lketa = -7.994668186e-08 wketa = 1.588186776e-22 pketa = -3.155443621e-29
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -3.277775429e+00 lags = 8.541882767e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.759880884e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.726830156e-8
+ nfactor = {2.114708772e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.835449655e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.893770899e-01 leta0 = 5.085585235e-08 peta0 = 6.310887242e-30
+ etab = -6.126409553e-02 letab = 8.850852274e-9
+ dsub = 1.292577563e-01 ldsub = 3.671865043e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.011325514e+00 lpclm = -1.644869450e-7
+ pdiblc1 = -1.270942857e+00 lpdiblc1 = 4.328417086e-7
+ pdiblc2 = 1.457542571e-02 lpdiblc2 = -1.653313411e-10
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 8.906043181e-03 lalpha0 = -1.574826721e-9
+ alpha1 = 0.0
+ beta0 = 3.744754421e+01 lbeta0 = -1.610294622e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.620297143e-01 lkt1 = -2.887976646e-8
+ kt2 = -3.810094857e-02 lkt2 = 4.288680798e-9
+ at = -1.210119714e+04 lat = 1.754286158e-2
+ ute = -1.022327429e+00 lute = -1.680277321e-7
+ ua1 = 1.775331440e-09 lua1 = -3.348974353e-16
+ ub1 = -2.283428800e-18 lub1 = 4.121646473e-25
+ uc1 = -1.411542557e-10 luc1 = 2.726299624e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.7 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {1.128974073e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope2/sqrt(l*w*mult))} lvth0 = 2.857099578e-8
+ k1 = 1.097236267e+00 lk1 = -7.599532043e-8
+ k2 = -2.061792656e-01 lk2 = 1.630271857e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.276902600e+05 lvsat = -6.339405556e-3
+ ua = -3.793134041e-09 lua = 2.670414910e-16
+ ub = 5.948734600e-18 lub = -5.675466848e-25
+ uc = 2.262694353e-10 luc = -3.524793157e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.199305800e-02 lu0 = -7.172007348e-10
+ a0 = 0.0
+ keta = 2.323739224e-01 lketa = -6.664958979e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 9.505873333e-01 lags = 4.826233427e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.286910051e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 8.253477489e-9
+ nfactor = {-2.225938087e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.290348373e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 6.493980999e-02 leta0 = 2.383051218e-9
+ etab = -9.420281110e-02 letab = 1.512897146e-8
+ dsub = 6.533059590e-01 ldsub = -6.316493702e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 6.990366667e-02 lpclm = 1.494805913e-8
+ pdiblc1 = 4.294484535e+00 lpdiblc1 = -6.279287523e-7
+ pdiblc2 = 7.877401933e-02 lpdiblc2 = -1.240158328e-8
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.974575979e-03 lalpha0 = -2.536890724e-10
+ alpha1 = 0.0
+ beta0 = 3.185758335e+01 lbeta0 = -5.448480825e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.900488667e-01 lkt1 = -4.479316013e-9
+ kt2 = 3.135944000e-02 lkt2 = -8.950469264e-9
+ at = 5.954280000e+04 lat = 3.887515720e-3
+ ute = -3.099299333e+00 lute = 2.278431129e-7
+ ua1 = -3.102292360e-09 lua1 = 5.947776610e-16 wua1 = -6.902532921e-31 pua1 = 1.410593221e-37
+ ub1 = 3.150130800e-18 lub1 = -6.234718125e-25 wub1 = -1.469367939e-39 pub1 = -1.751623080e-46
+ uc1 = 6.131370000e-12 luc1 = -8.096440220e-19
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.8 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 5.05e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {3.848415475e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 2.290173319e-7
+ k1 = 6.538401246e-01 wk1 = -1.250828899e-6
+ k2 = -9.550250718e-02 wk2 = 4.359319668e-7
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -4.584559308e+04 wvsat = 1.424816378e+0
+ ua = -1.392111445e-09 wua = 6.206418982e-16
+ ub = 2.718453416e-18 wub = -5.129931110e-25
+ uc = 6.942080777e-11 wuc = 5.033271399e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.100167215e-02 wu0 = 7.459865531e-9
+ a0 = 2.050288057e+00 wa0 = -5.990934010e-7
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.819561101e-01 wags = 2.266069348e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.072392592e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = -5.754683745e-8
+ nfactor = {1.408204040e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = -1.753514428e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 5.328417395e-01 wpclm = -2.291166040e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.706333615e-04 wpdiblc2 = 3.116274227e-8
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.122554897e-04 walpha0 = -8.804865197e-10
+ alpha1 = 0.0
+ beta0 = 1.853551744e+01 wbeta0 = -4.904844606e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.526532700e-01 wkt1 = -6.792303964e-9
+ kt2 = -3.374746946e-02 wkt2 = -4.650115791e-9
+ at = 1.003512433e+06 wat = -4.615022221e+0
+ ute = -7.761148308e-01 wute = -2.076006750e-6
+ ua1 = 2.067491308e-09 wua1 = 4.232127855e-15
+ ub1 = -3.438421692e-19 wub1 = -1.445193290e-23
+ uc1 = 3.977465385e-13 wuc1 = -1.350623519e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.9 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 5.05e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {3.848415475e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 2.290173319e-7
+ k1 = 6.538401246e-01 wk1 = -1.250828899e-6
+ k2 = -9.550250718e-02 wk2 = 4.359319668e-7
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -4.584559308e+04 wvsat = 1.424816378e+0
+ ua = -1.392111445e-09 wua = 6.206418982e-16
+ ub = 2.718453416e-18 wub = -5.129931110e-25
+ uc = 6.942080777e-11 wuc = 5.033271399e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.100167215e-02 wu0 = 7.459865531e-9
+ a0 = 2.050288057e+00 wa0 = -5.990934010e-7
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.819561101e-01 wags = 2.266069348e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.072392592e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = -5.754683745e-8
+ nfactor = {1.408204040e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = -1.753514428e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 5.328417395e-01 wpclm = -2.291166040e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.706333615e-04 wpdiblc2 = 3.116274227e-8
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.122554897e-04 walpha0 = -8.804865197e-10
+ alpha1 = 0.0
+ beta0 = 1.853551744e+01 wbeta0 = -4.904844606e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.526532700e-01 wkt1 = -6.792303964e-9
+ kt2 = -3.374746946e-02 wkt2 = -4.650115791e-9
+ at = 1.003512433e+06 wat = -4.615022221e+0
+ ute = -7.761148308e-01 wute = -2.076006750e-6
+ ua1 = 2.067491308e-09 wua1 = 4.232127855e-15
+ ub1 = -3.438421692e-19 wub1 = -1.445193290e-23
+ uc1 = 3.977465385e-13 wuc1 = -1.350623519e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.10 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 5.05e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {3.186186106e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.655937107e-07 wvth0 = 5.865315285e-07 pvth0 = -1.433846437e-12
+ k1 = 1.043546798e+00 lk1 = -1.562957583e-06 wk1 = -3.644586874e-06 pk1 = 9.600405734e-12
+ k2 = -2.374048848e-01 lk2 = 5.691136756e-07 wk2 = 1.308643546e-06 pk2 = -3.500097061e-12
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -1.297178753e+05 lvsat = 3.363781751e-01 wvsat = 2.802470315e+00 pvsat = -5.525218879e-6
+ ua = -1.629846028e-09 lua = 9.534583169e-16 wua = 1.724837350e-15 pua = -4.428486280e-21
+ ub = 2.613463154e-18 lub = 4.210739420e-25 wub = 3.056153890e-25 pub = -3.283111250e-30
+ uc = 1.253293868e-10 luc = -2.242269471e-16 wuc = -3.991497512e-16 puc = 1.621016430e-21
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.396846984e-02 lu0 = 2.820736117e-08 wu0 = 4.045335105e-08 pu0 = -1.323236730e-13
+ a0 = 2.043295005e+00 la0 = 2.804633571e-08 wa0 = -4.703658793e-07 pa0 = -5.162745983e-13
+ keta = 1.054644942e-01 lketa = -4.229759003e-07 wketa = 5.509915409e-07 pketa = -2.209806674e-12
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -6.179047199e-01 lags = 4.411101845e-06 wags = 1.480936464e-06 pags = -5.030614009e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-8.697351308e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.127780151e-08 wvoff = -1.949913009e-07 pvoff = 5.512347650e-13
+ nfactor = {2.163203045e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.027999010e-06 wnfactor = -8.528804583e-06 pnfactor = 2.717297870e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.717431654e-06 lcit = 5.100453139e-11 wcit = 8.754234840e-11 pcit = -3.510973425e-16
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.599213500e-01 leta0 = -3.205325663e-7
+ etab = -1.398683500e-01 letab = 2.802140045e-7
+ dsub = 1.190469989e+00 ldsub = -2.528562939e-06 wdsub = -2.422874560e-06 pdsub = 9.717180710e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.773409426e-01 lpclm = 6.236514962e-07 wpclm = -1.429048993e-06 ppclm = -3.457606629e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -7.961117476e-03 lpdiblc2 = 3.301425991e-08 wpdiblc2 = 6.088161870e-08 ppdiblc2 = -1.191905258e-13
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.076305106e-04 lalpha0 = -3.825110588e-10 walpha0 = -1.823743400e-09 palpha0 = 3.783026046e-15
+ alpha1 = 0.0
+ beta0 = 1.581270064e+01 lbeta0 = 1.092012908e-05 wbeta0 = -1.019986106e-05 pbeta0 = 2.123619298e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.795734084e-01 lkt1 = 1.079659070e-07 wkt1 = 1.784473053e-07 pkt1 = -7.429219767e-13
+ kt2 = -1.800463123e-02 lkt2 = -6.313822702e-08 wkt2 = -1.460135000e-07 pkt2 = 5.669519887e-13
+ at = 1.978121148e+06 lat = -3.908765710e+00 wat = -9.374472093e+00 pat = 1.908824966e-5
+ ute = -5.442381326e-01 lute = -9.299646858e-07 wute = -3.038972583e-06 pute = 3.862070768e-12
+ ua1 = -7.067160516e-10 lua1 = 1.112623604e-14 wua1 = 1.938570836e-14 pua1 = -6.077494999e-20
+ ub1 = 5.364266705e-18 lub1 = -2.289294145e-23 wub1 = -4.458576006e-23 pub1 = 1.208547272e-28
+ uc1 = 2.364566198e-11 luc1 = -9.323808965e-17 wuc1 = -1.876577948e-16 puc1 = 2.109392834e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.11 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 5.05e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.697118313e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.819431880e-08 wvth0 = -2.758315786e-07 pvth0 = 3.000208261e-13
+ k1 = 1.085111631e-01 lk1 = 3.170250637e-07 wk1 = 2.205892426e-06 pk1 = -2.162567947e-12
+ k2 = 1.046061518e-01 lk2 = -1.185337146e-07 wk2 = -8.110828382e-07 pk2 = 7.618248076e-13
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 6.306448244e+03 lvsat = 6.288767019e-02 wvsat = 8.221713681e-02 pvsat = -5.587783977e-8
+ ua = -8.695680040e-10 lua = -5.751566780e-16 wua = -4.905418394e-16 pua = 2.575511907e-23
+ ub = 2.878397213e-18 lub = -1.116024753e-25 wub = -2.138857611e-24 pub = 1.631746163e-30
+ uc = -8.624971096e-11 luc = 2.011739869e-16 wuc = 1.001181989e-15 puc = -1.194490566e-21
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 4.466544444e-02 lu0 = -1.340597595e-08 wu0 = -4.198712889e-08 pu0 = 3.343115594e-14
+ a0 = 2.528528788e+00 la0 = -9.475647080e-07 wa0 = -2.298574688e-06 pa0 = 3.159522033e-12
+ keta = 1.597890140e-01 lketa = -5.322007798e-07 wketa = -2.087802509e-06 pketa = 3.095752643e-12
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 7.776907494e-01 lags = 1.605117594e-06 wags = -2.576408636e-07 pags = -1.535030434e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.424255136e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.021399080e-08 wvoff = 1.742645438e-07 pvoff = -1.911910362e-13
+ nfactor = {-4.667114723e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.259707118e-06 wnfactor = 1.007616134e-05 pnfactor = -1.023416578e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 4.048786331e-05 lcit = -3.586403466e-11 wcit = -1.750846968e-10 pcit = 1.769405946e-16
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 7.633336395e-04 leta0 = -5.294586156e-10 weta0 = -1.162531212e-09 peta0 = 2.337385255e-15
+ etab = -5.914993773e-04 letab = 1.839686480e-10 wetab = 3.333586851e-10 petab = -6.702509723e-16
+ dsub = 1.896373989e-01 ldsub = -5.162889328e-07 wdsub = -1.741864502e-06 pdsub = 8.347941888e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.257307081e+00 lpclm = -1.145608421e-06 wpclm = -7.077125410e-06 ppclm = 7.898415814e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 1.062535902e-02 lpdiblc2 = -4.355709728e-09 wpdiblc2 = -2.525999779e-08 ppdiblc2 = 5.400580828e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.625105526e-04 lalpha0 = -9.073287141e-11 walpha0 = 1.806488263e-10 palpha0 = -2.470049650e-16
+ alpha1 = 0.0
+ beta0 = 2.066982985e+01 lbeta0 = 1.154385083e-06 wbeta0 = 3.604160624e-06 pbeta0 = -6.518173012e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.146409778e-01 lkt1 = -2.258723796e-08 wkt1 = -2.473778003e-07 pkt1 = 1.132419805e-13
+ kt2 = -1.442129240e-01 lkt2 = 1.906161663e-07 wkt2 = 6.724220243e-07 pkt2 = -1.078594477e-12
+ at = -7.658617393e+02 lat = 6.998451174e-02 wat = 2.136581109e-01 pat = -1.896449293e-7
+ ute = -1.419053002e+00 lute = 8.289380911e-07 wute = 6.137985649e-07 pute = -3.482190902e-12
+ ua1 = 3.748199640e-09 lua1 = 2.169182545e-15 wua1 = -3.259148076e-15 pua1 = -1.524520163e-20
+ ub1 = -4.708151405e-18 lub1 = -2.641337598e-24 wub1 = 5.471224181e-24 pub1 = 2.021015471e-29
+ uc1 = 1.746472790e-10 luc1 = -3.968419409e-16 wuc1 = -1.113357596e-15 puc1 = 2.072151303e-21
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.12 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 5.05e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.333120577e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.408707601e-09 wvth0 = 4.620995066e-08 pvth0 = -2.543434335e-14
+ k1 = 4.514845313e-01 lk1 = -2.958382216e-08 wk1 = -1.207392986e-07 pk1 = 1.887260738e-13
+ k2 = -8.231423878e-03 lk2 = -4.500060587e-09 wk2 = -4.100328710e-08 pk2 = -1.641758671e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.816690595e+05 lvsat = -1.143337848e-01 wvsat = -1.179859339e+00 pvsat = 1.219576647e-6
+ ua = -5.836471811e-10 lua = -8.641082616e-16 wua = -4.234667791e-15 pua = 3.809568806e-21
+ ub = 2.215394090e-18 lub = 5.584284799e-25 wub = 2.760556531e-24 pub = -3.319601768e-30
+ uc = 1.393033384e-10 luc = -2.676992478e-17 wuc = -2.089911051e-16 puc = 2.851036267e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 4.021542765e-02 lu0 = -8.908788978e-09 wu0 = -4.444005034e-08 pu0 = 3.591007836e-14
+ a0 = 2.002257724e+00 la0 = -4.157151709e-07 wa0 = -2.263143920e-07 pa0 = 1.065295778e-12
+ keta = -7.076898512e-01 lketa = 3.444733613e-07 wketa = 1.805147145e-06 pketa = -8.384622771e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.237255728e-01 lags = 2.266014802e-06 wags = 1.913000913e-05 pags = -2.112818951e-11
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.108157119e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.730874841e-09 wvoff = -2.873112141e-08 pvoff = 1.395638302e-14
+ nfactor = {6.156082103e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.165914847e-06 wnfactor = 3.984006410e-06 pnfactor = -4.077434013e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 4.478836202e-04 leta0 = -2.106647808e-10 weta0 = 2.502916291e-09 peta0 = -1.366915991e-15
+ etab = -7.654270721e-04 letab = 3.597399764e-10 wetab = -6.555919528e-10 petab = 3.291825424e-16
+ dsub = -1.670482755e+00 ldsub = 1.363548495e-06 wdsub = 1.317522724e-05 pdsub = -6.727271031e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -6.198471667e-01 lpclm = 7.514436613e-07 wpclm = 3.846263824e-06 ppclm = -3.140761346e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 3.901748210e-04 lpdiblc2 = 5.987967421e-09 wpdiblc2 = 6.818580219e-08 ppdiblc2 = -4.043051717e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.196680708e-04 lalpha0 = 1.944368455e-10 walpha0 = 5.839893905e-10 palpha0 = -6.546209392e-16
+ alpha1 = 0.0
+ beta0 = 1.805258342e+01 lbeta0 = 3.799374330e-06 wbeta0 = 2.076639166e-06 pbeta0 = -4.974459826e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.173339226e-01 lkt1 = -1.986574789e-08 wkt1 = -2.265626281e-07 pkt1 = 9.220616747e-14
+ kt2 = 9.152968183e-02 lkt2 = -4.762531107e-08 wkt2 = -6.334324475e-07 pkt2 = 2.411020527e-13
+ at = 8.178866141e+03 lat = 6.094496974e-02 wat = 4.418780298e-01 pat = -4.202839793e-7
+ ute = -2.481107479e-01 lute = -3.544161511e-07 wute = -5.207995930e-06 pute = 2.401314615e-12
+ ua1 = 9.514008115e-09 lua1 = -3.657743500e-15 wua1 = -3.734990977e-14 pua1 = 1.920692214e-20
+ ub1 = -1.237295257e-17 lub1 = 5.104710462e-24 wub1 = 5.237868831e-23 pub1 = -2.719452853e-29
+ uc1 = -5.389396767e-10 luc1 = 3.243090365e-16 wuc1 = 2.510006001e-15 puc1 = -1.589619948e-21
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.13 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 5.05e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {5.331111927e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -5.236614593e-08 wvth0 = -1.909103482e-07 pvth0 = 9.563928123e-14
+ k1 = 2.555436801e-01 lk1 = 7.046357643e-08 wk1 = 1.210685338e-07 pk1 = 6.525899454e-14
+ k2 = 3.010826017e-02 lk2 = -2.407630326e-08 wk2 = -2.236983086e-08 pk2 = -2.593182947e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -3.297686431e+05 lvsat = 1.468063062e-01 wvsat = 2.747416673e+00 pvsat = -7.856904850e-7
+ ua = -1.912290361e-09 lua = -1.857030541e-16 wua = 1.653843131e-15 pua = 8.028951290e-22
+ ub = 2.990337962e-18 lub = 1.627421392e-25 wub = -4.891466205e-26 pub = -1.885085777e-30
+ uc = 1.412058887e-10 luc = -2.774136697e-17 wuc = -4.530847367e-16 puc = 1.531445710e-22
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.893639592e-02 lu0 = -3.149715377e-09 wu0 = 2.873032417e-08 pu0 = -1.450714864e-15
+ a0 = 3.047767317e-01 la0 = 4.510186236e-07 wa0 = 6.828962900e-06 pa0 = -2.537128807e-12
+ keta = -1.437341228e-01 lketa = 5.651756640e-08 wketa = 8.911068031e-07 pketa = -3.717532787e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 9.316756318e+00 lags = -2.427946696e-06 wags = -4.544162742e-05 pags = 1.184208811e-11
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.244823715e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.247321578e-09 wvoff = 3.573234884e-08 pvoff = -1.895866489e-14
+ nfactor = {3.239326621e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.737557741e-07 wnfactor = -9.941220074e-06 pnfactor = 3.032786630e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.171196991e-02 leta0 = 5.998157005e-09 weta0 = 3.934463227e-08 peta0 = -2.017829617e-14
+ etab = -4.800475600e-02 letab = 2.448014133e-08 wetab = 5.254665845e-07 petab = -2.683088007e-13
+ dsub = 1.943666626e+00 ldsub = -4.818361791e-07 wdsub = -1.258878557e-06 pdsub = 6.427833910e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.376085782e+00 lpclm = -2.676797023e-07 wpclm = -4.931464028e-06 ppclm = 1.341146496e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 1.278808272e-02 lpdiblc2 = -3.424043515e-10 wpdiblc2 = -4.016013044e-08 ppdiblc2 = 1.489091603e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -5.138920428e-03 lalpha0 = 2.757267099e-09 walpha0 = 1.707685491e-08 palpha0 = -9.075878072e-15
+ alpha1 = 0.0
+ beta0 = 1.743969906e+01 lbeta0 = 4.112313081e-06 wbeta0 = -1.653425558e-06 pbeta0 = -3.069888778e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.672173493e-01 lkt1 = -4.545527026e-08 wkt1 = -5.875306704e-07 pkt1 = 2.765164499e-13
+ kt2 = 7.667981142e-03 lkt2 = -4.805526701e-09 wkt2 = -2.513038635e-07 pkt2 = 4.598719771e-14
+ at = 1.856314811e+05 lat = -2.966233548e-02 wat = -6.595863010e-01 pat = 1.421237080e-7
+ ute = 1.996209953e+00 lute = -1.500366301e-06 wute = -1.605739642e-05 pute = 7.941018503e-12
+ ua1 = 9.687473754e-09 lua1 = -3.746315055e-15 wua1 = -3.661407698e-14 pua1 = 1.883120591e-20
+ ub1 = -8.512256103e-18 lub1 = 3.133438844e-24 wub1 = 2.843426067e-23 pub1 = -1.496850378e-29
+ uc1 = 3.309565358e-10 luc1 = -1.198599696e-16 wuc1 = -1.895376652e-15 puc1 = 6.597684348e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.14 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.05e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {6.621173163e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -8.598514176e-08 wvth0 = -3.155254289e-07 pvth0 = 1.281139713e-13
+ k1 = 9.113905785e-02 lk1 = 1.133074210e-07 wk1 = 1.141141401e-06 pk1 = -2.005719946e-13
+ k2 = 4.644887520e-02 lk2 = -2.833466754e-08 wk2 = -1.082206399e-07 pk2 = -3.559108644e-15
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.024081324e+05 lvsat = -1.793896152e-02 wvsat = -7.361337813e-01 pvsat = 1.221227634e-7
+ ua = -3.572492586e-09 lua = 2.469456457e-16 wua = 1.978629571e-14 pua = -3.922422012e-21
+ ub = 4.262535660e-18 lub = -1.687925808e-25 wub = -1.950403152e-23 pub = 3.184917676e-30
+ uc = -2.180019591e-11 luc = 1.473801867e-17 wuc = 7.669034579e-16 puc = -1.647843525e-22
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = -1.178462721e-03 lu0 = 4.698216784e-09 wu0 = 1.844666042e-07 pu0 = -4.203558945e-14
+ a0 = 7.577763427e+00 la0 = -1.444321709e-06 wa0 = -1.082144394e-05 pa0 = 2.062567215e-12
+ keta = 8.184019325e-01 lketa = -1.942150896e-07 wketa = -3.553778092e-06 pketa = 7.865837251e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -3.359754981e+00 lags = 8.755521481e-07 wags = 5.643185463e-07 pags = -1.470614132e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.899302647e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.230304255e-08 wvoff = 9.597306212e-08 pvoff = -3.465739477e-14
+ nfactor = {1.333966648e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.227810349e-07 wnfactor = 5.374355517e-06 pnfactor = -9.584523694e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.302623816e-06 lcit = 1.642463767e-12 wcit = 4.338505643e-11 pcit = -1.130614571e-17
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -7.560291898e-02 leta0 = 2.264813803e-08 weta0 = -7.831815720e-07 peta0 = 1.941720327e-13
+ etab = 1.964671272e-01 letab = -3.922923143e-08 wetab = -1.774131531e-06 petab = 3.309664682e-13
+ dsub = -5.509021671e-01 ldsub = 1.682484483e-07 wdsub = 4.681982856e-06 pdsub = -9.054050933e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 8.185564234e-01 lpclm = -1.223875514e-07 wpclm = 1.326954952e-06 ppclm = -2.897974907e-13
+ pdiblc1 = -1.270952915e+00 lpdiblc1 = 4.328443297e-07 wpdiblc1 = 6.923572081e-11 ppdiblc1 = -1.804282884e-17
+ pdiblc2 = -1.920896613e-02 lpdiblc2 = 7.996026579e-09 wpdiblc2 = 2.325599289e-07 ppdiblc2 = -5.617993145e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.423466313e-02 lalpha0 = -4.897488775e-09 walpha0 = -1.055168547e-07 palpha0 = 2.287204265e-14
+ alpha1 = 0.0
+ beta0 = 5.429419371e+01 lbeta0 = -5.491968223e-06 wbeta0 = -1.159664388e-04 pbeta0 = 2.672008248e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -3.865147651e-01 lkt1 = 1.169363632e-08 wkt1 = 1.545276520e-06 pkt1 = -2.792931040e-13
+ kt2 = -1.051028938e-01 lkt2 = 2.458256332e-08 wkt2 = 4.612179405e-07 pkt2 = -1.396959844e-13
+ at = 7.102537653e+04 lat = 2.040153817e-04 wat = -5.722142389e-01 pat = 1.193545486e-7
+ ute = -6.648105127e+00 lute = 7.523422088e-07 wute = 3.872588465e-05 pute = -6.335504544e-12
+ ua1 = -1.564436843e-08 lua1 = 2.855163019e-15 wua1 = 1.199111170e-13 pua1 = -2.195925965e-20
+ ub1 = 1.306814430e-17 lub1 = -2.490413500e-24 wub1 = -1.056748562e-22 pub1 = 1.998033207e-29
+ uc1 = -4.982853807e-10 luc1 = 9.624047388e-17 wuc1 = 2.458365668e-15 puc1 = -4.748168139e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.15 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.05e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.468756752e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 6.820892244e-08 wvth0 = 1.788186980e-06 pvth0 = -2.728536138e-13
+ k1 = 1.828459196e+00 lk1 = -2.178257973e-07 wk1 = -5.033482715e-06 pk1 = 9.763113620e-13
+ k2 = -3.804817216e-01 lk2 = 5.303830422e-08 wk2 = 1.199837101e-06 pk2 = -2.528749141e-13
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.382701899e+05 lvsat = -2.477426968e-02 wvsat = -7.611935348e-01 pvsat = 1.268991525e-7
+ ua = -7.860820927e-09 lua = 1.064301028e-15 wua = 2.800053283e-14 pua = -5.488055609e-21
+ ub = 1.628561958e-17 lub = -2.460392375e-24 wub = -7.115549826e-23 pub = 1.302968724e-29
+ uc = 5.039079882e-10 luc = -8.546196121e-17 wuc = -1.911166624e-15 puc = 3.456558051e-22
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 5.632265940e-02 lu0 = -6.261497093e-09 wu0 = -2.363129607e-07 pu0 = 3.816499562e-14
+ a0 = 0.0
+ keta = 8.080350157e-01 lketa = -1.922391553e-07 wketa = -3.962649485e-06 pketa = 8.645146125e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.151353997e+00 lags = 1.573477678e-08 wags = -1.382007447e-06 pags = 2.239083211e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-5.093335580e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 8.318131024e-08 wvoff = 2.620210109e-06 pvoff = -5.157769759e-13
+ nfactor = {-4.017490158e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.342768702e-06 wnfactor = 2.612273825e-05 pnfactor = -4.913094119e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.970612224e-05 lcit = -2.361803231e-12 wcit = -1.012317983e-10 pcit = 1.625782681e-17
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -4.024696278e-01 leta0 = 8.494893274e-08 weta0 = 3.217482977e-06 peta0 = -5.683546303e-13
+ etab = -2.198226399e-01 letab = 4.011559818e-08 wetab = 8.647229346e-07 petab = -1.719991930e-13
+ dsub = 7.163498423e-01 ldsub = -7.328978467e-08 wdsub = -4.339720272e-07 pdsub = 6.969590756e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.677148020e+00 lpclm = -2.860351097e-07 wpclm = -1.106370759e-05 ppclm = 2.071862790e-12
+ pdiblc1 = 1.110385018e+01 lpdiblc1 = -1.925793140e-06 wpdiblc1 = -4.687328981e-05 ppdiblc1 = 8.934044192e-12
+ pdiblc2 = 1.548168627e-01 lpdiblc2 = -2.517329639e-08 wpdiblc2 = -5.234523186e-07 ppdiblc2 = 8.791600293e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -7.984633136e-03 lalpha0 = 1.243509092e-09 walpha0 = 6.855570983e-08 palpha0 = -1.030618815e-14
+ alpha1 = 0.0
+ beta0 = 1.903818858e+01 lbeta0 = 1.227826354e-06 wbeta0 = 8.824422678e-05 pbeta0 = -1.220247038e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = 2.000206238e-01 lkt1 = -1.001000088e-07 wkt1 = -3.373466848e-06 pkt1 = 6.582193820e-13
+ kt2 = 4.504385310e-01 lkt2 = -8.130363225e-08 wkt2 = -2.884793785e-06 pkt2 = 4.980538504e-13
+ at = -1.158710764e+05 lat = 3.582647931e-02 wat = 1.207487730e+00 pat = -2.198566467e-7
+ ute = -4.688617754e+00 lute = 3.788639155e-07 wute = 1.094031175e-05 pute = -1.039574348e-12
+ ua1 = -8.508617133e-09 lua1 = 1.495088821e-15 wua1 = 3.721524752e-14 pua1 = -6.197426918e-21
+ ub1 = 7.554705620e-18 lub1 = -1.439552088e-24 wub1 = -3.031955146e-23 pub1 = 5.617610989e-30
+ uc1 = -3.280166061e-10 luc1 = 6.378724544e-17 wuc1 = 2.300157716e-15 puc1 = -4.446623781e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.16 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 5.0e-06 wmax = 5.05e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.431261+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.40031
+ k2 = -0.007143591
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 242950.0
+ ua = -1.26631373e-9
+ ub = 2.614475e-18
+ uc = 7.0441e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.03251371
+ a0 = 1.928858
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.527887
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11890341+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.05278474+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.068446
+ pdiblc1 = 0.39
+ pdiblc2 = 0.006587
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.3789948e-5
+ alpha1 = 0.0
+ beta0 = 17.541356
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25403
+ kt2 = -0.03469
+ at = 68095.0
+ ute = -1.1969
+ ua1 = 2.9253e-9
+ ub1 = -3.2731e-18
+ uc1 = -2.6978e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.17 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 5.0e-06 wmax = 5.05e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.431261+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.40031
+ k2 = -0.007143591
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 242950.0
+ ua = -1.26631373e-9
+ ub = 2.614475e-18
+ uc = 7.0441e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.03251371
+ a0 = 1.928858
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.527887
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11890341+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.05278474+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.068446
+ pdiblc1 = 0.39
+ pdiblc2 = 0.006587
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.3789948e-5
+ alpha1 = 0.0
+ beta0 = 17.541356
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25403
+ kt2 = -0.03469
+ at = 68095.0
+ ute = -1.1969
+ ua1 = 2.9253e-9
+ ub1 = -3.2731e-18
+ uc1 = -2.6978e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.18 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 5.0e-06 wmax = 5.05e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.375025056e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.503218228e-8
+ k1 = 3.048266060e-01 lk1 = 3.829457000e-7
+ k2 = 2.784367289e-02 lk2 = -1.403199205e-7
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 4.383139702e+05 lvsat = -7.835267389e-1
+ ua = -1.280239276e-09 lua = 5.584979595e-17
+ ub = 2.675408244e-18 lub = -2.443788668e-25
+ uc = 4.442584660e-11 luc = 1.043363742e-16
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.216794712e-02 lu0 = 1.386716615e-9
+ a0 = 1.947956689e+00 la0 = -7.659720371e-8
+ keta = 2.171448000e-01 lketa = -8.708809349e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -3.177341639e-01 lags = 3.391448240e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.264962398e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.045180336e-8
+ nfactor = {4.345022689e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.479683679e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.502650000e-05 lcit = -2.015928090e-11
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.599213500e-01 leta0 = -3.205325663e-7
+ etab = -1.398683500e-01 letab = 2.802140045e-7
+ dsub = 6.993782904e-01 ldsub = -5.589905717e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 8.768744200e-02 lpclm = -7.716972729e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 4.378959080e-03 lpdiblc2 = 8.855568914e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.202347795e-05 lalpha0 = 3.842693261e-10 palpha0 = 1.262177448e-29
+ alpha1 = 0.0
+ beta0 = 1.374529394e+01 lbeta0 = 1.522448650e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.434039790e-01 lkt1 = -4.261671982e-8
+ kt2 = -4.760006260e-02 lkt2 = 5.177709706e-8
+ at = 7.801228450e+04 lat = -3.977426122e-2
+ ute = -1.160206550e+00 lute = -1.471627506e-7
+ ua1 = 3.222567210e-09 lua1 = -1.192219872e-15
+ ub1 = -3.672807280e-18 lub1 = 1.603066017e-24
+ uc1 = -1.439063870e-11 luc1 = -5.048287123e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.19 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 5.0e-06 wmax = 5.05e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.138036135e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.261681010e-8
+ k1 = 5.556228200e-01 lk1 = -1.213051679e-07 wk1 = -5.421010862e-20
+ k2 = -5.979197904e-02 lk2 = 3.588032122e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.297101440e+04 lvsat = 5.156180805e-2
+ ua = -9.689957784e-10 lua = -5.699363808e-16
+ ub = 2.444872822e-18 lub = 2.191356523e-25
+ uc = 1.166795582e-10 luc = -4.093693832e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.615508621e-02 lu0 = -6.629825244e-9
+ a0 = 2.062631391e+00 la0 = -3.071621595e-7
+ keta = -2.633870340e-01 lketa = 9.527637056e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 7.254696020e-01 lags = 1.293982748e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.071038869e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.538461481e-9
+ nfactor = {1.575622568e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.853472052e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 5.277005460e-04 leta0 = -5.569471779e-11
+ etab = -5.239310080e-04 letab = 4.811568468e-11
+ dsub = -1.634205809e-01 ldsub = 1.175752839e-06 pdsub = -5.169878828e-26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.771532904e-01 lpclm = 4.553190493e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 5.505417840e-03 lpdiblc2 = 6.590710931e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.991262076e-04 lalpha0 = -1.407982317e-10
+ alpha1 = 0.0
+ beta0 = 2.140035606e+01 lbeta0 = -1.667813984e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.647819080e-01 lkt1 = 3.657442248e-10
+ kt2 = -7.919910800e-03 lkt2 = -2.800381615e-8
+ at = 4.254043500e+04 lat = 3.154543939e-2
+ ute = -1.294642360e+00 lute = 1.231338890e-7
+ ua1 = 3.087603920e-09 lua1 = -9.208626816e-16
+ ub1 = -3.599190660e-18 lub1 = 1.455052441e-24 wub1 = 3.761581923e-37
+ uc1 = -5.101882940e-11 luc1 = 2.316176899e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.20 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 5.0e-06 wmax = 5.05e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.426783384e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -6.563986827e-9
+ k1 = 4.270119200e-01 lk1 = 8.669007648e-9
+ k2 = -1.654236752e-02 lk2 = -7.827736185e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -5.747626680e+04 lvsat = 1.328618304e-01 pvsat = -6.776263578e-21
+ ua = -1.441970692e-09 lua = -9.194793282e-17
+ ub = 2.774930444e-18 lub = -1.144205807e-25
+ uc = 9.694299559e-11 luc = -2.099116814e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.120788752e-02 lu0 = -1.630186248e-9
+ a0 = 1.956386129e+00 la0 = -1.997906976e-7
+ keta = -3.418051320e-01 lketa = 1.745257004e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.001181235e+00 lags = -2.016451428e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.166392140e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.097940139e-9
+ nfactor = {1.423125243e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.394610015e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 9.551990035e-04 leta0 = -4.877245624e-10
+ etab = -8.983088033e-04 letab = 4.264618846e-10
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.597508640e-01 lpclm = 1.148437108e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 1.421073408e-02 lpdiblc2 = -2.206881661e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.299440988e-06 lalpha0 = 6.175192876e-11
+ alpha1 = 0.0
+ beta0 = 1.847349677e+01 lbeta0 = 2.791102599e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.632558320e-01 lkt1 = -1.176508181e-9
+ kt2 = -3.686054600e-02 lkt2 = 1.243589788e-9
+ at = 9.774298800e+04 lat = -2.424226067e-2
+ ute = -1.303717840e+00 lute = 1.323055691e-7
+ ua1 = 1.943566400e-09 lua1 = 2.353016362e-16
+ ub1 = -1.756332360e-18 lub1 = -4.073401570e-25
+ uc1 = -3.018733280e-11 luc1 = 2.109458528e-18 wuc1 = 3.155443621e-30
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.21 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 5.0e-06 wmax = 5.05e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.600650913e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.378524963e-07 wvth0 = 2.616917201e-06 pvth0 = -1.336197923e-12
+ k1 = 2.800830240e-01 lk1 = 8.369090195e-8
+ k2 = 6.497932819e-02 lk2 = -4.945271402e-08 wk2 = -1.944114756e-07 pk2 = 9.926649944e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -2.356249646e+04 lvsat = 1.155454593e-01 wvsat = 1.236702718e+00 pvsat = -6.314604078e-7
+ ua = -1.134656613e-08 lua = 4.965338495e-15 wua = 4.819925776e-14 pua = -2.461054101e-20
+ ub = 1.144221286e-17 lub = -4.539934984e-24 wub = -4.174750727e-23 pub = 2.131627721e-29
+ uc = 4.937028284e-11 luc = 3.299458988e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = -6.081337997e-02 lu0 = 4.535587293e-08 wu0 = 4.715243060e-07 pu0 = -2.407603106e-13
+ a0 = 1.688937120e+00 la0 = -6.323123347e-8
+ keta = 3.688404081e-02 lketa = -1.883299124e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.062068424e-01 lags = -2.767750313e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.172397928e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.404595627e-9
+ nfactor = {-1.175698395e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.069224757e-06 wnfactor = 6.404532759e-05 pnfactor = -3.270154427e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -3.737219299e-03 leta0 = 1.908224365e-9
+ etab = 5.850190428e-02 letab = -2.990328692e-08 wetab = 1.111730743e-21 petab = -3.534096855e-28
+ dsub = 1.688504919e+00 ldsub = -3.515506114e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.765288560e-01 lpclm = 4.156868126e-9
+ pdiblc1 = 0.39
+ pdiblc2 = 4.648038240e-03 lpdiblc2 = 2.675830835e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.677617963e-03 lalpha0 = 9.176801660e-10 walpha0 = -2.646977960e-23 palpha0 = -2.524354897e-29
+ alpha1 = 0.0
+ beta0 = 1.710456674e+01 lbeta0 = 3.490078270e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.863037600e-01 lkt1 = 1.059176386e-8
+ kt2 = -4.326872160e-02 lkt2 = 4.515604249e-9
+ at = 5.194013680e+04 lat = -8.553248501e-4
+ ute = -1.258458784e+00 lute = 1.091962951e-7
+ ua1 = 2.266177760e-09 lua1 = 7.057627574e-17
+ ub1 = -2.748924560e-18 lub1 = 9.947742034e-26
+ uc1 = -5.321677440e-11 luc1 = 1.386829141e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.22 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.0e-06 wmax = 5.05e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {2.492528357e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -4.210836899e-07 wvth0 = -9.346132862e-06 pvth0 = 1.781372923e-12
+ k1 = 3.224366571e-01 lk1 = 7.265354515e-8
+ k2 = -1.162191978e-01 lk2 = -2.232378139e-09 wk2 = 6.943266986e-07 pk2 = -1.323386687e-13
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.048440307e+06 lvsat = -1.638184714e-01 wvsat = -4.416795421e+00 pvsat = 8.418412073e-7
+ ua = 3.532903103e-08 lua = -7.198322123e-15 wua = -1.721402063e-13 pua = 3.280992332e-20
+ ub = -2.991140691e-17 lub = 6.236818329e-24 wub = 1.490982402e-22 pub = -2.841812459e-29
+ uc = 1.336432299e-10 luc = -1.866207102e-17 wuc = 1.262177448e-29
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.775435753e-01 lu0 = -6.887994960e-08 wu0 = -1.684015379e-06 pu0 = 3.209733311e-13
+ a0 = 5.384368286e+00 la0 = -1.026260595e-6
+ keta = 9.808774473e-02 lketa = -3.478267648e-08 pketa = 1.615587134e-27
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -3.245373429e+00 lags = 8.457443155e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.704775143e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.527834587e-8
+ nfactor = {4.878517789e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -8.708062620e-06 wnfactor = -2.287333128e-04 pnfactor = 4.359656943e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 7.491079919e-06 lcit = -6.491754269e-13
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -2.343457508e-01 leta0 = 6.200480756e-08 peta0 = 1.615587134e-27
+ etab = -1.631310468e-01 letab = 2.785426014e-08 wetab = -1.355252716e-20
+ dsub = 3.980874970e-01 ldsub = -1.526783136e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.087516514e+00 lpclm = -1.811265156e-7
+ pdiblc1 = -1.270938882e+00 lpdiblc1 = 4.328406726e-7
+ pdiblc2 = 2.792853429e-02 lpdiblc2 = -3.391066435e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.847484325e-03 lalpha0 = -2.615614903e-10
+ alpha1 = 0.0
+ beta0 = 3.078899191e+01 lbeta0 = -7.608292872e-8
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -7.330314286e-02 lkt1 = -4.491619697e-8
+ kt2 = -1.161877143e-02 lkt2 = -3.732372766e-9
+ at = -4.495655143e+04 lat = 2.439595210e-2
+ ute = 1.201232514e+00 lute = -5.317992572e-7
+ ua1 = 8.660378971e-09 lua1 = -1.595752560e-15
+ ub1 = -8.351059771e-18 lub1 = 1.559393856e-24
+ uc1 = 0.0
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.23 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.0e-06 wmax = 5.05e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-7.386775378e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.947841537e-07 wvth0 = 4.707930239e-06 pvth0 = -8.973315036e-13
+ k1 = 8.082241333e-01 lk1 = -1.993754781e-8
+ k2 = -4.102284470e-01 lk2 = 5.380578475e-08 wk2 = 1.346597033e-06 pk2 = -2.566613945e-13
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 4.385330472e+04 lvsat = 2.765581132e-02 wvsat = 6.913563310e-01 pvsat = -1.317725167e-7
+ ua = -1.301021841e-08 lua = 2.015138821e-15 wua = 5.340585774e-14 pua = -1.017915649e-20
+ ub = -1.420528542e-18 lub = 8.064569121e-25 wub = 1.620043940e-23 pub = -3.087803749e-30
+ uc = 1.165342133e-10 luc = -1.540109246e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = -9.635991765e-02 lu0 = 2.144605615e-08 wu0 = 5.169694356e-07 pu0 = -9.853437442e-14
+ a0 = 0.0
+ keta = 4.846811240e-03 lketa = -1.701095456e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 8.712353333e-01 lags = 6.111868547e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {2.175602256e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.136136626e-8
+ nfactor = {-8.269658632e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.635236164e-05 wnfactor = 4.142978611e-04 pnfactor = -7.896517232e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -8.125198107e-07 lcit = 9.334906816e-13
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 2.496810064e-01 leta0 = -3.025069235e-8
+ etab = -4.455221445e-02 letab = 5.253134690e-9
+ dsub = 6.283881857e-01 ldsub = -5.916314262e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -5.653514667e-01 lpclm = 1.339101215e-7
+ pdiblc1 = 1.603117493e+00 lpdiblc1 = -1.149544725e-7
+ pdiblc2 = 4.871847333e-02 lpdiblc2 = -7.353628817e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.910902588e-03 lalpha0 = -8.454490111e-10
+ alpha1 = 0.0
+ beta0 = 3.692438375e+01 lbeta0 = -1.245488613e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -4.837463333e-01 lkt1 = 3.331427513e-8
+ kt2 = -1.342794333e-01 lkt2 = 1.964674939e-08 wkt2 = -1.355252716e-20
+ at = 1.288742400e+05 lat = -8.736196744e-3
+ ute = -2.471129333e+00 lute = 1.681529109e-7
+ ua1 = -9.654700667e-10 lua1 = 2.389342667e-16
+ ub1 = 1.409245067e-18 lub1 = -3.009202457e-25 pub1 = 1.121038771e-44
+ uc1 = 1.382016533e-10 luc1 = -2.634123513e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.24 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 3.01e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.396315006e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = -4.087859533e-8
+ k1 = 2.494330533e-01 wk1 = 7.368302009e-7
+ k2 = 5.272278487e-02 wk2 = -2.923664265e-7
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.493316251e+05 wvsat = -5.195306235e-1
+ ua = -1.506061110e-09 wua = 1.170842292e-15
+ ub = 2.915846466e-18 wub = -1.471792762e-24
+ uc = 7.252139330e-11 wuc = -1.015991275e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.257610524e-02 wu0 = -3.047164989e-10
+ a0 = 2.284318619e+00 wa0 = -1.735945252e-6
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 5.124209497e-01 wags = 7.553077663e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.248638928e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = 2.910891169e-8
+ nfactor = {5.307523946e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 2.549423263e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.727047739e-05 wcit = -3.550646689e-11
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.228460764e-01 wpclm = 9.342035491e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 6.405965113e-03 wpdiblc2 = 8.841110256e-10
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.647008226e-05 walpha0 = 3.574766232e-11
+ alpha1 = 0.0
+ beta0 = 1.717144284e+01 wbeta0 = 1.806526428e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.514562510e-01 wkt1 = -1.256928928e-8
+ kt2 = -3.455913141e-02 wkt2 = -6.391164040e-10
+ at = -2.959886961e+05 wat = 1.778057342e+0
+ ute = -1.103692480e+00 wute = -4.551929055e-7
+ ua1 = 4.147321839e-09 wua1 = -5.967926955e-15
+ ub1 = -4.995330683e-18 wub1 = 8.410771877e-24
+ uc1 = 1.877070653e-12 wuc1 = -1.409180658e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.25 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 3.01e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.396315006e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = -4.087859533e-8
+ k1 = 2.494330533e-01 wk1 = 7.368302009e-7
+ k2 = 5.272278487e-02 wk2 = -2.923664265e-7
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.493316251e+05 wvsat = -5.195306235e-1
+ ua = -1.506061110e-09 wua = 1.170842292e-15
+ ub = 2.915846466e-18 wub = -1.471792762e-24
+ uc = 7.252139330e-11 wuc = -1.015991275e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.257610524e-02 wu0 = -3.047164989e-10
+ a0 = 2.284318619e+00 wa0 = -1.735945252e-6
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 5.124209497e-01 wags = 7.553077663e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.248638928e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = 2.910891169e-8
+ nfactor = {5.307523946e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 2.549423263e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.727047739e-05 wcit = -3.550646689e-11
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.228460764e-01 wpclm = 9.342035491e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 6.405965113e-03 wpdiblc2 = 8.841110256e-10
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.647008226e-05 walpha0 = 3.574766232e-11
+ alpha1 = 0.0
+ beta0 = 1.717144284e+01 wbeta0 = 1.806526428e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.514562510e-01 wkt1 = -1.256928928e-8
+ kt2 = -3.455913141e-02 wkt2 = -6.391164040e-10
+ at = -2.959886961e+05 wat = 1.778057342e+0
+ ute = -1.103692480e+00 wute = -4.551929055e-7
+ ua1 = 4.147321839e-09 wua1 = -5.967926955e-15
+ ub1 = -4.995330683e-18 wub1 = 8.410771877e-24
+ uc1 = 1.877070653e-12 wuc1 = -1.409180658e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.26 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 3.01e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.688440581e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.171598829e-07 wvth0 = -1.530611728e-07 pvth0 = 4.499194452e-13
+ k1 = -7.492470859e-02 lk1 = 1.300869240e-06 wk1 = 1.854572508e-06 pk1 = -4.482817295e-12
+ k2 = 1.820446314e-01 lk2 = -5.186581976e-07 wk2 = -7.530635110e-07 pk2 = 1.847671727e-12
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 6.362877347e+05 lvsat = -1.150866173e+00 wvsat = -9.668345752e-01 pvsat = 1.793957228e-6
+ ua = -1.736282479e-09 lua = 9.233258244e-16 wua = 2.227155389e-15 pua = -4.236449307e-21
+ ub = 3.277098198e-18 lub = -1.448836194e-24 wub = -2.938443144e-24 pub = 5.882148025e-30
+ uc = 3.777155232e-11 luc = 1.393677122e-16 wuc = 3.249724426e-17 puc = -1.710807939e-22
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.149368176e-02 lu0 = 4.341167586e-09 wu0 = 3.292876003e-09 pu0 = -1.442850449e-14
+ a0 = 2.531747594e+00 la0 = -9.923386451e-07 wa0 = -2.851030449e-06 pa0 = 4.472160690e-12
+ keta = 1.647976638e-01 lketa = -6.609375105e-07 wketa = 2.556450916e-07 pketa = -1.025290205e-12
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.976295675e-01 lags = 1.262502317e-06 wags = -2.516856087e-06 pags = 1.039702675e-11
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.480268893e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 9.289751387e-08 wvoff = 1.051481562e-07 pvoff = -3.049629941e-13
+ nfactor = {-1.113825429e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.595743820e-06 wnfactor = 7.561490562e-06 pnfactor = -2.010139711e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.960598830e-05 lcit = -4.947280008e-11 wcit = -7.120111806e-11 pcit = 1.431569680e-16
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.599213500e-01 leta0 = -3.205325663e-7
+ etab = -1.398569041e-01 letab = 2.801680995e-07 wetab = -5.589782372e-11 petab = 2.241838118e-16
+ dsub = 5.866338881e-01 ldsub = -1.068178715e-07 wdsub = 5.506042007e-07 pdsub = -2.208253207e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -9.936540810e-02 lpclm = -9.417156841e-08 wpclm = 9.135006514e-07 ppclm = 8.303104142e-14
+ pdiblc1 = 0.39
+ pdiblc2 = 2.846049534e-03 lpdiblc2 = 1.427739742e-08 wpdiblc2 = 7.486193705e-09 ppdiblc2 = -2.647831279e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -5.782516840e-05 lalpha0 = 3.380745323e-10 walpha0 = -2.050307442e-11 palpha0 = 2.255992048e-16
+ alpha1 = 0.0
+ beta0 = 1.322558698e+01 lbeta0 = 1.582524948e-05 wbeta0 = 2.538066886e-06 pbeta0 = -2.933916164e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.219583638e-01 lkt1 = -1.183042264e-07 wkt1 = -1.047328786e-07 pkt1 = 3.696312913e-13
+ kt2 = -6.838465965e-02 lkt2 = 1.356606636e-07 wkt2 = 1.015046974e-07 pkt2 = -4.096579795e-13
+ at = -6.747470705e+05 lat = 1.519048337e+00 wat = 3.676213224e+00 pat = -7.612743980e-6
+ ute = -9.395298795e-01 lute = -6.583905251e-07 wute = -1.077707622e-06 pute = 2.496657521e-12
+ ua1 = 5.086904929e-09 lua1 = -3.768291938e-15 wua1 = -9.104772899e-15 pua1 = 1.258063434e-20
+ ub1 = -6.577051209e-18 lub1 = 6.343648340e-24 wub1 = 1.418331086e-23 pub1 = -2.315134486e-29
+ uc1 = 2.302620734e-11 luc1 = -8.482072760e-17 wuc1 = -1.827307802e-16 puc1 = 1.676940723e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.27 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 3.01e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {3.863920332e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.861815826e-08 wvth0 = 1.338685642e-07 pvth0 = -1.269814840e-13
+ k1 = 7.131484205e-01 lk1 = -2.836305937e-07 wk1 = -7.692998991e-07 pk1 = 7.927405659e-13
+ k2 = -1.265747776e-01 lk2 = 1.018519861e-07 wk2 = 3.261438144e-07 pk2 = -3.221825214e-13
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 5.978344050e+04 lvsat = 8.253360795e-03 wvsat = -1.797790047e-01 pvsat = 2.115032984e-7
+ ua = -9.537569882e-10 lua = -6.500199281e-16 wua = -7.442091797e-17 pua = 3.911000156e-22
+ ub = 2.214939918e-18 lub = 6.867392441e-25 wub = 1.122911827e-24 pub = -2.283612281e-30
+ uc = 1.344390431e-10 luc = -5.499194470e-17 wuc = -8.673110840e-17 puc = 6.863973193e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.512322968e-02 lu0 = -2.956401448e-09 wu0 = 5.039226164e-09 pu0 = -1.793971612e-14
+ a0 = 1.995617801e+00 la0 = 8.560391543e-08 wa0 = 3.272709196e-07 pa0 = -1.918132042e-12
+ keta = -1.827045369e-01 lketa = 3.775041422e-08 wketa = -3.940250771e-07 pketa = 2.809366367e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.976885917e-01 lags = 2.258389008e-06 wags = 4.996746513e-06 pags = -4.709822632e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-8.875202117e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.628053598e-08 wvoff = -8.962408901e-08 pvoff = 8.664608212e-14
+ nfactor = {2.807009285e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.287486457e-06 wnfactor = -6.013661742e-06 pnfactor = 7.192804115e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 5.177372757e-04 leta0 = -3.566256658e-11 weta0 = 4.865712486e-11 peta0 = -9.783001524e-17
+ etab = -5.415766835e-04 letab = 6.070225757e-11 wetab = 8.617530295e-11 petab = -6.146841665e-17
+ dsub = -2.534808307e-01 ldsub = 1.582316782e-06 wdsub = 4.398227389e-07 pdsub = -1.985516000e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -8.396780468e-01 lpclm = 1.394301023e-06 wpclm = 3.235539027e-06 ppclm = -4.585659316e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 9.610058591e-03 lpdiblc2 = 6.776808117e-10 wpdiblc2 = -2.004562880e-08 ppdiblc2 = 2.887716954e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.429512492e-04 lalpha0 = -6.560653286e-11 walpha0 = 2.743388360e-10 palpha0 = -3.672099403e-16
+ alpha1 = 0.0
+ beta0 = 2.033465129e+01 lbeta0 = 1.531764794e-06 wbeta0 = 5.204529110e-06 pbeta0 = -8.295105110e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.984823825e-01 lkt1 = 3.555496559e-08 wkt1 = 1.645813222e-07 pkt1 = -1.718518409e-13
+ kt2 = 5.574947439e-02 lkt2 = -1.139234263e-07 wkt2 = -3.109389930e-07 pkt2 = 4.196013043e-13
+ at = 9.282907453e+04 lat = -2.424026075e-02 wat = -2.455921144e-01 pat = 2.724378345e-7
+ ute = -1.264455280e+00 lute = -5.095515458e-09 wute = -1.474231346e-07 pute = 6.262275312e-13
+ ua1 = 5.028816322e-09 lua1 = -3.651498986e-15 wua1 = -9.480201947e-15 pua1 = 1.333547199e-20
+ ub1 = -6.020880034e-18 lub1 = 5.225410576e-24 wub1 = 1.182668331e-23 pub1 = -1.841310950e-29
+ uc1 = -9.789132403e-11 luc1 = 1.582960610e-16 wuc1 = 2.289088584e-16 puc1 = -6.599485851e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.28 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 3.01e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.462953823e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.192016635e-08 wvth0 = -1.766437675e-08 pvth0 = 2.615770613e-14
+ k1 = 4.013290284e-01 lk1 = 3.149408394e-08 wk1 = 1.254262534e-07 pk1 = -1.114696838e-13
+ k2 = -1.454307333e-02 lk2 = -1.136725423e-08 wk2 = -9.763853059e-09 pk2 = 1.728576730e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -9.163355237e+04 lvsat = 1.612753738e-01 wvsat = 1.668122277e-01 pvsat = -1.387618010e-7
+ ua = -1.034320785e-09 lua = -5.686021551e-16 wua = -1.990819471e-15 pua = 2.327812393e-21
+ ub = 2.583603010e-18 lub = 3.141683229e-25 wub = 9.343762224e-25 pub = -2.093078199e-30
+ uc = 9.363132046e-11 luc = -1.375166021e-17 wuc = 1.617306223e-17 puc = -3.535522291e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.813730840e-02 lu0 = -6.002429405e-09 wu0 = -3.384086627e-08 pu0 = 2.135250529e-14
+ a0 = 2.964782162e+00 la0 = -8.938335876e-07 wa0 = -4.924653286e-06 pa0 = 3.389462560e-12
+ keta = -3.117534833e-01 lketa = 1.681672794e-07 wketa = -1.467617344e-07 pketa = 3.105230257e-14
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.984823776e+00 lags = -3.080117991e-06 wags = -4.803765898e-06 pags = 5.194575210e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.100549538e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.751792266e-09 wvoff = -3.215522253e-08 pvoff = 2.856804566e-14
+ nfactor = {1.562156034e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.943776145e-08 wnfactor = -6.789777215e-07 pnfactor = 1.801572444e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 9.899747706e-04 leta0 = -5.129056788e-10 weta0 = -1.698326577e-10 peta0 = 1.229757590e-16
+ etab = -9.627047148e-04 letab = 4.862942460e-10 wetab = 3.144870931e-10 petab = -2.922003118e-16
+ dsub = 1.631098109e+00 ldsub = -3.222386945e-07 wdsub = -3.082062281e-06 pdsub = 1.573701000e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 5.642046070e-01 lpclm = -2.446278698e-08 wpclm = -1.975210522e-06 ppclm = 6.803241781e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 1.220658290e-02 lpdiblc2 = -1.946366655e-09 wpdiblc2 = 9.787572910e-09 ppdiblc2 = -1.272264110e-15
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.070122836e-05 lalpha0 = 5.793933817e-11 walpha0 = -1.074435689e-10 palpha0 = 1.861935806e-17
+ alpha1 = 0.0
+ beta0 = 1.942818654e+01 lbeta0 = 2.447838063e-06 wbeta0 = -4.662370716e-06 pbeta0 = 1.676383854e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.503310462e-01 lkt1 = -1.310677488e-08 wkt1 = -6.312013024e-08 pkt1 = 5.826324697e-14
+ kt2 = -6.589998840e-02 lkt2 = 9.015520761e-09 wkt2 = 1.418184729e-07 pkt2 = -3.795539070e-14
+ at = 1.198833680e+05 lat = -5.158132970e-02 wat = -1.081258666e-01 pat = 1.335144444e-7
+ ute = -2.238208352e+00 lute = 9.789793391e-07 wute = 4.563724588e-06 pute = -4.134858357e-12
+ ua1 = -2.726467352e-09 lua1 = 4.185990695e-15 wua1 = 2.280681033e-14 pua1 = -1.929378262e-20
+ ub1 = 4.584300525e-18 lub1 = -5.492184897e-24 wub1 = -3.096543179e-23 pub1 = 2.483260202e-29
+ uc1 = 1.840337005e-10 luc1 = -1.266173688e-16 wuc1 = -1.046180549e-15 puc1 = 6.286567704e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.29 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 3.01e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.986357867e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.864517681e-08 wvth0 = 5.911353450e-09 pvth0 = 1.411993829e-14
+ k1 = 3.022304018e-01 lk1 = 8.209384270e-08 wk1 = -1.081600416e-07 pk1 = 7.799478407e-15
+ k2 = 2.269182158e-02 lk2 = -3.037939157e-08 wk2 = 1.210590608e-08 pk2 = 6.119068285e-15
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.831693614e+05 lvsat = -3.009899396e-02 wvsat = -2.612683195e-01 pvsat = 7.981612636e-8
+ ua = -3.334837986e-09 lua = 6.060419277e-16 wua = 9.072781630e-15 pua = -3.321262329e-21
+ ub = 4.771594755e-18 lub = -8.030202619e-25 wub = -9.170543144e-24 pub = 3.066493629e-30
+ uc = 4.954613784e-11 luc = 8.758234036e-18 wuc = -8.588142757e-19 puc = -2.665874676e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.453324036e-02 lu0 = 9.438077358e-10 wu0 = 5.472128360e-08 pu0 = -2.386732843e-14
+ a0 = 1.045429869e+00 la0 = 8.618769327e-08 wa0 = 3.142664187e-06 pa0 = -7.297097416e-13
+ keta = 7.608545142e-02 lketa = -2.986328062e-08 wketa = -1.914459690e-07 pketa = 5.386807273e-14
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.139467883e+00 lags = 5.575453303e-07 wags = 1.096708937e-05 pags = -2.858023490e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.254556026e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.111779014e-09 wvoff = 4.012313980e-08 pvoff = -8.337286147e-15
+ nfactor = {-2.786158941e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 9.104603851e-07 wnfactor = 7.988995421e-06 pnfactor = -2.624294643e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 3.238031453e-03 leta0 = -1.660763306e-09 weta0 = -3.406468358e-08 peta0 = 1.742968664e-14
+ etab = 1.156574142e-01 letab = -5.905993846e-08 wetab = -2.791275059e-07 petab = 1.423908813e-13
+ dsub = 1.574327190e+00 ldsub = -2.932514631e-07 wdsub = 5.576040647e-07 pdsub = -2.847126354e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 5.996401639e-01 lpclm = -4.255618234e-08 wpclm = -1.089597539e-06 ppclm = 2.281301889e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 4.902668738e-03 lpdiblc2 = 1.783011916e-09 wpdiblc2 = -1.243526231e-09 ppdiblc2 = 4.360215111e-15
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.396392408e-03 lalpha0 = 7.815073487e-10 walpha0 = -1.373407182e-09 palpha0 = 6.650203792e-16
+ alpha1 = 0.0
+ beta0 = 1.764033415e+01 lbeta0 = 3.360715495e-06 wbeta0 = -2.616500484e-06 pbeta0 = 6.317625134e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -3.460514846e-01 lkt1 = 3.576808097e-08 wkt1 = 2.917869752e-07 pkt1 = -1.229523211e-13
+ kt2 = -6.032463105e-02 lkt2 = 6.168743301e-09 wkt2 = 8.329509220e-08 pkt2 = -8.073352529e-15
+ at = -4.768550074e+02 lat = 9.874600155e-03 wat = 2.559862420e-01 pat = -5.240119825e-8
+ ute = -1.072179475e+00 lute = 3.836049946e-07 wute = -9.097229479e-07 pute = -1.340116045e-12
+ ua1 = 4.705219949e-09 lua1 = 3.913711593e-16 wua1 = -1.191142839e-14 pua1 = -1.566649933e-21
+ ub1 = -6.455251943e-18 lub1 = 1.446105931e-25 wub1 = 1.810040573e-23 pub1 = -2.204146190e-31
+ uc1 = -1.763003973e-10 luc1 = 5.736922150e-17 wuc1 = 6.010973348e-16 puc1 = -2.124433172e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.30 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.01e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {6.226325442e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -7.095873181e-08 wvth0 = -2.142161733e-07 pvth0 = 7.148517175e-14
+ k1 = 3.376497671e-01 lk1 = 7.286355611e-08 wk1 = -7.429550421e-08 pk1 = -1.025620028e-15
+ k2 = 1.583106600e-02 lk2 = -2.859147867e-08 wk2 = 4.943942772e-08 pk2 = -3.610047456e-15
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 9.902217631e+04 lvsat = 1.788976246e-02 wvsat = 2.198304345e-01 pvsat = -4.555820893e-8
+ ua = 3.581993886e-09 lua = -1.196484458e-15 wua = -1.709878833e-14 pua = 3.499048803e-21
+ ub = -2.255406308e-18 lub = 1.028216215e-24 wub = 1.403601290e-23 pub = -2.981134876e-30
+ uc = 2.251955405e-10 luc = -3.701600029e-17 wuc = -4.471094413e-16 puc = 8.963416665e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 6.493074078e-02 lu0 = -9.583780873e-09 wu0 = -1.573237093e-07 pu0 = 3.139159673e-14
+ a0 = 5.123238816e+00 la0 = -9.764893183e-07 wa0 = 1.275264936e-06 pa0 = -2.430654968e-13
+ keta = -1.877737008e-02 lketa = -5.142029332e-09 wketa = 5.707283180e-07 pketa = -1.447545464e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -3.444921859e+00 lags = 8.977466365e-07 wags = 9.745246929e-07 pags = -2.539611350e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.849812979e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.862417520e-08 wvoff = 7.083140257e-08 pvoff = -1.633985942e-14
+ nfactor = {3.978877490e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.990423907e-07 wnfactor = -9.915023876e-06 pnfactor = 2.041492786e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.111334796e-05 lcit = -1.593138479e-12 wcit = -1.768988933e-11 pcit = 4.609985160e-18
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -3.020870465e-01 leta0 = 7.790695193e-08 weta0 = 3.308247791e-07 peta0 = -7.766050733e-14
+ etab = -3.582479906e-01 letab = 6.443981004e-08 wetab = 9.528828627e-07 petab = -1.786710207e-13
+ dsub = 8.749634155e-01 ldsub = -1.109972635e-07 wdsub = -2.328895079e-06 pdsub = 4.675090415e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.544024081e+00 lpclm = -2.886626311e-07 wpclm = -2.229423178e-06 ppclm = 5.251687504e-13
+ pdiblc1 = -1.282696956e+00 lpdiblc1 = 4.359048268e-07 wpdiblc1 = 5.742232066e-08 ppdiblc1 = -1.496425676e-14
+ pdiblc2 = 2.474131487e-02 lpdiblc2 = -3.386939267e-09 wpdiblc2 = 1.556526409e-08 ppdiblc2 = -2.015564563e-17
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.734655581e-03 lalpha0 = 8.696587316e-10 walpha0 = 2.237756755e-08 palpha0 = -5.524483637e-15
+ alpha1 = 0.0
+ beta0 = 2.404367742e+01 lbeta0 = 1.692004240e-06 wbeta0 = 3.294175513e-05 pbeta0 = -8.634718900e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = 8.962210664e-02 lkt1 = -7.776845691e-08 wkt1 = -7.956698947e-07 pkt1 = 1.604389392e-13
+ kt2 = -1.442438218e-02 lkt2 = -5.792861556e-09 wkt2 = 1.370162094e-08 pkt2 = 1.006270608e-14
+ at = -1.366801920e+05 lat = 4.536918978e-02 wat = 4.479461574e-01 pat = -1.024259522e-7
+ ute = 5.281135183e+00 lute = -1.272068805e-06 wute = -1.992481667e-05 pute = 3.615217379e-12
+ ua1 = 2.108401453e-08 lua1 = -3.876942709e-15 wua1 = -6.067268780e-14 pua1 = 1.114053427e-20
+ ub1 = -1.991916571e-17 lub1 = 3.653306520e-24 wub1 = 5.649458055e-23 pub1 = -1.022593658e-29
+ uc1 = 1.395520365e-10 luc1 = -2.494192275e-17 wuc1 = -6.815233032e-16 puc1 = 1.218076210e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.31 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.01e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {2.912482682e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 4.216383911e-08 wvth0 = 9.582522211e-07 pvth0 = -1.519873042e-13
+ k1 = 6.328128152e-01 lk1 = 1.660547912e-08 wk1 = 8.566474836e-07 pk1 = -1.784633535e-13
+ k2 = -4.952030899e-02 lk2 = -1.613550659e-08 wk2 = -4.149752653e-07 pk2 = 8.490739304e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.209299539e+05 lvsat = -5.345859952e-03 wvsat = -1.734240469e-01 pvsat = 2.939609521e-8
+ ua = -2.749930259e-09 lua = 1.038028388e-17 wua = 3.298201498e-15 pua = -3.886174584e-22
+ ub = 1.134235365e-18 lub = 3.821505122e-25 wub = 3.723866645e-24 pub = -1.015639799e-30
+ uc = 1.421713030e-10 luc = -2.119158063e-17 wuc = -1.252025730e-16 puc = 2.827871754e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = -1.894861081e-02 lu0 = 6.403623539e-09 wu0 = 1.389197069e-07 pu0 = -2.507239841e-14
+ a0 = 0.0
+ keta = -3.322027448e-01 lketa = 5.459684708e-08 wketa = 1.646032064e-06 pketa = -3.497074405e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.302597604e+00 lags = -7.130573124e-09 wags = -2.106622352e-06 pags = 3.333054917e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {2.660304154e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.733865735e-08 wvoff = -1.192950639e-06 pvoff = 2.245369976e-13
+ nfactor = {4.313979636e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.629128598e-07 wnfactor = -1.063128940e-05 pnfactor = 2.178012994e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.965681037e-05 lcit = -5.127522413e-12 wcit = -1.488015443e-10 pcit = 2.959986660e-17
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 4.880749005e-01 leta0 = -7.269791517e-08 weta0 = -1.164232341e-06 peta0 = 2.072973797e-13
+ etab = 2.751040814e-02 letab = -9.085740771e-09 wetab = -3.519286268e-07 petab = 7.002604915e-14
+ dsub = 4.671587816e-01 ldsub = -3.326970032e-08 wdsub = 7.873879794e-07 pdsub = -1.264545095e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.031472604e+00 lpclm = 3.928270371e-07 wpclm = 7.160022495e-06 ppclm = -1.264459595e-12
+ pdiblc1 = 2.507556907e+00 lpdiblc1 = -2.865175596e-07 wpdiblc1 = -4.416965545e-06 ppdiblc1 = 8.378540705e-13
+ pdiblc2 = 5.120972761e-02 lpdiblc2 = -8.431818735e-09 wpdiblc2 = -1.216641397e-08 ppdiblc2 = 5.265502192e-15
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.207572646e-02 lalpha0 = -1.762600085e-09 walpha0 = -3.010684210e-08 palpha0 = 4.479044843e-15
+ alpha1 = 0.0
+ beta0 = 4.361902425e+01 lbeta0 = -2.039056867e-06 wbeta0 = -3.269428110e-05 pbeta0 = 3.875509605e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.162162527e+00 lkt1 = 1.608216943e-07 wkt1 = 3.313147246e-06 pkt1 = -6.227016078e-13
+ kt2 = -2.184832330e-01 lkt2 = 3.310075541e-08 wkt2 = 4.112218863e-07 pkt2 = -6.570465650e-14
+ at = 3.433907901e+05 lat = -4.613233941e-02 wat = -1.047623750e+00 pat = 1.826296721e-7
+ ute = -3.088572202e+00 lute = 3.231974223e-07 wute = 3.015374865e-06 pute = -7.571831279e-13
+ ua1 = -9.483701753e-10 lua1 = 3.224298162e-16 wua1 = -8.350988455e-17 pua1 = -4.077630403e-22
+ ub1 = 7.072011298e-19 lub1 = -2.780789993e-25 wub1 = 3.428536872e-24 pub1 = -1.115486532e-31
+ uc1 = 8.917805351e-11 luc1 = -1.534064158e-17 wuc1 = 2.394141033e-16 puc1 = -5.372304865e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.32 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 3.0e-06 wmax = 3.01e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.4255045+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.50407
+ k2 = -0.048314461
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 169790.0
+ ua = -1.1014364e-9
+ ub = 2.407218e-18
+ uc = 6.9010287e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0324708
+ a0 = 1.6844032
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.5385232
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11480431+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.41179304+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0067115
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.8823913e-5
+ alpha1 = 0.0
+ beta0 = 17.79575
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.2558
+ kt2 = -0.03478
+ at = 318480.0
+ ute = -1.261
+ ua1 = 2.0849e-9
+ ub1 = -2.0887e-18
+ uc1 = -4.6822e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.33 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 3.0e-06 wmax = 3.01e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.4255045+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.50407
+ k2 = -0.048314461
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 169790.0
+ ua = -1.1014364e-9
+ ub = 2.407218e-18
+ uc = 6.9010287e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0324708
+ a0 = 1.6844032
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.5385232
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11480431+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.41179304+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0067115
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.8823913e-5
+ alpha1 = 0.0
+ beta0 = 17.79575
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.2558
+ kt2 = -0.03478
+ at = 318480.0
+ ute = -1.261
+ ua1 = 2.0849e-9
+ ub1 = -2.0887e-18
+ uc1 = -4.6822e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.34 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 3.0e-06 wmax = 3.01e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.159485203e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.832521210e-8
+ k1 = 5.659864270e-01 lk1 = -2.483220221e-7
+ k2 = -7.820229238e-02 lk2 = 1.198681365e-7
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.021648881e+05 lvsat = -5.309027262e-1
+ ua = -9.666125508e-10 lua = -5.407245295e-16
+ ub = 2.261618390e-18 lub = 5.839417943e-25
+ uc = 4.900208962e-11 luc = 8.024487641e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.263164800e-02 lu0 = -6.450969888e-10
+ a0 = 1.546476241e+00 la0 = 5.531698615e-7
+ keta = 2.531445930e-01 lketa = -1.015261705e-6
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -6.721563730e-01 lags = 4.855551496e-06 pags = 2.067951531e-25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.116893377e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.249290797e-8
+ nfactor = {1.499306969e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.509833617e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.599213500e-01 leta0 = -3.205325663e-7
+ etab = -1.398762215e-01 letab = 2.802455739e-7
+ dsub = 7.769140535e-01 ldsub = -8.699555029e-07 wdsub = -1.084202172e-19
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.163260720e-01 lpclm = -6.547734436e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 5.433160520e-03 lpdiblc2 = 5.126908318e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.491070895e-05 lalpha0 = 4.160380748e-10 palpha0 = 2.524354897e-29
+ alpha1 = 0.0
+ beta0 = 1.410270304e+01 lbeta0 = 1.481133413e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.581524020e-01 lkt1 = 9.434543461e-9
+ kt2 = -3.330623020e-02 lkt2 = -5.910701160e-9
+ at = 5.956944909e+05 lat = -1.111796437e+0
+ ute = -1.311968710e+00 lute = 2.044151083e-7
+ ua1 = 1.940438390e-09 lua1 = 5.793777331e-16
+ ub1 = -1.675521700e-18 lub1 = -1.657092890e-24
+ uc1 = -4.012268080e-11 luc1 = -2.686828958e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.35 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 3.0e-06 wmax = 3.01e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.326549068e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.735351436e-9
+ k1 = 4.472904560e-01 lk1 = -9.671902834e-9
+ k2 = -1.386459694e-02 lk2 = -9.489233912e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -2.345360400e+03 lvsat = 8.134557942e-2
+ ua = -9.794756888e-10 lua = -5.148619043e-16
+ ub = 2.603000612e-18 lub = -1.024412999e-25
+ uc = 1.044661340e-10 luc = -3.127113122e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.686470711e-02 lu0 = -9.156085626e-9
+ a0 = 2.108717492e+00 la0 = -5.772723972e-7
+ keta = -3.188734160e-01 lketa = 1.348377042e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.429108537e+00 lags = 6.307482667e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.197246989e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.662989369e-9
+ nfactor = {7.287822219e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.198233694e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 5.345524140e-04 leta0 = -6.947108359e-11
+ etab = -5.117958520e-04 letab = 3.945973803e-11
+ dsub = -1.014849988e-01 ldsub = 8.961536316e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.784734320e-01 lpclm = -1.904308264e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.682604060e-03 lpdiblc2 = 1.065717714e-8
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.377584428e-04 lalpha0 = -1.925085218e-10
+ alpha1 = 0.0
+ beta0 = 2.213325482e+01 lbeta0 = -1.334893272e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.416056620e-01 lkt1 = -2.383433198e-8
+ kt2 = -5.170615880e-02 lkt2 = 3.108419528e-8
+ at = 7.956296400e+03 lat = 6.990997666e-2
+ ute = -1.315402400e+00 lute = 2.113188854e-7
+ ua1 = 1.752607400e-09 lua1 = 9.570307216e-16
+ ub1 = -1.933764000e-18 lub1 = -1.137870922e-24
+ uc1 = -1.878401720e-11 luc1 = -6.977180662e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.36 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 3.0e-06 wmax = 3.01e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.401908511e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.880473876e-9
+ k1 = 4.446743720e-01 lk1 = -7.028088343e-9
+ k2 = -1.791730762e-02 lk2 = -5.393564496e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -3.398586600e+04 lvsat = 1.133214744e-1
+ ua = -1.722316731e-09 lua = 2.358532534e-16
+ ub = 2.906508760e-18 lub = -4.091666343e-25
+ uc = 9.922047680e-11 luc = -2.596987005e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.644243643e-02 lu0 = 1.376661119e-9
+ a0 = 1.262899320e+00 la0 = 2.775114472e-7
+ keta = -3.624720340e-01 lketa = 1.788984676e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 3.324717717e+00 lags = -1.284954370e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.211672938e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.120875700e-9
+ nfactor = {1.327511996e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.931573843e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 9.312831720e-04 leta0 = -4.704071876e-10
+ etab = -8.540229139e-04 letab = 3.853144068e-10
+ dsub = 5.659857836e-01 ldsub = 2.216076589e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.183971320e-01 lpclm = 2.106465656e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 1.558901440e-02 lpdiblc2 = -2.386041153e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.642958181e-05 lalpha0 = 6.437389593e-11
+ alpha1 = 0.0
+ beta0 = 1.781694444e+01 lbeta0 = 3.027169998e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.721443720e-01 lkt1 = 7.028088343e-9
+ kt2 = -1.688975120e-02 lkt2 = -4.101266237e-9
+ at = 8.251676640e+04 lat = -5.440834324e-3
+ ute = -6.610568000e-01 lute = -4.499627779e-7
+ ua1 = 5.155208156e-09 lua1 = -2.481637602e-15
+ ub1 = -6.116866440e-18 lub1 = 3.089572404e-24
+ uc1 = -1.775098688e-10 luc1 = 9.063653901e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.37 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 3.0e-06 wmax = 3.01e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {5.006786576e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.376554787e-8
+ k1 = 2.648519899e-01 lk1 = 8.478921996e-8
+ k2 = 2.687543262e-02 lk2 = -2.826473766e-08 pk2 = -1.615587134e-27
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.928791329e+05 lvsat = -2.515794073e-3
+ ua = -1.994271278e-10 lua = -5.417341782e-16
+ ub = 1.602399052e-18 lub = 2.567117822e-25
+ uc = 4.924934511e-11 luc = -4.546102142e-19
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 4.344405666e-02 lu0 = -7.304366173e-9
+ a0 = 2.131485262e+00 la0 = -1.659885345e-7
+ keta = 9.924730893e-03 lketa = -1.124732059e-08 pketa = 8.077935669e-28
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.650585984e+00 lags = -4.301427074e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.115896756e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.305438449e-10
+ nfactor = {2.482255469e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.545366745e-9
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -8.534188585e-03 leta0 = 4.362662692e-09 weta0 = -2.911675756e-22 peta0 = 1.443615457e-28
+ etab = 1.919533138e-02 letab = -9.851885895e-09 wetab = -3.705769144e-22 petab = 4.985600921e-28
+ dsub = 1.767026398e+00 ldsub = -3.916436790e-07 wdsub = -2.168404345e-19 pdsub = 5.169878828e-26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.230923648e-01 lpclm = 3.628202854e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 4.472925600e-03 lpdiblc2 = 3.289833789e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.871020363e-03 lalpha0 = 1.011327949e-09 walpha0 = -2.646977960e-23 palpha0 = 2.524354897e-29
+ alpha1 = 0.0
+ beta0 = 1.673611267e+01 lbeta0 = 3.579042699e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.452144880e-01 lkt1 = -6.722310427e-9
+ kt2 = -3.153915520e-02 lkt2 = 3.378719445e-9
+ at = 8.798797040e+04 lat = -8.234431086e-3
+ ute = -1.386565440e+00 lute = -7.951806634e-8
+ ua1 = 5.888173480e-10 lua1 = -1.500384559e-16
+ ub1 = -2.000359616e-19 lub1 = 6.843876199e-26 pub1 = 5.605193857e-45
+ uc1 = 3.142940240e-11 luc1 = -1.604785287e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.38 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.0e-06 wmax = 3.01e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {5.486027986e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -4.625457901e-8
+ k1 = 3.119744075e-01 lk1 = 7.250911793e-8
+ k2 = 3.291655585e-02 lk2 = -2.983905438e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.749921224e+05 lvsat = 2.145560871e-3
+ ua = -2.327078853e-09 lua = 1.273186146e-17
+ ub = 2.595219338e-18 lub = -2.017184277e-27
+ uc = 7.068153865e-11 luc = -6.039839851e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 1.056213734e-02 lu0 = 1.264662003e-9
+ a0 = 5.563950352e+00 la0 = -1.060488937e-6
+ keta = 1.784573743e-01 lketa = -5.516692745e-08 wketa = 1.355252716e-20 pketa = -3.231174268e-27
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -3.108141429e+00 lags = 8.099816563e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.605030774e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.297737638e-8
+ nfactor = {5.524009374e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.064654578e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.877591979e-01 leta0 = 5.106870013e-08 weta0 = -3.388131789e-21 peta0 = -2.423380701e-27
+ etab = -2.894663676e-02 letab = 2.693911001e-9
+ dsub = 7.013384757e-02 ldsub = 5.056651973e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 7.735704401e-01 lpclm = -1.071725579e-7
+ pdiblc1 = -1.262852704e+00 lpdiblc1 = 4.307334147e-7
+ pdiblc2 = 3.012042571e-02 lpdiblc2 = -3.393904741e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.998680363e-03 lalpha0 = -1.039516060e-9
+ alpha1 = 0.0
+ beta0 = 3.542783069e+01 lbeta0 = -1.292019018e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.853489143e-01 lkt1 = -2.232327894e-8
+ kt2 = -9.689317143e-03 lkt2 = -2.315348353e-9
+ at = 1.812296571e+04 lat = 9.972389135e-3
+ ute = -1.604568571e+00 lute = -2.270645029e-8
+ ua1 = 1.164863914e-10 lua1 = -2.694900861e-17 wua1 = 6.310887242e-30 pua1 = -1.504632769e-36
+ ub1 = -3.955258229e-19 lub1 = 1.193834198e-25
+ uc1 = -9.597171486e-11 luc1 = 1.715287829e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.39 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.0e-06 wmax = 3.01e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.018908126e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 6.337130033e-07 wvth0 = 9.778192776e-06 pvth0 = -1.863723543e-12
+ k1 = 9.288567333e-01 lk1 = -4.506865337e-8
+ k2 = 9.463316632e-01 lk2 = -2.039359738e-07 wk2 = -3.296622325e-06 pk2 = 6.283362151e-13
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 6.272560921e+06 lvsat = -1.160051052e+00 wvsat = -1.768472599e+01 pvsat = 3.370708774e-6
+ ua = -8.710916099e-09 lua = 1.229491240e-15 wua = 2.054720817e-14 pua = -3.916297878e-21
+ ub = 2.688314546e-17 lub = -4.631295903e-24 wub = -7.078446705e-23 pub = 1.349151942e-29
+ uc = 9.890325989e-11 luc = -1.141889992e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = -9.967044928e-02 lu0 = 2.227499301e-08 wu0 = 3.725004548e-07 pu0 = -7.099858669e-14
+ a0 = 0.0
+ keta = 2.366400884e-01 lketa = -6.625655277e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 5.745820000e-01 lags = 1.080545708e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.462345920e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.025780305e-8
+ nfactor = {-7.839818213e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.555444659e-05 wnfactor = 2.287087575e-04 pnfactor = -4.359188918e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.176666667e-05 lcit = 5.101726667e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 8.573448585e-02 leta0 = -1.059196002e-9
+ etab = -9.411059882e-02 letab = 1.511416217e-8
+ dsub = 7.392677026e-01 ldsub = -7.697039304e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 4.429187333e-01 lpclm = -4.415034257e-8
+ pdiblc1 = 9.811229760e-01 lpdiblc1 = 3.031650054e-9
+ pdiblc2 = 4.700520600e-02 lpdiblc2 = -6.612143864e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.671274608e-03 lalpha0 = -2.147125235e-10
+ alpha1 = 0.0
+ beta0 = 3.232039411e+01 lbeta0 = -6.997416058e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.719086667e-02 lkt1 = -5.437420281e-8
+ kt2 = -7.637140667e-02 lkt2 = 1.039425791e-8
+ at = -1.865152667e+04 lat = 1.698160738e-2
+ ute = -2.046506000e+00 lute = 6.152682360e-8
+ ua1 = -9.772298800e-10 lua1 = 1.815133127e-16 wua1 = 2.524354897e-29 pua1 = -6.018531076e-36
+ ub1 = 1.892049633e-18 lub1 = -3.166284621e-25 wub1 = 1.880790961e-37 pub1 = 2.242077543e-44
+ uc1 = 1.719158080e-10 luc1 = -3.390648356e-17 wuc1 = 6.310887242e-30 puc1 = 2.256949154e-36
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.40 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 1.65e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.300018434e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = -1.296876436e-8
+ k1 = 4.709090789e-01 wk1 = 9.562449016e-8
+ k2 = -3.781288124e-02 wk2 = -3.028288049e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.348455007e+05 wvsat = 1.007677053e-1
+ ua = -1.240718153e-09 wua = 4.016398280e-16
+ ub = 2.717296924e-18 wub = -8.941590880e-25
+ uc = 1.220174343e-10 wuc = -1.528540604e-16
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.620449933e-02 wu0 = -1.076668206e-8
+ a0 = 1.421338942e+00 wa0 = 7.585852476e-7
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.957823058e-01 wags = 1.232497797e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.199962492e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = 1.497173544e-8
+ nfactor = {9.409661708e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 1.357699901e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.801851852e-07 wcit = 1.637966601e-11
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 5.737234637e-03 wpdiblc2 = 2.809440314e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.551688192e-05 walpha0 = 9.536320173e-12
+ alpha1 = 0.0
+ beta0 = 1.779846172e+01 wbeta0 = -7.819652553e-9
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.537210522e-01 wkt1 = -5.994957759e-9
+ kt2 = -3.298051733e-02 wkt2 = -5.189078192e-9
+ at = 6.141336389e+05 wat = -8.525616158e-1
+ ute = -1.352110170e+00 wute = 2.627298428e-7
+ ua1 = 2.222701293e-09 wua1 = -3.973706974e-16
+ ub1 = -2.796110263e-18 wub1 = 2.039923605e-24
+ uc1 = -1.720587230e-10 wuc1 = 3.611388762e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.41 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1.65e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.300018434e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = -1.296876436e-8
+ k1 = 4.709090789e-01 wk1 = 9.562449016e-8
+ k2 = -3.781288124e-02 wk2 = -3.028288049e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.348455007e+05 wvsat = 1.007677053e-1
+ ua = -1.240718153e-09 wua = 4.016398280e-16
+ ub = 2.717296924e-18 wub = -8.941590880e-25
+ uc = 1.220174343e-10 wuc = -1.528540604e-16
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.620449933e-02 wu0 = -1.076668206e-8
+ a0 = 1.421338942e+00 wa0 = 7.585852476e-7
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.957823058e-01 wags = 1.232497797e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.199962492e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = 1.497173544e-8
+ nfactor = {9.409661708e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 1.357699901e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.801851852e-07 wcit = 1.637966601e-11
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 5.737234637e-03 wpdiblc2 = 2.809440314e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.551688192e-05 walpha0 = 9.536320173e-12
+ alpha1 = 0.0
+ beta0 = 1.779846172e+01 wbeta0 = -7.819652553e-9
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.537210522e-01 wkt1 = -5.994957759e-9
+ kt2 = -3.298051733e-02 wkt2 = -5.189078192e-9
+ at = 6.141336389e+05 wat = -8.525616158e-1
+ ute = -1.352110170e+00 wute = 2.627298428e-7
+ ua1 = 2.222701293e-09 wua1 = -3.973706974e-16
+ ub1 = -2.796110263e-18 wub1 = 2.039923605e-24
+ uc1 = -1.720587230e-10 wuc1 = 3.611388762e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.42 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1.65e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.274691780e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.015750782e-08 wvth0 = -3.322154460e-08 pvth0 = 8.122580045e-14
+ k1 = 5.171336285e-01 lk1 = -1.853881787e-07 wk1 = 1.408743724e-07 pk1 = -1.814791776e-13
+ k2 = -6.818409211e-02 lk2 = 1.218067783e-07 wk2 = -2.888898322e-08 pk2 = -5.590364362e-15
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.373270198e+05 lvsat = -4.110123804e-01 wvsat = 1.869697189e-01 pvsat = -3.457217957e-7
+ ua = -1.099315171e-09 lua = -5.671108029e-16 wua = 3.826679092e-16 pua = 7.608877742e-23
+ ub = 2.576465292e-18 lub = 5.648193414e-25 wub = -9.079082680e-25 pub = 5.514246131e-32
+ uc = 1.125295329e-10 luc = 3.805217733e-17 wuc = -1.831909119e-16 puc = 1.216689767e-22
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.670739371e-02 lu0 = -2.016908204e-09 wu0 = -1.175302411e-08 pu0 = 3.955823412e-15
+ a0 = 1.047262819e+00 la0 = 1.500269699e-06 wa0 = 1.439556785e-06 pa0 = -2.731104446e-12
+ keta = 3.337510490e-01 lketa = -1.338541957e-06 wketa = -2.324408068e-07 pketa = 9.322270998e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -1.104604928e+00 lags = 6.418513039e-06 wags = 1.247030275e-06 pags = -4.507034054e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.211150345e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.487000252e-09 wvoff = 2.718041053e-08 pvoff = -4.896411234e-14
+ nfactor = {5.147423325e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.709413326e-06 wnfactor = 2.839139813e-06 pnfactor = -5.941462908e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.801851852e-07 wcit = 1.637966601e-11
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.599213500e-01 leta0 = -3.205325663e-7
+ etab = -1.398851638e-01 letab = 2.802814380e-07 wetab = 2.578650492e-11 petab = -1.034193566e-16
+ dsub = 8.431688943e-01 ldsub = -1.135677168e-06 wdsub = -1.910557717e-07 pdsub = 7.662482781e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.743083584e-01 lpclm = -2.980211020e-07 wpclm = -1.672006200e-07 ppclm = 6.705748067e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 7.779200477e-03 lpdiblc2 = -8.189508199e-09 wpdiblc2 = -6.765158123e-09 ppdiblc2 = 3.839988449e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -9.161597834e-05 lalpha0 = 5.098790493e-10 walpha0 = 7.700865005e-11 palpha0 = -2.706045262e-16
+ alpha1 = 0.0
+ beta0 = 1.379054365e+01 lbeta0 = 1.607415620e-05 wbeta0 = 9.001584240e-07 pbeta0 = -3.641536874e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.711828820e-01 lkt1 = 7.003241452e-08 wkt1 = 3.757534366e-08 pkt1 = -1.747430509e-13
+ kt2 = -3.066048253e-02 lkt2 = -9.304731580e-09 wkt2 = -7.629410267e-09 pkt2 = 9.787195820e-15
+ at = 1.195929297e+06 lat = -2.333349666e+00 wat = -1.730867099e+00 pat = 3.522531969e-6
+ ute = -1.391201477e+00 lute = 1.567795937e-07 wute = 2.284795681e-07 pute = 1.373641519e-13
+ ua1 = 2.008574143e-09 lua1 = 8.587783479e-16 wua1 = -1.964796629e-16 pua1 = -8.056935830e-22
+ ub1 = -2.402689567e-18 lub1 = -1.577853043e-24 wub1 = 2.096897620e-24 pub1 = -2.284999834e-31
+ uc1 = -2.406713929e-10 luc1 = 2.751779741e-16 wuc1 = 5.783122937e-16 puc1 = -8.709957083e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.43 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1.65e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.331664104e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.297347584e-09 wvth0 = -1.474997343e-09 pvth0 = 1.739619253e-14
+ k1 = 4.346869044e-01 lk1 = -1.962079521e-08 wk1 = 3.634423158e-08 pk1 = 2.868912349e-14
+ k2 = -2.014123538e-03 lk2 = -1.123456048e-08 wk2 = -3.417261763e-08 pk2 = 5.032910968e-15
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -5.988110418e+03 lvsat = 7.819702044e-02 wvsat = 1.050441609e-02 pvsat = 9.079342099e-9
+ ua = -1.298002379e-09 lua = -1.676303024e-16 wua = 9.185194890e-16 pua = -1.001294409e-21
+ ub = 3.021893421e-18 lub = -3.307584541e-25 wub = -1.207940249e-24 pub = 6.583867616e-31
+ uc = 1.567189014e-10 luc = -5.079496688e-17 wuc = -1.506786927e-16 puc = 5.629990870e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.968348320e-02 lu0 = -8.000633730e-09 wu0 = -8.128363673e-09 pu0 = -3.331918858e-15
+ a0 = 2.001871513e+00 la0 = -4.190665418e-07 wa0 = 3.081064060e-07 pa0 = -4.562103148e-13
+ keta = -3.963454436e-01 lketa = 1.293900508e-07 wketa = 2.234022123e-07 pketa = 1.570912563e-14
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.761241475e+00 lags = 6.564422623e-07 wags = -9.577551442e-07 pags = -7.409249040e-14
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.206054905e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.462511108e-09 wvoff = 2.539894532e-09 pvoff = 5.781091358e-16
+ nfactor = {1.003696977e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.263211185e-07 wnfactor = -7.927579322e-07 pnfactor = 1.360830698e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.420580333e-06 lcit = 1.154163848e-11 wcit = 3.293295648e-11 pcit = -3.328204582e-17
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 4.974350190e-04 leta0 = 5.157150855e-12 weta0 = 1.070335762e-10 peta0 = -2.152017083e-16
+ etab = -4.929468368e-04 letab = 1.944653690e-11 wetab = -5.435396264e-11 petab = 5.771106745e-17
+ dsub = -4.780043780e-01 ldsub = 1.520673814e-06 wdsub = 1.085750108e-06 pdsub = -1.800897623e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.024367314e-01 lpclm = -3.545760089e-07 wpclm = -6.910176839e-08 ppclm = 4.733372556e-13
+ pdiblc1 = 0.39
+ pdiblc2 = -4.234928741e-03 lpdiblc2 = 1.596610001e-08 wpdiblc2 = 1.994774346e-08 ppdiblc2 = -1.530907543e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.776641528e-04 lalpha0 = -2.325955823e-10 walpha0 = -1.150741005e-10 palpha0 = 1.155970520e-16
+ alpha1 = 0.0
+ beta0 = 2.272318965e+01 lbeta0 = -1.885821843e-06 wbeta0 = -1.701165583e-06 pbeta0 = 1.588685175e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.121895370e-01 lkt1 = -4.857960489e-08 wkt1 = -8.482580879e-08 pkt1 = 7.135670623e-14
+ kt2 = -5.180815652e-02 lkt2 = 3.321478175e-08 wkt2 = 2.941257314e-10 pkt2 = -6.143865658e-15
+ at = -5.134559428e+03 lat = 8.150932334e-02 wat = 3.774944641e-02 pat = -3.344845605e-8
+ ute = -1.506959057e+00 lute = 3.895217836e-07 wute = 5.523823529e-07 pute = -5.138747874e-13
+ ua1 = 1.360754122e-09 lua1 = 2.161285281e-15 wua1 = 1.129967705e-15 pua1 = -3.472648661e-21
+ ub1 = -1.784915633e-18 lub1 = -2.819949314e-24 wub1 = -4.292265925e-25 pub1 = 4.850525357e-30
+ uc1 = -7.648668546e-11 luc1 = -5.493179869e-17 wuc1 = 1.663942993e-16 puc1 = -4.279338887e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.44 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 1.65e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.296327147e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.273805270e-09 wvth0 = 3.044596999e-08 pvth0 = -1.486313706e-14
+ k1 = 4.480041693e-01 lk1 = -3.307922308e-08 wk1 = -9.601969874e-09 pk1 = 7.512235469e-14
+ k2 = -1.005872965e-02 lk2 = -3.104681549e-09 wk2 = -2.266138838e-08 pk2 = -6.600337309e-15
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -3.604682031e+04 lvsat = 1.085743527e-01 wvsat = 5.943070909e-03 pvsat = 1.368903754e-8
+ ua = -2.361542113e-09 lua = 9.071829528e-16 wua = 1.843302270e-15 pua = -1.935879888e-21
+ ub = 3.627576490e-18 lub = -9.428617641e-25 wub = -2.079306961e-24 pub = 1.538989961e-30
+ uc = 1.755322420e-10 luc = -6.980772890e-17 wuc = -2.200564217e-16 puc = 1.264130417e-22
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.514450765e-02 lu0 = 6.692454956e-09 wu0 = 3.742772324e-09 pu0 = -1.532888890e-14
+ a0 = 4.024488986e-01 la0 = 1.197309952e-06 wa0 = 2.481237858e-06 pa0 = -2.652376960e-12
+ keta = -5.159129463e-01 lketa = 2.502249691e-07 wketa = 4.424698867e-07 pketa = -2.056806661e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 3.372605206e+00 lags = -9.720019247e-07 wags = -1.380907569e-07 pags = -9.024453202e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.369106805e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.994053618e-08 wvoff = 4.539841727e-08 pvoff = -4.273471394e-14
+ nfactor = {3.509115586e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.386026062e-06 wnfactor = 2.816173851e-06 pnfactor = -2.286355762e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 4.138029529e-03 leta0 = -3.674027661e-09 weta0 = -9.247134133e-09 peta0 = 9.238120179e-15
+ etab = -8.856597526e-04 letab = 4.163222095e-10 wetab = 9.122956984e-11 petab = -8.941565048e-17
+ dsub = 1.054005179e+00 ldsub = -2.757504423e-08 wdsub = -1.407277128e-06 pdsub = 7.185557018e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -3.626371609e-01 lpclm = 3.175476667e-07 wpclm = 7.043027593e-07 ppclm = -3.082653601e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 8.083046745e-03 lpdiblc2 = 3.517553981e-09 wpdiblc2 = 2.164458363e-08 ppdiblc2 = -1.702390211e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.024104834e-05 lalpha0 = 2.755620706e-11 walpha0 = -1.057452626e-10 palpha0 = 1.061693285e-16
+ alpha1 = 0.0
+ beta0 = 1.853258551e+01 lbeta0 = 2.349202699e-06 wbeta0 = -2.063658386e-06 pbeta0 = 1.955020401e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.764485346e-01 lkt1 = 1.636053805e-08 wkt1 = 1.241169847e-08 pkt1 = -2.691151860e-14
+ kt2 = -2.545105218e-02 lkt2 = 6.578292103e-09 wkt2 = 2.468779558e-08 pkt2 = -3.079610841e-14
+ at = 9.031797590e+04 lat = -1.495500887e-02 wat = -2.249595778e-02 pat = 2.743554943e-8
+ ute = -2.125793237e-01 lute = -9.185783745e-07 wute = -1.293252074e-06 pute = 1.351323365e-12
+ ua1 = 8.124323333e-09 lua1 = -4.673977764e-15 wua1 = -8.561888981e-15 pua1 = 6.321941706e-21
+ ub1 = -1.060259529e-17 lub1 = 6.091197749e-24 wub1 = 1.293527200e-23 pub1 = -8.655636925e-30
+ uc1 = -2.780388627e-10 luc1 = 1.487568316e-16 wuc1 = 2.898904333e-16 puc1 = -1.675985819e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.45 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 1.65e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.909045710e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.901160454e-08 wvth0 = 2.818504486e-08 pvth0 = -1.370870869e-14
+ k1 = 1.796413484e-01 lk1 = 1.039468333e-07 wk1 = 2.457176665e-07 pk1 = -5.524385163e-14
+ k2 = 5.994307163e-02 lk2 = -3.884760128e-08 wk2 = -9.535549725e-08 pk2 = 3.051727468e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.406173147e+05 lvsat = 1.836964531e-02 wvsat = 1.507047920e-01 pvsat = -6.022629727e-8
+ ua = 1.255936096e-09 lua = -9.399014207e-16 wua = -4.196758162e-15 pua = 1.148174969e-21
+ ub = 4.733019163e-19 lub = 6.677108333e-25 wub = 3.255920957e-24 pub = -1.185177414e-30
+ uc = 2.303437926e-11 luc = 8.057679817e-18 wuc = 7.559478627e-17 puc = -2.454646515e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 5.858375227e-02 lu0 = -1.038162335e-08 wu0 = -4.365758324e-08 pu0 = 8.873732653e-15
+ a0 = 4.077171639e+00 la0 = -6.790034786e-07 wa0 = -5.610678522e-06 pa0 = 1.479355543e-12
+ keta = -1.089994895e-02 lketa = -7.634667343e-09 wketa = 6.005108802e-08 pketa = -1.041762753e-14
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 3.000201174e+00 lags = -7.818524259e-07 wags = -3.891817843e-06 pags = 1.014207730e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-8.555414408e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.282111335e-09 wvoff = -7.507736035e-08 pvoff = 1.878021811e-14
+ nfactor = {3.237936554e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -8.808890083e-08 wnfactor = -2.179119760e-06 pnfactor = 2.642411557e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.092102504e-05 lcit = -3.023275384e-12 wcit = -1.707416385e-11 pcit = 8.718068061e-18
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -2.112008228e-02 leta0 = 9.222764226e-09 weta0 = 3.629331234e-08 peta0 = -1.401483179e-14
+ etab = 3.109951072e-02 letab = -1.591530583e-08 wetab = -3.432748675e-08 petab = 1.748478090e-14
+ dsub = 1.867905010e+00 ldsub = -4.431522980e-07 wdsub = -2.908986079e-07 pdsub = 1.485328292e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.845129998e-01 lpclm = -6.394720537e-08 wpclm = -4.654806140e-07 ppclm = 2.890260304e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 7.094249450e-03 lpdiblc2 = 4.022433880e-09 wpdiblc2 = -7.558980520e-09 ppdiblc2 = -2.112562252e-15
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.646910139e-03 lalpha0 = 1.389403603e-09 walpha0 = 2.237394554e-09 palpha0 = -1.090237862e-15
+ alpha1 = 0.0
+ beta0 = 1.484878072e+01 lbeta0 = 4.230153425e-06 wbeta0 = 5.442404770e-06 pbeta0 = -1.877575446e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.169360360e-01 lkt1 = -1.402654375e-08 wkt1 = -8.154515824e-08 pkt1 = 2.106285243e-14
+ kt2 = -1.330754297e-02 lkt2 = 3.778162990e-10 wkt2 = -5.257358861e-08 pkt2 = 8.653554357e-15
+ at = 6.201579623e+04 lat = -5.039159296e-04 wat = 7.489466004e-02 pat = -2.229210003e-8
+ ute = -1.549745346e+00 lute = -2.358214037e-07 wute = 4.705537347e-07 pute = 4.507241187e-13
+ ua1 = -7.840437999e-10 lua1 = -1.253655055e-16 wua1 = 3.958851049e-15 pua1 = -7.114815344e-23
+ ub1 = 1.553314475e-18 lub1 = -1.156097782e-25 wub1 = -5.056048986e-24 pub1 = 5.307315730e-31
+ uc1 = 1.028517127e-10 luc1 = -4.572589614e-17 wuc1 = -2.059569450e-16 puc1 = 8.558108948e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.46 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.65e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {5.564652574e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -4.609671942e-08 wvth0 = -2.267257935e-08 pvth0 = -4.552118188e-16
+ k1 = 3.856932875e-01 lk1 = 5.024969793e-08 wk1 = -2.125794483e-07 pk1 = 6.418837648e-14
+ k2 = -8.770342405e-03 lk2 = -2.094088558e-08 wk2 = 1.202104242e-07 pk2 = -2.565920444e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.852664659e+05 lvsat = -1.932592348e-02 wvsat = -3.179926105e-01 pvsat = 6.191624584e-8
+ ua = -2.630988136e-09 lua = 7.303103427e-17 wua = 8.763680030e-16 pua = -1.738817097e-22
+ ub = 3.492522958e-18 lub = -1.190981702e-25 wub = -2.587509583e-24 pub = 3.376205850e-31
+ uc = 6.952147748e-11 luc = -4.056857978e-18 wuc = 3.345210410e-18 puc = -5.718225678e-24
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 1.664838189e-02 lu0 = 5.467341739e-10 wu0 = -1.755059909e-08 pu0 = 2.070252584e-15
+ a0 = 5.478677864e+00 la0 = -1.044236001e-06 wa0 = 2.458960098e-07 pa0 = -4.686777947e-14
+ keta = 1.775565937e-01 lketa = -5.674644235e-08 wketa = 2.597535920e-09 pketa = 4.554768147e-15
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -3.253524957e+00 lags = 8.478686038e-07 wags = 4.192352116e-07 pags = -1.092526961e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.429053962e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 8.663624962e-09 wvoff = -5.074555358e-08 pvoff = 1.243934926e-14
+ nfactor = {2.358253406e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.411565275e-07 wnfactor = -5.207446472e-06 pnfactor = 1.053423097e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.614651799e-05 lcit = 4.030526329e-12 wcit = 6.097915660e-11 pcit = -1.162262725e-17
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.831542407e-01 leta0 = 5.144886590e-08 weta0 = -1.327908505e-08 peta0 = -1.096265031e-15
+ etab = -8.724984675e-02 letab = 1.492653672e-08 wetab = 1.681260515e-07 petab = -3.527461117e-14
+ dsub = -2.794295123e-01 ldsub = 1.164430784e-07 wdsub = 1.008018383e-06 pdsub = -1.899649385e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 4.224245586e-02 lpclm = 2.524849837e-08 wpclm = 2.108893942e-06 ppclm = -3.818559788e-13
+ pdiblc1 = -1.253661990e+00 lpdiblc1 = 4.283383147e-07 wpdiblc1 = -2.650280129e-08 ppdiblc1 = 6.906630016e-15
+ pdiblc2 = 5.680678936e-02 lpdiblc2 = -8.932654022e-09 wpdiblc2 = -7.695413254e-08 ppdiblc2 = 1.597181436e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 8.286584906e-03 lalpha0 = -1.459865205e-09 walpha0 = -6.597515935e-09 palpha0 = 1.212139812e-15
+ alpha1 = 0.0
+ beta0 = 3.675506836e+01 lbeta0 = -1.478625132e-06 wbeta0 = -3.827288887e-06 pbeta0 = 5.381067209e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.897079533e-01 lkt1 = -2.112218209e-08 wkt1 = 1.256994289e-08 pkt1 = -3.463542920e-15
+ kt2 = 1.834263369e-02 lkt2 = -7.870219739e-09 wkt2 = -8.083433502e-08 pkt2 = 1.601830487e-14
+ at = 4.297921589e+04 lat = 4.457016907e-03 wat = -7.167672583e-02 pat = 1.590440313e-8
+ ute = -4.555707811e+00 lute = 5.475324147e-07 wute = 8.510052667e-06 pute = -1.644369303e-12
+ ua1 = -5.302841914e-09 lua1 = 1.052233283e-15 wua1 = 1.562744607e-14 pua1 = -3.111984015e-21
+ ub1 = 4.158888082e-18 lub1 = -7.946222602e-25 wub1 = -1.313333566e-23 pub1 = 2.635672479e-30
+ uc1 = -2.025037471e-10 luc1 = 3.384973666e-17 wuc1 = 3.072010946e-16 puc1 = -4.814789564e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.47 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.65e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {6.364032786e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -6.133290625e-08 wvth0 = -7.624459567e-07 pvth0 = 1.405455939e-13
+ k1 = 6.552366842e-01 lk1 = -1.125273490e-09 wk1 = 7.890244545e-07 pk1 = -1.267173274e-13
+ k2 = -1.283558755e-01 lk2 = 1.852117018e-09 wk2 = -1.975996037e-07 pk2 = 3.491538688e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.284493351e+05 lvsat = 1.056342164e-02 wvsat = 3.274137990e-02 pvsat = -4.933652737e-9
+ ua = -1.472883926e-09 lua = -1.477036282e-16 wua = -3.247433018e-16 pua = 5.505010503e-23
+ ub = 3.354447214e-18 lub = -9.278093336e-26 wub = -2.935936356e-24 pub = 4.040307277e-31
+ uc = 1.576324003e-10 luc = -2.085079987e-17 wuc = -1.693542858e-16 puc = 2.719829830e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 4.020213322e-02 lu0 = -3.942610829e-09 wu0 = -3.084311770e-08 pu0 = 4.603806631e-15
+ a0 = 0.0
+ keta = 1.782666324e-01 lketa = -5.688177573e-08 wketa = 1.683286164e-07 pketa = -2.703357580e-14
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 9.138102328e-01 lags = 5.357451661e-08 wags = -9.782154936e-07 pags = 1.571014083e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.782223708e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.539504033e-08 wvoff = 9.224155843e-08 pvoff = -1.481399428e-14
+ nfactor = {-2.025308647e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 9.766634548e-07 wnfactor = 8.476120878e-06 pnfactor = -1.554664840e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.176666667e-05 lcit = 5.101726667e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.276635068e-01 leta0 = -7.792996772e-09 weta0 = -1.209086214e-07 peta0 = 1.941792459e-14
+ etab = -5.677613555e-02 letab = 9.118247369e-09 wetab = -1.076595250e-07 petab = 1.729011972e-14
+ dsub = 7.142604469e-01 ldsub = -7.295422777e-08 wdsub = 7.211217301e-08 pdsub = -1.158121499e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.105834819e-01 lpclm = -6.837301201e-09 wpclm = 6.699735477e-07 ppclm = -1.075977518e-13
+ pdiblc1 = 9.596779776e-01 lpdiblc1 = 6.475716800e-09 wpdiblc1 = 6.183986967e-08 ppdiblc1 = -9.931483070e-15
+ pdiblc2 = 3.192759369e-02 lpdiblc2 = -4.190679327e-09 wpdiblc2 = 4.347855673e-08 ppdiblc2 = -6.982656210e-15
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.195456641e-03 lalpha0 = -2.988961581e-10 walpha0 = -1.511557521e-09 palpha0 = 2.427561378e-16
+ alpha1 = 0.0
+ beta0 = 3.453257360e+01 lbeta0 = -1.055017631e-06 wbeta0 = -6.379151365e-06 pbeta0 = 1.024491709e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -4.848733089e-03 lkt1 = -5.635634947e-08 wkt1 = -3.559039349e-08 pkt1 = 5.715817195e-15
+ kt2 = -8.343745858e-02 lkt2 = 1.152906585e-08 wkt2 = 2.037602060e-08 pkt2 = -3.272388909e-15
+ at = -4.457722480e+04 lat = 2.114527450e-02 wat = 7.476063943e-02 pat = -1.200655869e-8
+ ute = -1.788115133e+00 lute = 2.002925041e-08 wute = -7.451088228e-07 pute = 1.196644769e-13
+ ua1 = 5.647140083e-10 lua1 = -6.612287574e-17 wua1 = -4.446426494e-15 pua1 = 7.140960949e-22
+ ub1 = 3.609033075e-19 lub1 = -7.072636218e-26 wub1 = 4.415290103e-24 pub1 = -7.090955905e-31
+ uc1 = 5.164424245e-11 luc1 = -1.459087014e-17 wuc1 = 3.468211000e-16 puc1 = -5.569946866e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.48 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 1e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.4215457+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.53326
+ k2 = -0.057558508
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200550.0
+ ua = -9.7883322e-10
+ ub = 2.1342701e-18
+ uc = 2.2350587e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0291842
+ a0 = 1.9159663
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.576146
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.8262398+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0075691
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.1734937e-5
+ alpha1 = 0.0
+ beta0 = 17.793363
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25763
+ kt2 = -0.036364
+ at = 58230.0
+ ute = -1.1808
+ ua1 = 1.9636e-9
+ ub1 = -1.466e-18
+ uc1 = 6.3418e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.49 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.4215457+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.53326
+ k2 = -0.057558508
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200550.0
+ ua = -9.7883322e-10
+ ub = 2.1342701e-18
+ uc = 2.2350587e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0291842
+ a0 = 1.9159663
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.576146
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.8262398+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0075691
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.1734937e-5
+ alpha1 = 0.0
+ beta0 = 17.793363
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25763
+ kt2 = -0.036364
+ at = 58230.0
+ ute = -1.1808
+ ua1 = 1.9636e-9
+ ub1 = -1.466e-18
+ uc1 = 6.3418e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.50 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.058074269e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.311991805e-8
+ k1 = 6.089892490e-01 lk1 = -3.037197260e-7
+ k2 = -8.702084314e-02 lk2 = 1.181616413e-7
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.592386156e+05 lvsat = -6.364365617e-1
+ ua = -8.498006729e-10 lua = -5.174979333e-16
+ ub = 1.984473463e-18 lub = 6.007743906e-25
+ uc = -6.918132389e-12 luc = 1.173851260e-16 puc = 2.350988702e-38
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.904396065e-02 lu0 = 5.624439371e-10
+ a0 = 1.985910349e+00 la0 = -2.805176033e-7
+ keta = 1.821905190e-01 lketa = -7.306932955e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.914922392e-01 lags = 3.479749922e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.033923399e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.743952297e-8
+ nfactor = {2.365972934e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.164653709e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.599213500e-01 leta0 = -3.205325663e-7
+ etab = -1.398683500e-01 letab = 2.802140045e-7
+ dsub = 7.185930317e-01 ldsub = -6.360532128e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.652869910e-01 lpclm = 1.392199939e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 3.368051830e-03 lpdiblc2 = 1.684872379e-8
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -4.140331570e-05 lalpha0 = 3.334342763e-10 palpha0 = 4.930380658e-32
+ alpha1 = 0.0
+ beta0 = 1.437748228e+01 lbeta0 = 1.369973122e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.466822830e-01 lkt1 = -4.390691380e-8
+ kt2 = -3.563515750e-02 lkt2 = -2.923095730e-9
+ at = 6.733600740e+04 lat = -3.652055328e-2
+ ute = -1.242223830e+00 lute = 2.463464126e-7
+ ua1 = 1.880461690e-09 lua1 = 3.334345061e-16
+ ub1 = -1.035430010e-18 lub1 = -1.726844002e-24
+ uc1 = 1.364109229e-10 luc1 = -2.927454167e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.51 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.322046542e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.004565279e-8
+ k1 = 4.583847700e-01 lk1 = -9.143605620e-10
+ k2 = -2.429601160e-02 lk2 = -7.952904977e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 8.611812000e+02 lvsat = 8.411710788e-2
+ ua = -6.990916173e-10 lua = -8.205135605e-16
+ ub = 2.234268964e-18 lub = 9.853555799e-26
+ uc = 5.847047920e-11 luc = -1.408521648e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.438347102e-02 lu0 = -1.017317561e-8
+ a0 = 2.202768984e+00 la0 = -7.165335746e-7
+ keta = -2.506784320e-01 lketa = 1.396330174e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.136747526e+00 lags = 6.081310502e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.189493795e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.839460957e-9
+ nfactor = {4.867876868e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.613636150e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.505300000e-05 lcit = -1.015956180e-11
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 5.672251120e-04 leta0 = -1.351628102e-10
+ etab = -5.283877540e-04 letab = 5.707641819e-11
+ dsub = 2.299473109e-01 ldsub = 3.464178733e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.573796660e-01 lpclm = -4.594153846e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 8.771783000e-03 lpdiblc2 = 5.983981900e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.026313223e-04 lalpha0 = -1.572217669e-10
+ alpha1 = 0.0
+ beta0 = 2.161396292e+01 lbeta0 = -8.499367487e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.674992940e-01 lkt1 = -2.052231484e-9
+ kt2 = -5.161637500e-02 lkt2 = 2.920874017e-8
+ at = 1.947956140e+04 lat = 5.969961705e-2
+ ute = -1.146784080e+00 lute = 5.445525125e-8
+ ua1 = 2.097537420e-09 lua1 = -1.030179567e-16
+ ub1 = -2.064788220e-18 lub1 = 3.427836151e-25
+ uc1 = 3.200892914e-11 luc1 = -8.283476799e-17 wuc1 = -6.162975822e-33
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.52 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 1e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.494846822e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.417543512e-9
+ k1 = 4.417433080e-01 lk1 = 1.590350094e-8
+ k2 = -2.483484439e-02 lk2 = -7.408360556e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -3.217170480e+04 lvsat = 1.175001425e-01 pvsat = 2.646977960e-23
+ ua = -1.159636678e-09 lua = -3.550867226e-16
+ ub = 2.271786733e-18 lub = 6.062010003e-26
+ uc = 3.204681721e-11 luc = 1.261853632e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.758494212e-02 lu0 = -3.302582306e-9
+ a0 = 2.020313377e+00 la0 = -5.321439384e-7
+ keta = -2.274052120e-01 lketa = 1.161131012e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 3.282564612e+00 lags = -1.560431697e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.073091305e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.924174767e-9
+ nfactor = {2.187167452e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.047676407e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.891464901e-03 leta0 = 2.349589317e-09 weta0 = 4.135903063e-25 peta0 = -1.972152263e-31
+ etab = -8.261744920e-04 letab = 3.580196956e-10
+ dsub = 1.364052514e-01 ldsub = 4.409514786e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 9.659588400e-02 lpclm = 1.165465516e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.219616488e-02 lpdiblc2 = -7.582698428e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -4.870901370e-05 lalpha0 = 9.678277668e-11 palpha0 = -1.232595164e-32
+ alpha1 = 0.0
+ beta0 = 1.718699924e+01 lbeta0 = 3.623952740e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.683556200e-01 lkt1 = -1.186828428e-9
+ kt2 = -9.353640400e-03 lkt2 = -1.350197941e-8
+ at = 7.564972840e+04 lat = 2.934046279e-3
+ ute = -1.055830440e+00 lute = -3.746249734e-8
+ ua1 = 2.541635640e-09 lua1 = -5.518236178e-16
+ ub1 = -2.168290200e-18 lub1 = 4.473827161e-25
+ uc1 = -8.901892120e-11 luc1 = 3.947597756e-17 wuc1 = 2.465190329e-32
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.53 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 1e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {5.092823266e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.795022070e-8
+ k1 = 3.398589120e-01 lk1 = 6.792567353e-8
+ k2 = -2.232455539e-03 lk2 = -1.894914030e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.388827547e+05 lvsat = -2.090026456e-2
+ ua = -1.480514959e-09 lua = -1.912462720e-16
+ ub = 2.596290184e-18 lub = -1.050713620e-25
+ uc = 7.232514722e-11 luc = -7.947578976e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.011729432e-02 lu0 = -4.595601340e-9
+ a0 = 4.187890080e-01 la0 = 2.855944045e-7
+ keta = 2.825571761e-02 lketa = -1.442736941e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.625831760e-01 lags = -1.205491757e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.345075300e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.963328048e-9
+ nfactor = {1.817064934e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.420670488e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.120000000e-07 lcit = 2.661247200e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 2.544581982e-03 leta0 = 8.454377845e-11
+ etab = 8.716641908e-03 letab = -4.514542358e-09 wetab = 7.237830360e-25 petab = -3.451266460e-31
+ dsub = 1.678227699e+00 ldsub = -3.463030631e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 8.100136800e-02 lpclm = 1.245091115e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.165497440e-03 lpdiblc2 = 2.644960367e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.188041066e-03 lalpha0 = 6.785257227e-10 walpha0 = 1.033975766e-25 palpha0 = 7.395570986e-32
+ alpha1 = 0.0
+ beta0 = 1.839744226e+01 lbeta0 = 3.005900535e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.701066800e-01 lkt1 = -2.927371920e-10
+ kt2 = -4.758758640e-02 lkt2 = 6.020273416e-9
+ at = 1.108500544e+05 lat = -1.503924018e-2
+ ute = -1.242925840e+00 lute = 5.806841390e-8
+ ua1 = 1.797282480e-09 lua1 = -1.717568943e-16
+ ub1 = -1.743427928e-18 lub1 = 2.304480400e-25 wub1 = 7.346839693e-40
+ uc1 = -3.144029984e-11 luc1 = 1.007633350e-17 puc1 = 1.469367939e-39
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.54 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {5.416818457e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -4.639353539e-8
+ k1 = 2.470831429e-01 lk1 = 9.210303897e-8
+ k2 = 6.961157274e-02 lk2 = -3.767169407e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 7.792280171e+04 lvsat = 2.104589919e-2
+ ua = -2.059561798e-09 lua = -4.034666577e-17
+ ub = 1.805365143e-18 lub = 1.010437038e-25
+ uc = 7.170268597e-11 luc = -7.785365576e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 5.204702371e-03 lu0 = 1.896620122e-9
+ a0 = 5.639011714e+00 la0 = -1.074795633e-6
+ keta = 1.792502891e-01 lketa = -5.377655473e-08 wketa = 2.646977960e-23 pketa = -6.310887242e-30
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.980167143e+00 lags = 7.766315574e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.759934890e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.677456896e-8
+ nfactor = {-1.037206100e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.280297364e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.361428571e-05 lcit = -3.547882857e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.918127253e-01 leta0 = 5.073405807e-08 weta0 = 3.308722450e-24 peta0 = -2.366582716e-30
+ etab = 2.237493824e-02 letab = -8.073894383e-9
+ dsub = 3.778380407e-01 ldsub = -7.421518127e-9
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.417324086e+00 lpclm = -2.237365887e-07 ppclm = -1.009741959e-28
+ pdiblc1 = -1.270942857e+00 lpdiblc1 = 4.328417086e-7
+ pdiblc2 = 6.629674286e-03 lpdiblc2 = 1.481595881e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.984745545e-03 lalpha0 = -6.695024682e-10
+ alpha1 = 0.0
+ beta0 = 3.425952577e+01 lbeta0 = -1.127758428e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.815118571e-01 lkt1 = -2.338054803e-8
+ kt2 = -3.436452571e-02 lkt2 = 2.574343801e-9
+ at = -3.756822857e+03 lat = 1.482731204e-2
+ ute = 9.931805714e-01 lute = -5.246609169e-7
+ ua1 = 4.886866343e-09 lua1 = -9.769024489e-16 pua1 = 1.880790961e-37
+ ub1 = -4.404562286e-18 lub1 = 9.239396537e-25
+ uc1 = -2.196574857e-12 luc1 = 2.455418768e-18
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.55 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {2.473098676e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 9.713763628e-09 wvth0 = -1.657128471e-07 pvth0 = 3.158486865e-14
+ k1 = 1.274291442e+00 lk1 = -1.036828628e-07 wk1 = -1.603888740e-07 pk1 = 3.057011938e-14
+ k2 = -2.987896926e-01 lk2 = 3.254558710e-08 wk2 = 6.378621990e-08 pk2 = -1.215765351e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.439540464e+05 lvsat = 8.460343950e-03 wvsat = 8.962579389e-03 pvsat = -1.708267632e-9
+ ua = 8.570943735e-10 lua = -5.962613321e-16 wua = -3.898114521e-15 pua = 7.429806277e-22
+ ub = -1.705663686e-19 lub = 4.776562499e-25 wub = 2.470200726e-24 pub = -4.708202583e-31
+ uc = -8.480010875e-11 luc = 2.204406710e-17 wuc = 2.024523317e-16 puc = -3.858741443e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 6.205559967e-02 lu0 = -8.939160902e-09 wu0 = -6.435868652e-08 pu0 = 1.226676565e-14
+ a0 = 0.0
+ keta = 1.568280748e+00 lketa = -3.185257602e-07 wketa = -1.963466532e-06 pketa = 3.742367210e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 2.643310921e-01 lags = 1.582301938e-07 wags = 1.785819056e-08 pags = -3.403771121e-15
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-3.404510258e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.812017548e-08 wvoff = 3.410435352e-07 pvoff = -6.500289780e-14
+ nfactor = {4.881776332e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.001283151e-07 wnfactor = -2.116930000e-06 pnfactor = 4.034868580e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.176666667e-05 lcit = 5.101726667e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.776689040e-01 leta0 = 4.803824572e-08 weta0 = 3.473644306e-07 peta0 = -6.620766046e-14
+ etab = -2.120138302e-01 letab = 3.660060488e-08 wetab = 1.304207654e-07 petab = -2.485819788e-14
+ dsub = 7.612804143e-01 ldsub = -8.050563453e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.828959136e+00 lpclm = -3.021942293e-07 wpclm = -1.812048274e-06 ppclm = 3.453764010e-13
+ pdiblc1 = 6.359752562e-01 lpdiblc1 = 6.938311616e-08 wpdiblc1 = 5.582865483e-07 ppdiblc1 = -1.064094161e-13
+ pdiblc2 = 7.268571389e-02 lpdiblc2 = -1.110868527e-08 wpdiblc2 = -1.903013432e-08 ppdiblc2 = 3.627143601e-15
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.287806108e-04 lalpha0 = 6.544444824e-11 walpha0 = 1.658000174e-09 palpha0 = -3.160148331e-16
+ alpha1 = 0.0
+ beta0 = 2.253272867e+01 lbeta0 = 1.107369100e-06 wbeta0 = 1.202441081e-05 pbeta0 = -2.291852700e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = 4.280353070e-01 lkt1 = -1.395602375e-07 wkt1 = -6.994830016e-07 pkt1 = 1.333214601e-13
+ kt2 = -4.304151645e-02 lkt2 = 4.228178236e-09 wkt2 = -4.157721604e-08 pkt2 = 7.924617378e-15
+ at = -9.260127561e+04 lat = 3.176106473e-02 wat = 1.484127250e-01 pat = -2.828746538e-8
+ ute = -2.207728711e+00 lute = 8.543239238e-08 wute = -1.015684588e-07 pute = 1.935894825e-14
+ ua1 = -4.255684850e-09 lua1 = 7.656678084e-16 wua1 = 2.946378216e-15 pua1 = -5.615796879e-22
+ ub1 = 6.546191676e-18 lub1 = -1.163274051e-24 wub1 = -5.070777404e-24 pub1 = 9.664901731e-31
+ uc1 = 4.677318984e-10 luc1 = -8.711294824e-17 wuc1 = -2.913117336e-16 puc1 = 5.552401642e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.56 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.4215457+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.53326
+ k2 = -0.057558508
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200550.0
+ ua = -9.7883322e-10
+ ub = 2.1342701e-18
+ uc = 2.2350587e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0291842
+ a0 = 1.9159663
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.576146
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.8262398+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0075691
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.1734937e-5
+ alpha1 = 0.0
+ beta0 = 17.793363
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25763
+ kt2 = -0.036364
+ at = 58230.0
+ ute = -1.1808
+ ua1 = 1.9636e-9
+ ub1 = -1.466e-18
+ uc1 = 6.3418e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.57 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.4215457+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.53326
+ k2 = -0.057558508
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200550.0
+ ua = -9.7883322e-10
+ ub = 2.1342701e-18
+ uc = 2.2350587e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0291842
+ a0 = 1.9159663
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.576146
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.8262398+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0075691
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.1734937e-5
+ alpha1 = 0.0
+ beta0 = 17.793363
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25763
+ kt2 = -0.036364
+ at = 58230.0
+ ute = -1.1808
+ ua1 = 1.9636e-9
+ ub1 = -1.466e-18
+ uc1 = 6.3418e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.58 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.058074269e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.311991805e-8
+ k1 = 6.089892490e-01 lk1 = -3.037197260e-7
+ k2 = -8.702084314e-02 lk2 = 1.181616413e-7
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.592386156e+05 lvsat = -6.364365617e-01 pvsat = 4.235164736e-22
+ ua = -8.498006729e-10 lua = -5.174979333e-16
+ ub = 1.984473463e-18 lub = 6.007743906e-25
+ uc = -6.918132389e-12 luc = 1.173851260e-16 puc = 4.701977403e-38
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.904396065e-02 lu0 = 5.624439371e-10
+ a0 = 1.985910349e+00 la0 = -2.805176033e-7
+ keta = 1.821905190e-01 lketa = -7.306932955e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.914922392e-01 lags = 3.479749922e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.033923399e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.743952297e-8
+ nfactor = {2.365972934e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.164653709e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.599213500e-01 leta0 = -3.205325663e-7
+ etab = -1.398683500e-01 letab = 2.802140045e-7
+ dsub = 7.185930317e-01 ldsub = -6.360532128e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.652869910e-01 lpclm = 1.392199939e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 3.368051830e-03 lpdiblc2 = 1.684872379e-8
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -4.140331570e-05 lalpha0 = 3.334342763e-10
+ alpha1 = 0.0
+ beta0 = 1.437748228e+01 lbeta0 = 1.369973122e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.466822830e-01 lkt1 = -4.390691380e-8
+ kt2 = -3.563515750e-02 lkt2 = -2.923095731e-9
+ at = 6.733600740e+04 lat = -3.652055328e-2
+ ute = -1.242223830e+00 lute = 2.463464126e-7
+ ua1 = 1.880461690e-09 lua1 = 3.334345061e-16
+ ub1 = -1.035430010e-18 lub1 = -1.726844002e-24
+ uc1 = 1.364109229e-10 luc1 = -2.927454167e-16 puc1 = -1.880790961e-37
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.59 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.322046542e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.004565279e-8
+ k1 = 4.583847700e-01 lk1 = -9.143605620e-10
+ k2 = -2.429601160e-02 lk2 = -7.952904977e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 8.611812000e+02 lvsat = 8.411710788e-2
+ ua = -6.990916173e-10 lua = -8.205135605e-16
+ ub = 2.234268964e-18 lub = 9.853555799e-26
+ uc = 5.847047920e-11 luc = -1.408521648e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.438347102e-02 lu0 = -1.017317561e-8
+ a0 = 2.202768984e+00 la0 = -7.165335746e-7
+ keta = -2.506784320e-01 lketa = 1.396330174e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.136747526e+00 lags = 6.081310502e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.189493795e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.839460957e-9
+ nfactor = {4.867876868e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.613636150e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.505300000e-05 lcit = -1.015956180e-11
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 5.672251120e-04 leta0 = -1.351628102e-10
+ etab = -5.283877540e-04 letab = 5.707641819e-11
+ dsub = 2.299473109e-01 ldsub = 3.464178733e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.573796660e-01 lpclm = -4.594153846e-08 wpclm = 2.117582368e-22
+ pdiblc1 = 0.39
+ pdiblc2 = 8.771783000e-03 lpdiblc2 = 5.983981900e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.026313223e-04 lalpha0 = -1.572217669e-10
+ alpha1 = 0.0
+ beta0 = 2.161396292e+01 lbeta0 = -8.499367487e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.674992940e-01 lkt1 = -2.052231484e-9
+ kt2 = -5.161637500e-02 lkt2 = 2.920874017e-8
+ at = 1.947956140e+04 lat = 5.969961705e-2
+ ute = -1.146784080e+00 lute = 5.445525125e-8
+ ua1 = 2.097537420e-09 lua1 = -1.030179567e-16
+ ub1 = -2.064788220e-18 lub1 = 3.427836151e-25
+ uc1 = 3.200892914e-11 luc1 = -8.283476799e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.60 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.494846822e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.417543512e-9
+ k1 = 4.417433080e-01 lk1 = 1.590350094e-8
+ k2 = -2.483484439e-02 lk2 = -7.408360556e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -3.217170480e+04 lvsat = 1.175001425e-1
+ ua = -1.159636678e-09 lua = -3.550867226e-16
+ ub = 2.271786733e-18 lub = 6.062010003e-26
+ uc = 3.204681721e-11 luc = 1.261853632e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.758494212e-02 lu0 = -3.302582306e-9
+ a0 = 2.020313377e+00 la0 = -5.321439384e-7
+ keta = -2.274052120e-01 lketa = 1.161131012e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 3.282564612e+00 lags = -1.560431697e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.073091305e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.924174767e-9
+ nfactor = {2.187167452e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.047676407e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.891464901e-03 leta0 = 2.349589317e-09 weta0 = -4.135903063e-25 peta0 = -3.944304526e-31
+ etab = -8.261744920e-04 letab = 3.580196956e-10
+ dsub = 1.364052514e-01 ldsub = 4.409514786e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 9.659588400e-02 lpclm = 1.165465516e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.219616488e-02 lpdiblc2 = -7.582698428e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -4.870901370e-05 lalpha0 = 9.678277668e-11 palpha0 = 2.465190329e-32
+ alpha1 = 0.0
+ beta0 = 1.718699924e+01 lbeta0 = 3.623952740e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.683556200e-01 lkt1 = -1.186828428e-9
+ kt2 = -9.353640400e-03 lkt2 = -1.350197941e-8
+ at = 7.564972840e+04 lat = 2.934046279e-3
+ ute = -1.055830440e+00 lute = -3.746249734e-8
+ ua1 = 2.541635640e-09 lua1 = -5.518236178e-16
+ ub1 = -2.168290200e-18 lub1 = 4.473827161e-25
+ uc1 = -8.901892120e-11 luc1 = 3.947597756e-17 wuc1 = 4.930380658e-32
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.61 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {5.092823266e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.795022070e-08 wvth0 = 4.235164736e-22
+ k1 = 3.398589120e-01 lk1 = 6.792567353e-8
+ k2 = -2.232455539e-03 lk2 = -1.894914030e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.388827547e+05 lvsat = -2.090026456e-2
+ ua = -1.480514959e-09 lua = -1.912462720e-16
+ ub = 2.596290184e-18 lub = -1.050713620e-25
+ uc = 7.232514722e-11 luc = -7.947578976e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.011729432e-02 lu0 = -4.595601340e-9
+ a0 = 4.187890080e-01 la0 = 2.855944045e-7
+ keta = 2.825571761e-02 lketa = -1.442736941e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.625831760e-01 lags = -1.205491757e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.345075300e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.963328048e-9
+ nfactor = {1.817064934e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.420670488e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.120000000e-07 lcit = 2.661247200e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 2.544581982e-03 leta0 = 8.454377845e-11
+ etab = 8.716641908e-03 letab = -4.514542358e-09 wetab = 6.203854594e-25 petab = -1.380506584e-30
+ dsub = 1.678227699e+00 ldsub = -3.463030631e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 8.100136800e-02 lpclm = 1.245091115e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.165497440e-03 lpdiblc2 = 2.644960367e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.188041066e-03 lalpha0 = 6.785257227e-10 palpha0 = 1.479114197e-31
+ alpha1 = 0.0
+ beta0 = 1.839744226e+01 lbeta0 = 3.005900535e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.701066800e-01 lkt1 = -2.927371920e-10
+ kt2 = -4.758758640e-02 lkt2 = 6.020273416e-9
+ at = 1.108500544e+05 lat = -1.503924018e-2
+ ute = -1.242925840e+00 lute = 5.806841390e-8
+ ua1 = 1.797282480e-09 lua1 = -1.717568943e-16
+ ub1 = -1.743427928e-18 lub1 = 2.304480400e-25
+ uc1 = -3.144029984e-11 luc1 = 1.007633350e-17 wuc1 = -1.232595164e-32
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.62 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {5.416818457e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -4.639353539e-8
+ k1 = 2.470831429e-01 lk1 = 9.210303897e-8
+ k2 = 6.961157274e-02 lk2 = -3.767169407e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 7.792280171e+04 lvsat = 2.104589919e-2
+ ua = -2.059561798e-09 lua = -4.034666577e-17
+ ub = 1.805365143e-18 lub = 1.010437038e-25
+ uc = 7.170268597e-11 luc = -7.785365576e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 5.204702371e-03 lu0 = 1.896620122e-9
+ a0 = 5.639011714e+00 la0 = -1.074795633e-6
+ keta = 1.792502891e-01 lketa = -5.377655473e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.980167143e+00 lags = 7.766315574e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.759934890e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.677456896e-8
+ nfactor = {-1.037206100e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.280297364e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.361428571e-05 lcit = -3.547882857e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.918127253e-01 leta0 = 5.073405807e-08 weta0 = -1.323488980e-23 peta0 = 7.888609052e-30
+ etab = 2.237493824e-02 letab = -8.073894383e-09 petab = 3.155443621e-30
+ dsub = 3.778380407e-01 ldsub = -7.421518127e-9
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.417324086e+00 lpclm = -2.237365887e-7
+ pdiblc1 = -1.270942857e+00 lpdiblc1 = 4.328417086e-7
+ pdiblc2 = 6.629674286e-03 lpdiblc2 = 1.481595881e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.984745545e-03 lalpha0 = -6.695024682e-10
+ alpha1 = 0.0
+ beta0 = 3.425952577e+01 lbeta0 = -1.127758428e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.815118571e-01 lkt1 = -2.338054803e-8
+ kt2 = -3.436452571e-02 lkt2 = 2.574343801e-9
+ at = -3.756822857e+03 lat = 1.482731204e-2
+ ute = 9.931805714e-01 lute = -5.246609169e-7
+ ua1 = 4.886866343e-09 lua1 = -9.769024489e-16 pua1 = -3.761581923e-37
+ ub1 = -4.404562286e-18 lub1 = 9.239396537e-25 pub1 = -3.503246161e-46
+ uc1 = -2.196574857e-12 luc1 = 2.455418768e-18
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.63 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.306389030e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.389307993e-07 wvth0 = 4.333565841e-07 pvth0 = -8.259776493e-14
+ k1 = 2.436557022e+00 lk1 = -3.252106824e-07 wk1 = -1.187424854e-06 pk1 = 2.263231772e-13
+ k2 = -2.287639682e-01 lk2 = 1.919868402e-08 wk2 = 1.907988488e-09 pk2 = -3.636626057e-16
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -1.269818083e+05 lvsat = 6.010071786e-02 wvsat = 2.483750474e-01 pvsat = -4.734028403e-8
+ ua = -1.087373226e-08 lua = 1.639634225e-15 wua = 6.467830437e-15 pua = -1.232768481e-21
+ ub = 3.109054962e-18 lub = -1.474395758e-25 wub = -4.278366632e-25 pub = 8.154566800e-32
+ uc = 2.809811888e-11 luc = 5.256649126e-19 wuc = 1.026898129e-16 puc = -1.957267834e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = -1.777391381e-01 lu0 = 3.676571611e-08 wu0 = 1.475359335e-07 pu0 = -2.812034892e-14
+ a0 = 0.0
+ keta = -3.264023960e+00 lketa = 6.025115171e-07 wketa = 2.306599523e-06 pketa = -4.396378690e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 2.191679348e-01 lags = 1.668382916e-07 wags = 5.776661452e-08 pags = -1.101031673e-14
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {7.795543868e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.653528562e-07 wvoff = -6.486492477e-07 pvoff = 1.236325466e-13
+ nfactor = {1.350922436e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.944519909e-06 wnfactor = -9.740574448e-06 pnfactor = 1.856553490e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.176666667e-05 lcit = 5.101726667e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -2.408013377e-01 leta0 = 6.007128758e-08 weta0 = 4.031514056e-07 peta0 = -7.684065790e-14
+ etab = 1.682800638e-01 letab = -3.588341132e-08 wetab = -2.056259341e-07 petab = 3.919230303e-14
+ dsub = 7.622193604e-01 ldsub = -8.068459766e-08 wdsub = -8.296997449e-10 pdsub = 1.581407714e-16
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.303974976e-01 lpclm = 9.031914504e-08 wpclm = 7.702215270e-09 ppclm = -1.468042230e-15
+ pdiblc1 = 2.478850522e+00 lpdiblc1 = -2.818689094e-07 wpdiblc1 = -1.070170180e-06 ppdiblc1 = 2.039744363e-13
+ pdiblc2 = 3.226476839e-01 lpdiblc2 = -5.875143675e-08 wpdiblc2 = -2.399090291e-07 ppdiblc2 = 4.572666095e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.308769144e-03 lalpha0 = 5.300414315e-10 walpha0 = 3.811941014e-09 palpha0 = -7.265559573e-16
+ alpha1 = 0.0
+ beta0 = -1.160575948e+02 lbeta0 = 2.752268474e-05 wbeta0 = 1.344897501e-04 pbeta0 = -2.563374637e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -9.494818413e-01 lkt1 = 1.229945309e-07 wkt1 = 5.177600265e-07 pkt1 = -9.868506104e-14
+ kt2 = -3.701330302e-01 lkt2 = 6.657182076e-08 wkt2 = 2.474572001e-07 pkt2 = -4.716534234e-14
+ at = 1.642598353e+05 lat = -1.719666302e-02 wat = -7.856259575e-02 pat = 1.497403075e-8
+ ute = -4.010255634e+00 lute = 4.289940238e-07 wute = 1.491234456e-06 pute = -2.842292874e-13
+ ua1 = -3.736743319e-09 lua1 = 6.667575527e-16 wua1 = 2.487815532e-15 pua1 = -4.741776404e-22
+ ub1 = 1.637036637e-19 lub1 = 5.322816369e-26 wub1 = 5.691081282e-25 pub1 = -1.084720092e-31
+ uc1 = 9.158292378e-10 luc1 = -1.725203011e-16 wuc1 = -6.872729475e-16 puc1 = 1.309942238e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.64 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.4215457+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.53326
+ k2 = -0.057558508
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200550.0
+ ua = -9.7883322e-10
+ ub = 2.1342701e-18
+ uc = 2.2350587e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0291842
+ a0 = 1.9159663
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.576146
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.8262398+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0075691
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.1734937e-5
+ alpha1 = 0.0
+ beta0 = 17.793363
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25763
+ kt2 = -0.036364
+ at = 58230.0
+ ute = -1.1808
+ ua1 = 1.9636e-9
+ ub1 = -1.466e-18
+ uc1 = 6.3418e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.65 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.4215457+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.53326
+ k2 = -0.057558508
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200550.0
+ ua = -9.7883322e-10
+ ub = 2.1342701e-18
+ uc = 2.2350587e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0291842
+ a0 = 1.9159663
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.576146
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.8262398+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0075691
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.1734937e-5
+ alpha1 = 0.0
+ beta0 = 17.793363
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25763
+ kt2 = -0.036364
+ at = 58230.0
+ ute = -1.1808
+ ua1 = 1.9636e-9
+ ub1 = -1.466e-18
+ uc1 = 6.3418e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.66 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.058074269e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.311991805e-8
+ k1 = 6.089892490e-01 lk1 = -3.037197260e-7
+ k2 = -8.702084314e-02 lk2 = 1.181616413e-7
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.592386156e+05 lvsat = -6.364365617e-1
+ ua = -8.498006729e-10 lua = -5.174979333e-16
+ ub = 1.984473463e-18 lub = 6.007743906e-25
+ uc = -6.918132389e-12 luc = 1.173851260e-16
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.904396065e-02 lu0 = 5.624439371e-10
+ a0 = 1.985910349e+00 la0 = -2.805176033e-7
+ keta = 1.821905190e-01 lketa = -7.306932955e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.914922392e-01 lags = 3.479749922e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.033923399e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.743952297e-8
+ nfactor = {2.365972934e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.164653709e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.599213500e-01 leta0 = -3.205325663e-7
+ etab = -1.398683500e-01 letab = 2.802140045e-7
+ dsub = 7.185930317e-01 ldsub = -6.360532128e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.652869910e-01 lpclm = 1.392199939e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 3.368051830e-03 lpdiblc2 = 1.684872379e-8
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -4.140331570e-05 lalpha0 = 3.334342763e-10 palpha0 = -4.930380658e-32
+ alpha1 = 0.0
+ beta0 = 1.437748228e+01 lbeta0 = 1.369973122e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.466822830e-01 lkt1 = -4.390691380e-8
+ kt2 = -3.563515750e-02 lkt2 = -2.923095731e-9
+ at = 6.733600740e+04 lat = -3.652055328e-2
+ ute = -1.242223830e+00 lute = 2.463464126e-7
+ ua1 = 1.880461690e-09 lua1 = 3.334345061e-16
+ ub1 = -1.035430010e-18 lub1 = -1.726844002e-24
+ uc1 = 1.364109229e-10 luc1 = -2.927454167e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.67 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.322046542e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.004565279e-8
+ k1 = 4.583847700e-01 lk1 = -9.143605620e-10
+ k2 = -2.429601160e-02 lk2 = -7.952904977e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 8.611812000e+02 lvsat = 8.411710788e-2
+ ua = -6.990916173e-10 lua = -8.205135605e-16
+ ub = 2.234268964e-18 lub = 9.853555799e-26
+ uc = 5.847047920e-11 luc = -1.408521648e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.438347102e-02 lu0 = -1.017317561e-08 wu0 = 1.323488980e-23
+ a0 = 2.202768984e+00 la0 = -7.165335746e-7
+ keta = -2.506784320e-01 lketa = 1.396330174e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.136747526e+00 lags = 6.081310502e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.189493795e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.839460957e-9
+ nfactor = {4.867876868e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.613636150e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.505300000e-05 lcit = -1.015956180e-11
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 5.672251120e-04 leta0 = -1.351628102e-10
+ etab = -5.283877540e-04 letab = 5.707641819e-11
+ dsub = 2.299473109e-01 ldsub = 3.464178733e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.573796660e-01 lpclm = -4.594153846e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 8.771783000e-03 lpdiblc2 = 5.983981900e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.026313223e-04 lalpha0 = -1.572217669e-10
+ alpha1 = 0.0
+ beta0 = 2.161396292e+01 lbeta0 = -8.499367487e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.674992940e-01 lkt1 = -2.052231484e-9
+ kt2 = -5.161637500e-02 lkt2 = 2.920874017e-8
+ at = 1.947956140e+04 lat = 5.969961705e-2
+ ute = -1.146784080e+00 lute = 5.445525125e-8
+ ua1 = 2.097537420e-09 lua1 = -1.030179567e-16
+ ub1 = -2.064788220e-18 lub1 = 3.427836151e-25
+ uc1 = 3.200892914e-11 luc1 = -8.283476799e-17 puc1 = 5.877471754e-39
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.68 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.494846822e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.417543512e-9
+ k1 = 4.417433080e-01 lk1 = 1.590350094e-8
+ k2 = -2.483484439e-02 lk2 = -7.408360556e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -3.217170480e+04 lvsat = 1.175001425e-1
+ ua = -1.159636678e-09 lua = -3.550867226e-16
+ ub = 2.271786733e-18 lub = 6.062010003e-26
+ uc = 3.204681721e-11 luc = 1.261853632e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.758494212e-02 lu0 = -3.302582306e-9
+ a0 = 2.020313377e+00 la0 = -5.321439384e-7
+ keta = -2.274052120e-01 lketa = 1.161131012e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 3.282564612e+00 lags = -1.560431697e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.073091305e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.924174767e-9
+ nfactor = {2.187167452e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.047676407e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.891464901e-03 leta0 = 2.349589317e-09 weta0 = 2.067951531e-25 peta0 = -2.958228395e-31
+ etab = -8.261744920e-04 letab = 3.580196956e-10
+ dsub = 1.364052514e-01 ldsub = 4.409514786e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 9.659588400e-02 lpclm = 1.165465516e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.219616488e-02 lpdiblc2 = -7.582698428e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -4.870901370e-05 lalpha0 = 9.678277668e-11 palpha0 = -1.232595164e-32
+ alpha1 = 0.0
+ beta0 = 1.718699924e+01 lbeta0 = 3.623952740e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.683556200e-01 lkt1 = -1.186828428e-9
+ kt2 = -9.353640400e-03 lkt2 = -1.350197941e-8
+ at = 7.564972840e+04 lat = 2.934046279e-3
+ ute = -1.055830440e+00 lute = -3.746249734e-8
+ ua1 = 2.541635640e-09 lua1 = -5.518236178e-16
+ ub1 = -2.168290200e-18 lub1 = 4.473827161e-25
+ uc1 = -8.901892120e-11 luc1 = 3.947597756e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.69 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {5.092823266e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.795022070e-8
+ k1 = 3.398589120e-01 lk1 = 6.792567353e-8
+ k2 = -2.232455539e-03 lk2 = -1.894914030e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.388827547e+05 lvsat = -2.090026456e-2
+ ua = -1.480514959e-09 lua = -1.912462720e-16
+ ub = 2.596290184e-18 lub = -1.050713620e-25
+ uc = 7.232514722e-11 luc = -7.947578976e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.011729432e-02 lu0 = -4.595601340e-9
+ a0 = 4.187890080e-01 la0 = 2.855944045e-7
+ keta = 2.825571761e-02 lketa = -1.442736941e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.625831760e-01 lags = -1.205491757e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.345075300e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.963328048e-9
+ nfactor = {1.817064934e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.420670488e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.120000000e-07 lcit = 2.661247200e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 2.544581982e-03 leta0 = 8.454377845e-11
+ etab = 8.716641908e-03 letab = -4.514542358e-09 wetab = 6.203854594e-25 petab = -5.176899691e-31
+ dsub = 1.678227699e+00 ldsub = -3.463030631e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 8.100136800e-02 lpclm = 1.245091115e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.165497440e-03 lpdiblc2 = 2.644960367e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.188041066e-03 lalpha0 = 6.785257227e-10 palpha0 = 7.395570986e-32
+ alpha1 = 0.0
+ beta0 = 1.839744226e+01 lbeta0 = 3.005900535e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.701066800e-01 lkt1 = -2.927371920e-10
+ kt2 = -4.758758640e-02 lkt2 = 6.020273416e-9
+ at = 1.108500544e+05 lat = -1.503924018e-2
+ ute = -1.242925840e+00 lute = 5.806841390e-8
+ ua1 = 1.797282480e-09 lua1 = -1.717568943e-16
+ ub1 = -1.743427928e-18 lub1 = 2.304480400e-25
+ uc1 = -3.144029984e-11 luc1 = 1.007633350e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.70 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {5.416818457e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -4.639353539e-8
+ k1 = 2.470831429e-01 lk1 = 9.210303897e-8
+ k2 = 6.961157274e-02 lk2 = -3.767169407e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 7.792280171e+04 lvsat = 2.104589919e-2
+ ua = -2.059561798e-09 lua = -4.034666577e-17
+ ub = 1.805365143e-18 lub = 1.010437038e-25
+ uc = 7.170268597e-11 luc = -7.785365576e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 5.204702371e-03 lu0 = 1.896620122e-9
+ a0 = 5.639011714e+00 la0 = -1.074795633e-6
+ keta = 1.792502891e-01 lketa = -5.377655473e-08 pketa = -6.310887242e-30
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.980167143e+00 lags = 7.766315574e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.759934890e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.677456896e-8
+ nfactor = {-1.037206100e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.280297364e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.361428571e-05 lcit = -3.547882857e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.918127253e-01 leta0 = 5.073405807e-08 weta0 = -9.926167351e-24 peta0 = 1.577721810e-30
+ etab = 2.237493824e-02 letab = -8.073894383e-09 petab = 1.577721810e-30
+ dsub = 3.778380407e-01 ldsub = -7.421518127e-9
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.417324086e+00 lpclm = -2.237365887e-7
+ pdiblc1 = -1.270942857e+00 lpdiblc1 = 4.328417086e-7
+ pdiblc2 = 6.629674286e-03 lpdiblc2 = 1.481595881e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.984745545e-03 lalpha0 = -6.695024682e-10 walpha0 = -1.654361225e-24
+ alpha1 = 0.0
+ beta0 = 3.425952577e+01 lbeta0 = -1.127758428e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.815118571e-01 lkt1 = -2.338054803e-8
+ kt2 = -3.436452571e-02 lkt2 = 2.574343801e-9
+ at = -3.756822857e+03 lat = 1.482731204e-2
+ ute = 9.931805714e-01 lute = -5.246609169e-7
+ ua1 = 4.886866343e-09 lua1 = -9.769024489e-16
+ ub1 = -4.404562286e-18 lub1 = 9.239396537e-25 wub1 = 7.346839693e-40 pub1 = -1.751623080e-46
+ uc1 = -2.196574857e-12 luc1 = 2.455418768e-18
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.71 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {1.627290146e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 2.583487421e-08 wvth0 = 3.965890530e-09 pvth0 = -7.558987350e-16
+ k1 = 7.956742000e-01 lk1 = -1.245841652e-8
+ k2 = -2.177876132e-01 lk2 = 1.710659076e-08 wk2 = -6.035050807e-09 pk2 = 1.150280684e-15
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.138888240e+05 lvsat = -4.869224657e-03 wvsat = 1.704014345e-03 pvsat = -3.247851342e-10
+ ua = -1.962922755e-09 lua = -5.876606748e-17 wua = 1.952313579e-17 pua = -3.721109681e-24
+ ub = 1.063189351e-19 lub = 4.248819110e-25 wub = 1.745093263e-24 pub = -3.326147759e-31
+ uc = 1.700034777e-10 luc = -2.652149647e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 1.685249332e-02 lu0 = -3.234488330e-10 wu0 = 6.719699428e-09 pu0 = -1.280774711e-15
+ a0 = 0.0
+ keta = 5.508284089e-01 lketa = -1.245993444e-07 wketa = -4.540183936e-07 pketa = 8.653590583e-14
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 2.989946667e-01 lags = 1.516233165e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.168059176e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.493417848e-09 wvoff = 1.886587311e-12 pvoff = -3.595835415e-19
+ nfactor = {7.137654675e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.942945556e-07 wnfactor = -4.811406220e-07 pnfactor = 9.170540255e-14
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.176666667e-05 lcit = 5.101726667e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 3.163069406e-01 leta0 = -4.611355026e-08 weta0 = -1.058791184e-22
+ etab = -1.158710231e-01 letab = 1.827578585e-8
+ dsub = 7.610728120e-01 ldsub = -8.046606554e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -4.493419920e-01 lpclm = 1.320499657e-07 wpclm = 1.661413987e-07 ppclm = -3.166655059e-14
+ pdiblc1 = 1.0
+ pdiblc2 = -1.873215126e-02 lpdiblc2 = 6.315559830e-09 wpdiblc2 = 7.130488600e-09 ppdiblc2 = -1.359071127e-15
+ pdiblcb = 0.0
+ drout = -3.079223206e+01 ldrout = 6.535070191e-06 wdrout = 2.481166602e-05 pdrout = -4.729103544e-12
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.923300322e-03 lalpha0 = -4.671910087e-10 walpha0 = 2.575394538e-11 palpha0 = -4.908701990e-18
+ alpha1 = 0.0
+ beta0 = 6.162003200e+01 lbeta0 = -6.342670916e-06 wbeta0 = 5.913335496e-06 pbeta0 = -1.127081746e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -4.302269100e-01 lkt1 = 2.402454105e-08 wkt1 = 1.420011955e-07 pkt1 = -2.706542785e-14
+ kt2 = -2.817600667e-02 lkt2 = 1.394812071e-9
+ at = 1.193017444e+05 lat = -8.627650877e-03 wat = -4.602867321e-02 pat = 8.773065114e-9
+ ute = -1.949543333e+00 lute = 3.622225933e-8
+ ua1 = -2.988720667e-10 lua1 = 1.149929191e-17
+ ub1 = 9.501448000e-19 lub1 = -9.666751688e-26
+ uc1 = -3.390191333e-11 luc1 = 8.498456281e-18
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.72 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.4215457+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.53326
+ k2 = -0.057558508
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200550.0
+ ua = -9.7883322e-10
+ ub = 2.1342701e-18
+ uc = 2.2350587e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0291842
+ a0 = 1.9159663
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.576146
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.8262398+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0075691
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.1734937e-5
+ alpha1 = 0.0
+ beta0 = 17.793363
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25763
+ kt2 = -0.036364
+ at = 58230.0
+ ute = -1.1808
+ ua1 = 1.9636e-9
+ ub1 = -1.466e-18
+ uc1 = 6.3418e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.73 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.4215457+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.53326
+ k2 = -0.057558508
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200550.0
+ ua = -9.7883322e-10
+ ub = 2.1342701e-18
+ uc = 2.2350587e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0291842
+ a0 = 1.9159663
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.576146
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11023409+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.8262398+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0075691
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.1734937e-5
+ alpha1 = 0.0
+ beta0 = 17.793363
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25763
+ kt2 = -0.036364
+ at = 58230.0
+ ute = -1.1808
+ ua1 = 1.9636e-9
+ ub1 = -1.466e-18
+ uc1 = 6.3418e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.74 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.058074269e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.311991805e-8
+ k1 = 6.089892490e-01 lk1 = -3.037197260e-7
+ k2 = -8.702084314e-02 lk2 = 1.181616413e-7
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.592386156e+05 lvsat = -6.364365617e-1
+ ua = -8.498006729e-10 lua = -5.174979333e-16
+ ub = 1.984473463e-18 lub = 6.007743906e-25
+ uc = -6.918132389e-12 luc = 1.173851260e-16
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.904396065e-02 lu0 = 5.624439371e-10
+ a0 = 1.985910349e+00 la0 = -2.805176033e-7
+ keta = 1.821905190e-01 lketa = -7.306932955e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.914922392e-01 lags = 3.479749922e-06 pags = 8.077935669e-28
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.033923399e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.743952297e-8
+ nfactor = {2.365972934e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.164653709e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.599213500e-01 leta0 = -3.205325663e-7
+ etab = -1.398683500e-01 letab = 2.802140045e-7
+ dsub = 7.185930317e-01 ldsub = -6.360532128e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.652869910e-01 lpclm = 1.392199939e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 3.368051830e-03 lpdiblc2 = 1.684872379e-8
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -4.140331570e-05 lalpha0 = 3.334342763e-10 palpha0 = -4.930380658e-32
+ alpha1 = 0.0
+ beta0 = 1.437748228e+01 lbeta0 = 1.369973122e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.466822830e-01 lkt1 = -4.390691380e-8
+ kt2 = -3.563515750e-02 lkt2 = -2.923095730e-9
+ at = 6.733600740e+04 lat = -3.652055328e-2
+ ute = -1.242223830e+00 lute = 2.463464126e-7
+ ua1 = 1.880461690e-09 lua1 = 3.334345061e-16
+ ub1 = -1.035430010e-18 lub1 = -1.726844002e-24
+ uc1 = 1.364109229e-10 luc1 = -2.927454167e-16 puc1 = -9.403954807e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.75 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {3.219859039e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.316514723e-07 wvth0 = 5.771604863e-08 pvth0 = -1.160438874e-13
+ k1 = 5.665343143e-01 lk1 = -2.183598343e-07 wk1 = -5.663250886e-08 pk1 = 1.138653223e-13
+ k2 = -7.557525680e-02 lk2 = 9.514914542e-08 wk2 = 2.685237675e-08 pk2 = -5.398938869e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.769825020e+04 lvsat = 1.005249695e-02 wvsat = -1.928973118e-02 pvsat = 3.878393351e-8
+ ua = 8.877692621e-10 lua = -4.011056045e-15 wua = -8.309596995e-16 pua = 1.670727572e-21
+ ub = 1.373510707e-19 lub = 4.314598673e-24 wub = 1.098051055e-24 pub = -2.207741450e-30
+ uc = -3.571360389e-11 luc = 1.752813010e-16 wuc = 4.931949511e-17 puc = -9.916177687e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.660410533e-02 lu0 = 5.468017040e-09 wu0 = 4.073664843e-09 pu0 = -8.190510533e-15
+ a0 = 2.524388491e+00 la0 = -1.363181755e-06 wa0 = -1.684160548e-07 pa0 = 3.386173198e-13
+ keta = -3.358443721e-01 lketa = 3.108676565e-07 wketa = 4.459714453e-08 pketa = -8.966701879e-14
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.235109561e+00 lags = 4.103643429e-07 wags = -5.150727956e-08 pags = 1.035605363e-13
+ b0 = 2.717129478e-07 lb0 = -5.463060528e-13 wb0 = -1.422824851e-13 pb0 = 2.860731646e-19
+ b1 = 7.646430859e-08 lb1 = -1.537391389e-13 wb1 = -4.004053519e-14 pb1 = 8.050550006e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.920230222e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.507613269e-07 wvoff = 3.826501297e-08 pvoff = -7.693563508e-14
+ nfactor = {-1.879069637e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.370428885e-06 wnfactor = 1.238881187e-06 pnfactor = -2.490894515e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 3.940003833e-05 lcit = -5.911171707e-11 wcit = -1.274932662e-11 pcit = 2.563379611e-17
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.231202960e-03 leta0 = 3.480756672e-09 weta0 = 9.417468601e-10 peta0 = -1.893476237e-15
+ etab = 1.769534418e-03 letab = -4.563125901e-09 wetab = -1.203306945e-09 petab = 2.419368944e-15
+ dsub = -1.292870681e+00 ldsub = 3.408195727e-06 wdsub = 7.974236413e-07 pdsub = -1.603299973e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 4.149536981e-01 lpclm = -3.627598874e-07 wpclm = -8.251364191e-08 ppclm = 1.659019284e-13
+ pdiblc1 = 0.39
+ pdiblc2 = -6.849276795e-03 lpdiblc2 = 3.739168472e-08 wpdiblc2 = 8.179967961e-09 ppdiblc2 = -1.644664358e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.039801412e-04 lalpha0 = -5.620537021e-10 walpha0 = -1.054363090e-10 palpha0 = 2.119902429e-16
+ alpha1 = 0.0
+ beta0 = 2.710697128e+01 lbeta0 = -1.189417936e-05 wbeta0 = -2.876413827e-06 pbeta0 = 5.783317641e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.993762807e-01 lkt1 = -1.390203619e-07 wkt1 = -3.567261589e-08 pkt1 = 7.172336151e-14
+ kt2 = -9.562608149e-02 lkt2 = 1.176946560e-07 wkt2 = 2.304568280e-08 pkt2 = -4.633564985e-14
+ at = 5.107714775e+04 lat = -3.830490064e-03 wat = -1.654607609e-02 pat = 3.326754059e-8
+ ute = -9.690507002e-01 lute = -3.028954822e-07 wute = -9.307008435e-08 pute = 1.871267116e-13
+ ua1 = 2.644858842e-09 lua1 = -1.203462407e-15 wua1 = -2.866048625e-16 pua1 = 5.762477365e-22
+ ub1 = -2.896969990e-18 lub1 = 2.015968282e-24 wub1 = 4.357719840e-25 pub1 = -8.761631510e-31
+ uc1 = 4.594796200e-10 luc1 = -9.423073390e-16 wuc1 = -2.238450273e-16 puc1 = 4.500628118e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.76 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {6.699221830e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.199729314e-07 wvth0 = -1.154320973e-07 pvth0 = 5.893962886e-14
+ k1 = 2.254442194e-01 lk1 = 1.263458156e-07 wk1 = 1.132650177e-07 pk1 = -5.783311805e-14
+ k2 = 7.772364600e-02 lk2 = -5.977472575e-08 wk2 = -5.370475349e-08 pk2 = 2.742164713e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -1.058458428e+05 lvsat = 1.551181573e-01 wvsat = 3.857946236e-02 pvsat = -1.969867348e-8
+ ua = -4.333358436e-09 lua = 1.265415607e-15 wua = 1.661919399e-15 pua = -8.485760451e-22
+ ub = 6.465622519e-18 lub = -2.080752452e-24 wub = -2.196102109e-24 pub = 1.121329737e-30
+ uc = 2.204149834e-10 luc = -8.356224933e-17 wuc = -9.863899022e-17 puc = 5.036506841e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 4.314367350e-02 lu0 = -1.124687055e-08 wu0 = -8.147329685e-09 pu0 = 4.160026537e-15
+ a0 = 1.377074363e+00 la0 = -2.037060979e-07 wa0 = 3.368321097e-07 pa0 = -1.719864752e-13
+ keta = -5.707333182e-02 lketa = 2.914164323e-08 wketa = -8.919428906e-08 pketa = 4.554260399e-14
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 3.085840542e+00 lags = -1.459984387e-06 wags = 1.030145591e-07 pags = -5.259923388e-14
+ b0 = -5.434258956e-07 lb0 = 2.774732623e-13 wb0 = 2.845649702e-13 pb0 = -1.452988738e-19
+ b1 = -1.529286172e-07 lb1 = 7.808535193e-14 wb1 = 8.008107039e-14 pb1 = -4.088939454e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {3.883815482e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.254697863e-08 wvoff = -7.653002594e-08 pvoff = 3.907623125e-14
+ nfactor = {6.918882099e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.520781139e-06 wnfactor = -2.477762375e-06 pnfactor = 1.265145469e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -4.369407667e-05 lcit = 2.486319555e-11 wcit = 2.549865325e-11 pcit = -1.301961235e-17
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.705391244e-03 leta0 = 5.130345696e-10 weta0 = -1.883493720e-09 peta0 = 9.617118935e-16
+ etab = -5.422018836e-03 letab = 2.704657818e-09 wetab = 2.406613891e-09 petab = -1.228817053e-15
+ dsub = 3.182041234e+00 ldsub = -1.114150254e-06 wdsub = -1.594847283e-06 pdsub = 8.143290224e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.185521802e-01 lpclm = 2.774611532e-07 wpclm = 1.650272838e-07 ppclm = -8.426293111e-14
+ pdiblc1 = 0.39
+ pdiblc2 = 5.343828447e-02 lpdiblc2 = -2.353492469e-08 wpdiblc2 = -1.635993592e-08 ppdiblc2 = 8.353383282e-15
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -4.514066515e-04 lalpha0 = 3.024001905e-10 walpha0 = 2.108726180e-10 palpha0 = -1.076715588e-16
+ alpha1 = 0.0
+ beta0 = 6.200982523e+00 lbeta0 = 9.233412877e-06 wbeta0 = 5.752827655e-06 pbeta0 = -2.937393801e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -4.046016465e-01 lkt1 = 6.838039271e-08 wkt1 = 7.134523178e-08 pkt1 = -3.642887535e-14
+ kt2 = 7.866577258e-02 lkt2 = -5.844469168e-08 wkt2 = -4.609136561e-08 pkt2 = 2.353425128e-14
+ at = 1.245455570e+04 lat = 3.520150146e-02 wat = 3.309215218e-02 pat = -1.689685290e-8
+ ute = -1.411297200e+00 lute = 1.440388301e-07 wute = 1.861401687e-07 pute = -9.504317014e-14
+ ua1 = 1.446992797e-09 lua1 = 7.101018090e-18 wua1 = 5.732097250e-16 pua1 = -2.926808856e-22
+ ub1 = -5.039266595e-19 lub1 = -4.024413076e-25 wub1 = -8.715439680e-25 pub1 = 4.450103500e-31
+ uc1 = -9.439603029e-10 luc1 = 4.760090470e-16 wuc1 = 4.476900545e-16 puc1 = -2.285905418e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.77 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {5.092823266e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.795022070e-8
+ k1 = 3.398589120e-01 lk1 = 6.792567353e-8
+ k2 = -2.232455539e-03 lk2 = -1.894914030e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.388827547e+05 lvsat = -2.090026456e-2
+ ua = -1.480514959e-09 lua = -1.912462720e-16
+ ub = 2.596290184e-18 lub = -1.050713620e-25
+ uc = 7.232514722e-11 luc = -7.947578976e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.011729432e-02 lu0 = -4.595601340e-9
+ a0 = 4.187890080e-01 la0 = 2.855944045e-7
+ keta = 2.825571761e-02 lketa = -1.442736941e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.625831760e-01 lags = -1.205491757e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.345075300e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.963328048e-9
+ nfactor = {1.817064934e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.420670488e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.120000000e-07 lcit = 2.661247200e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 2.544581982e-03 leta0 = 8.454377845e-11
+ etab = 8.716641908e-03 letab = -4.514542358e-09 wetab = 2.067951531e-25 petab = 4.437342592e-31
+ dsub = 1.678227699e+00 ldsub = -3.463030631e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 8.100136800e-02 lpclm = 1.245091115e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.165497440e-03 lpdiblc2 = 2.644960367e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.188041066e-03 lalpha0 = 6.785257227e-10 palpha0 = 9.860761315e-32
+ alpha1 = 0.0
+ beta0 = 1.839744226e+01 lbeta0 = 3.005900535e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.701066800e-01 lkt1 = -2.927371920e-10
+ kt2 = -4.758758640e-02 lkt2 = 6.020273416e-09 wkt2 = 2.646977960e-23
+ at = 1.108500544e+05 lat = -1.503924018e-2
+ ute = -1.242925840e+00 lute = 5.806841390e-8
+ ua1 = 1.797282480e-09 lua1 = -1.717568943e-16
+ ub1 = -1.743427928e-18 lub1 = 2.304480400e-25
+ uc1 = -3.144029984e-11 luc1 = 1.007633350e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.78 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {1.377874796e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -2.643054182e-07 wvth0 = -4.378724383e-07 pvth0 = 1.141095574e-13
+ k1 = -2.655009315e-01 lk1 = 2.256824487e-07 wk1 = 2.684146505e-07 pk1 = -6.994885793e-14
+ k2 = 3.237384768e-01 lk2 = -1.038971653e-07 wk2 = -1.330735533e-07 pk2 = 3.467896800e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.154821572e+05 lvsat = -1.480206885e-02 wvsat = -7.203295651e-02 pvsat = 1.877178847e-8
+ ua = 3.991792983e-09 lua = -1.617329722e-15 wua = -3.168791931e-15 pua = 8.257871773e-22
+ ub = -5.136743648e-19 lub = 7.053853995e-25 wub = 1.214365038e-24 pub = -3.164635289e-31
+ uc = -2.469399757e-10 luc = 7.525291205e-17 wuc = 1.668572298e-16 puc = -4.348299408e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 1.064451081e-01 lu0 = -2.448662961e-08 wu0 = -5.301453847e-08 pu0 = 1.381558872e-14
+ a0 = 5.639011714e+00 la0 = -1.074795633e-6
+ keta = 1.529171739e+00 lketa = -4.055660846e-07 wketa = -7.068863673e-07 pketa = 1.842145873e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.915880940e+00 lags = 7.598785728e-07 wags = -3.366347038e-08 pags = 8.772700380e-15
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-6.259212383e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.340257404e-07 wvoff = 2.356046659e-07 pvoff = -6.139857594e-14
+ nfactor = {-9.490229151e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.030887544e-06 wnfactor = 4.426425521e-06 pnfactor = -1.153526491e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 8.921245238e-05 lcit = -2.064276509e-11 wcit = -3.435047997e-11 pcit = 8.951735081e-18
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -2.139505585e-01 leta0 = 5.650317738e-08 weta0 = 1.159247632e-08 peta0 = -3.020999329e-15
+ etab = -1.274041225e-01 letab = 3.095852884e-08 wetab = 7.843180514e-08 petab = -2.043932842e-14
+ dsub = 1.048788213e-01 ldsub = 6.371165444e-08 wdsub = 1.429350952e-07 pdsub = -3.724888581e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.305785655e+00 lpclm = -4.552696737e-07 wpclm = -4.652429008e-07 ppclm = 1.212422999e-13
+ pdiblc1 = -1.387891049e+01 lpdiblc1 = 3.718478074e-06 wpdiblc1 = 6.602162251e-06 ppdiblc1 = -1.720523483e-12
+ pdiblc2 = -2.039677038e-02 lpdiblc2 = 8.524687361e-09 wpdiblc2 = 1.415239775e-08 ppdiblc2 = -3.688114854e-15
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.409091295e-03 lalpha0 = -7.800869707e-10 walpha0 = -2.222086520e-10 palpha0 = 5.790757471e-17
+ alpha1 = 0.0
+ beta0 = 3.758882952e+01 lbeta0 = -1.995374986e-06 wbeta0 = -1.743389910e-06 pbeta0 = 4.543274106e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = 2.792496655e-01 lkt1 = -1.434550008e-07 wkt1 = -2.412777713e-07 pkt1 = 6.287698721e-14
+ kt2 = -1.537138301e-01 lkt2 = 3.367677254e-08 wkt2 = 6.249726327e-08 pkt2 = -1.628678681e-14
+ at = -6.024996399e+04 lat = 2.954942462e-02 wat = 2.958263335e-02 pat = -7.709234252e-9
+ ute = 1.226710045e+00 lute = -5.855186977e-07 wute = -1.222877087e-07 pute = 3.186817689e-14
+ ua1 = 6.937202640e-09 lua1 = -1.511220088e-15 wua1 = -1.073658602e-15 pua1 = 2.797954317e-22
+ ub1 = -7.751643142e-18 lub1 = 1.796188925e-24 wub1 = 1.752698890e-24 pub1 = -4.567533308e-31
+ uc1 = -2.179568168e-10 luc1 = 5.868253782e-17 wuc1 = 1.129828507e-16 puc1 = -2.944333089e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.79 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.644595440e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 3.117774088e-07 wvth0 = 9.503713413e-07 pvth0 = -1.504897070e-13
+ k1 = 1.991703707e+00 lk1 = -2.045407553e-07 wk1 = -6.263008512e-07 pk1 = 1.005839167e-13
+ k2 = -7.645738587e-01 lk2 = 1.035351659e-07 wk2 = 2.802895667e-07 pk2 = -4.410804268e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 9.561298815e+05 lvsat = -1.559695251e-01 wvsat = -3.869705154e-01 pvsat = 7.879888719e-8
+ ua = -1.474738778e-08 lua = 1.954358132e-15 wua = 6.714108247e-15 pua = -1.057893597e-21
+ ub = 2.238879825e-17 lub = -3.659825882e-24 wub = -9.923127033e-24 pub = 1.806342460e-30
+ uc = 1.522724601e-09 luc = -2.620451564e-16 wuc = -7.083524165e-16 puc = 1.233319645e-22
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = -1.521959802e-01 lu0 = 2.481036182e-08 wu0 = 9.524193260e-08 pu0 = -1.444209466e-14
+ a0 = 0.0
+ keta = -3.464776626e+00 lketa = 5.462804737e-07 wketa = 1.648753183e-06 pketa = -2.647703109e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.489935256e-01 lags = 1.757134998e-07 wags = 7.854809754e-08 pags = -1.261482447e-14
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {9.330548943e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.631151105e-07 wvoff = -5.497577276e-07 pvoff = 8.829149626e-14
+ nfactor = {1.228340739e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.119167582e-06 wnfactor = -6.539583617e-06 pnfactor = 9.365948509e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.748290556e-04 lcit = 2.968354632e-11 wcit = 8.015111994e-11 pcit = -1.287226986e-17
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 3.679618846e-01 leta0 = -5.440933426e-08 weta0 = -2.704911141e-08 peta0 = 4.344087293e-15
+ etab = 2.336134519e-01 letab = -3.785142083e-08 wetab = -1.830075453e-07 petab = 2.939101178e-14
+ dsub = 1.397977657e+00 ldsub = -1.827529837e-07 wdsub = -3.335152222e-07 pdsub = 5.356254468e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -8.475975063e-01 lpclm = 1.457651569e-07 wpclm = 3.746878987e-07 ppclm = -3.884851045e-14
+ pdiblc1 = 3.041859114e+01 lpdiblc1 = -4.724625738e-06 wpdiblc1 = -1.540504525e-05 ppdiblc1 = 2.474050268e-12
+ pdiblc2 = -1.053046893e-01 lpdiblc2 = 2.470813671e-08 wpdiblc2 = 5.246419814e-08 ppdiblc2 = -1.099034401e-14
+ pdiblcb = 0.0
+ drout = 7.968756014e+01 ldrout = -1.452237820e-05 wdrout = -3.304107716e-05 pdrout = 6.297629308e-12
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.926154455e-03 lalpha0 = -3.068392089e-10 walpha0 = 5.479093787e-10 palpha0 = -8.887692195e-17
+ alpha1 = 0.0
+ beta0 = 3.798295661e+01 lbeta0 = -2.070495609e-06 wbeta0 = 1.829089003e-05 pbeta0 = -3.364206345e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -8.730433307e-01 lkt1 = 7.617204424e-08 wkt1 = 3.738820141e-07 pkt1 = -5.437246790e-14
+ kt2 = 2.503057037e-01 lkt2 = -4.332935061e-08 wkt2 = -1.458269476e-07 pkt2 = 2.341980779e-14
+ at = 2.383061371e+05 lat = -2.735536826e-02 wat = -1.083453235e-01 pat = 1.857983432e-8
+ ute = -2.494445438e+00 lute = 1.237335373e-07 wute = 2.853379870e-07 pute = -4.582528071e-14
+ ua1 = -7.896873311e-09 lua1 = 1.316154788e-15 wua1 = 3.978693352e-15 pua1 = -6.831828507e-22
+ ub1 = 8.760000131e-18 lub1 = -1.350930283e-24 wub1 = -4.089630744e-24 pub1 = 6.567946975e-31
+ uc1 = 4.695386512e-10 luc1 = -7.235409838e-17 wuc1 = -2.636266516e-16 puc1 = 4.233844025e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.80 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.263006254e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = -2.061973410e-9
+ k1 = 6.583871577e-01 wk1 = -5.426139193e-8
+ k2 = -9.227296257e-02 wk2 = 1.505392322e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 4.548895758e+05 wvsat = -1.102943570e-1
+ ua = -4.970061183e-10 wua = -2.089443227e-16
+ ub = 2.678808214e-18 wub = -2.361389533e-25
+ uc = 1.571603771e-11 wuc = 2.877072299e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 4.428448092e-02 wu0 = -6.548236822e-9
+ a0 = 2.747888585e+00 wa0 = -3.607630987e-7
+ keta = 3.036500000e-01 wketa = -1.316778225e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.186027247e+00 wags = 1.197816429e-6
+ b0 = -1.303359231e-07 wb0 = 5.652017304e-14
+ b1 = -3.667858423e-08 wb1 = 1.590566805e-14
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-6.369907348e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = -2.017990991e-8
+ nfactor = {2.360202532e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = -2.315529389e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 2.667117035e-01 weta0 = -8.096753024e-8
+ etab = -2.335038462e-01 wetab = 7.090344288e-8
+ dsub = 1.260730769e+00 wdsub = -3.038718981e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 9.657213846e-02 wpclm = 4.485149216e-8
+ pdiblc1 = 0.39
+ pdiblc2 = -1.577538731e-03 wpdiblc2 = 3.966439886e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.728345973e-05 walpha0 = 4.727582774e-11
+ alpha1 = 0.0
+ beta0 = 8.198856870e+00 wbeta0 = 4.160657583e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.625117577e-01 wkt1 = 2.116974223e-9
+ kt2 = -4.713656769e-02 wkt2 = 4.671523980e-9
+ at = -4.396644615e+03 wat = 2.715804444e-2
+ ute = -1.471369692e+00 wute = 1.260055471e-7
+ ua1 = 1.626314923e-09 wua1 = 1.462636736e-16
+ ub1 = -4.604513462e-19 wub1 = -4.360561737e-25
+ uc1 = 1.231856631e-10 wuc1 = -2.591824709e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.81 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.263006254e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} wvth0 = -2.061973410e-9
+ k1 = 6.583871577e-01 wk1 = -5.426139193e-8
+ k2 = -9.227296257e-02 wk2 = 1.505392322e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 4.548895758e+05 wvsat = -1.102943570e-1
+ ua = -4.970061183e-10 wua = -2.089443227e-16
+ ub = 2.678808214e-18 wub = -2.361389533e-25
+ uc = 1.571603771e-11 wuc = 2.877072299e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 4.428448092e-02 wu0 = -6.548236822e-9
+ a0 = 2.747888585e+00 wa0 = -3.607630987e-7
+ keta = 3.036500000e-01 wketa = -1.316778225e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.186027247e+00 wags = 1.197816429e-6
+ b0 = -1.303359231e-07 wb0 = 5.652017304e-14
+ b1 = -3.667858423e-08 wb1 = 1.590566805e-14
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-6.369907348e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} wvoff = -2.017990991e-8
+ nfactor = {2.360202532e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = -2.315529389e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 2.667117035e-01 weta0 = -8.096753024e-8
+ etab = -2.335038462e-01 wetab = 7.090344288e-8
+ dsub = 1.260730769e+00 wdsub = -3.038718981e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 9.657213846e-02 wpclm = 4.485149216e-8
+ pdiblc1 = 0.39
+ pdiblc2 = -1.577538731e-03 wpdiblc2 = 3.966439886e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.728345972e-05 walpha0 = 4.727582774e-11
+ alpha1 = 0.0
+ beta0 = 8.198856870e+00 wbeta0 = 4.160657583e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.625117577e-01 wkt1 = 2.116974223e-9
+ kt2 = -4.713656769e-02 wkt2 = 4.671523980e-9
+ at = -4.396644615e+03 wat = 2.715804444e-2
+ ute = -1.471369692e+00 wute = 1.260055471e-7
+ ua1 = 1.626314923e-09 wua1 = 1.462636736e-16
+ ub1 = -4.604513462e-19 wub1 = -4.360561737e-25
+ uc1 = 1.231856631e-10 wuc1 = -2.591824709e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.82 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {3.738013783e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.105534805e-07 wvth0 = 1.387942298e-08 pvth0 = -6.393456435e-14
+ k1 = 9.110024564e-01 lk1 = -1.013138917e-06 wk1 = -1.309680274e-07 pk1 = 3.076396321e-13
+ k2 = -1.905525136e-01 lk2 = 3.941599674e-07 wk2 = 4.489650890e-08 pk2 = -1.196866741e-13
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 9.842381770e+05 lvsat = -2.123005500e+00 wvsat = -2.710310598e-01 pvsat = 6.446506201e-7
+ ua = -6.658331792e-11 lua = -1.726253683e-15 wua = -3.396422060e-16 pua = 5.241769308e-22
+ ub = 2.179121203e-18 lub = 2.004044727e-24 wub = -8.440899235e-26 pub = -6.085281813e-31
+ uc = -8.191765585e-11 luc = 3.915696914e-16 wuc = 3.252354335e-17 puc = -1.189001368e-22
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 4.381667481e-02 lu0 = 1.876183179e-09 wu0 = -6.406187497e-09 pu0 = -5.697030224e-16
+ a0 = 2.981205791e+00 la0 = -9.357419897e-07 wa0 = -4.316098686e-07 pa0 = 2.841380552e-13
+ keta = 9.113955274e-01 lketa = -2.437424212e-06 wketa = -3.162197519e-07 pketa = 7.401238621e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -5.080268189e+00 lags = 1.160764272e-05 wags = 2.076652690e-06 pags = -3.524660712e-12
+ b0 = -1.303359231e-07 wb0 = 5.652017304e-14
+ b1 = -3.667858423e-08 wb1 = 1.590566805e-14
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-4.087657400e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -9.153191642e-08 wvoff = -2.710996188e-08 pvoff = 2.779366642e-14
+ nfactor = {4.160627715e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.220785238e-06 wnfactor = -7.782520456e-07 pnfactor = 2.192591437e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 5.333108837e-01 leta0 = -1.069222672e-06 weta0 = -1.619203713e-07 peta0 = 3.246694644e-13
+ etab = -4.665685383e-01 letab = 9.347292543e-07 wetab = 1.416735367e-07 petab = -2.838305381e-13
+ dsub = 1.789760525e+00 ldsub = -2.121726737e-06 wdsub = -4.645117833e-07 pdsub = 6.442623235e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.922244887e-02 lpclm = 4.644057719e-07 wpclm = 8.001251860e-08 ppclm = -1.410168127e-13
+ pdiblc1 = 0.39
+ pdiblc2 = -1.559126595e-02 lpdiblc2 = 5.620345440e-08 wpdiblc2 = 8.221708157e-09 ppdiblc2 = -1.706617893e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.446134850e-04 lalpha0 = 1.112259799e-09 walpha0 = 1.314870899e-10 palpha0 = -3.377376880e-16
+ alpha1 = 0.0
+ beta0 = -3.195732937e+00 lbeta0 = 4.569914188e-05 wbeta0 = 7.620624778e-06 pbeta0 = -1.387654443e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.259927002e-01 lkt1 = -1.464633321e-07 wkt1 = -8.972037591e-09 pkt1 = 4.447359078e-14
+ kt2 = -4.470531731e-02 lkt2 = -9.750772796e-09 wkt2 = 3.933274800e-09 pkt2 = 2.960822160e-15
+ at = 2.597889468e+04 lat = -1.218241379e-01 wat = 1.793451193e-02 pat = 3.699189948e-8
+ ute = -1.676265414e+00 lute = 8.217547833e-07 wute = 1.882221331e-07 pute = -2.495258399e-13
+ ua1 = 1.348984707e-09 lua1 = 1.112260566e-15 wua1 = 2.304749938e-16 pua1 = -3.377379208e-22
+ ub1 = 9.758307782e-19 lub1 = -5.760353088e-24 wub1 = -8.721832408e-25 pub1 = 1.749131215e-30
+ uc1 = 3.666732095e-10 luc1 = -9.765311535e-16 wuc1 = -9.985324055e-17 puc1 = 2.965236848e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.83 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {5.381617257e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.199094340e-07 wvth0 = -3.602859651e-08 pvth0 = 3.641049964e-14
+ k1 = 3.337479079e-01 lk1 = 1.474890783e-07 wk1 = 4.431531627e-08 pk1 = -4.478505862e-14
+ k2 = 5.418406536e-02 lk2 = -9.790739830e-08 wk2 = -2.941775331e-08 pk2 = 2.972958149e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -2.367288279e+05 lvsat = 3.318707601e-01 wvsat = 9.971557125e-02 pvsat = -1.007725563e-7
+ ua = -6.624486809e-10 lua = -5.282067842e-16 wua = -1.587076885e-16 pua = 1.603899900e-22
+ ub = 4.464093734e-18 lub = -2.590121044e-24 wub = -7.782409013e-25 pub = 7.864902549e-31
+ uc = 2.014080279e-10 luc = -1.780849284e-16 wuc = -5.350830054e-17 puc = 5.407548852e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 6.701376392e-02 lu0 = -4.476388418e-08 wu0 = -1.344998360e-08 pu0 = 1.359255343e-14
+ a0 = 3.481936494e+00 la0 = -1.942511141e-06 wa0 = -5.836567466e-07 pa0 = 5.898435081e-13
+ keta = -4.735943648e-01 lketa = 3.472364651e-07 wketa = 1.043324289e-07 pketa = -1.054383526e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -3.840867191e-01 lags = 2.165500258e-06 wags = 6.506571873e-07 pags = -6.575541535e-13
+ b0 = -3.184448869e-07 lb0 = 3.782118827e-13 wb0 = 1.136394599e-13 pb0 = -1.148440382e-19
+ b1 = -8.961541325e-08 lb1 = 1.064347884e-13 wb1 = 3.197993618e-14 pb1 = -3.231892351e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-4.218182329e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.890758221e-08 wvoff = -2.671362293e-08 pvoff = 2.699678734e-14
+ nfactor = {-4.699993891e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.089553618e-06 wnfactor = 6.278378746e-07 pnfactor = -6.344929560e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 2.987362739e-03 leta0 = -2.954200816e-09 weta0 = -8.876341556e-10 peta0 = 8.970430777e-16
+ etab = -3.353448808e-03 letab = 3.388995365e-09 wetab = 1.018274730e-09 petab = -1.029068443e-15
+ dsub = 1.214009774e+00 ldsub = -9.641222777e-07 wdsub = -2.896850679e-07 pdsub = 2.927557296e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.788877482e-01 lpclm = 6.608540962e-08 wpclm = 1.985635724e-08 ppclm = -2.006683463e-14
+ pdiblc1 = 0.39
+ pdiblc2 = 1.324891407e-02 lpdiblc2 = -1.782611562e-09 wpdiblc2 = -5.356125082e-10 ppdiblc2 = 5.412900008e-16
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.300344155e-04 lalpha0 = -2.441872695e-10 walpha0 = -7.336974508e-11 palpha0 = 7.414746438e-17
+ alpha1 = 0.0
+ beta0 = 1.714064457e+01 lbeta0 = 4.810821258e-06 wbeta0 = 1.445483747e-06 pbeta0 = -1.460805875e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -3.425955310e-01 lkt1 = 8.797831968e-08 wkt1 = 2.643441200e-08 pkt1 = -2.671461677e-14
+ kt2 = -6.754671257e-02 lkt2 = 3.617413653e-08 wkt2 = 1.086906447e-08 pkt2 = -1.098427656e-14
+ at = -1.555344175e+05 lat = 2.431265275e-01 wat = 7.305102916e-02 pat = -7.382537007e-8
+ ute = -1.480946619e+00 lute = 4.290468132e-07 wute = 1.289135809e-07 pute = -1.302800648e-13
+ ua1 = 1.694184417e-09 lua1 = 4.182020280e-16 wua1 = 1.256551017e-16 pua1 = -1.269870458e-22
+ ub1 = -1.881744825e-18 lub1 = -1.491157961e-26 wub1 = -4.480408814e-27 pub1 = 4.527901147e-33
+ uc1 = -2.775289966e-10 luc1 = 3.187018019e-16 wuc1 = 9.575875931e-17 puc1 = -9.677380216e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.84 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.037349415e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.594227410e-8
+ k1 = 4.866341600e-01 lk1 = -7.017768096e-9
+ k2 = -4.611989947e-02 lk2 = 3.459788568e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -1.688132680e+04 lvsat = 1.096928755e-1
+ ua = -5.009604218e-10 lua = -6.914068188e-16
+ ub = 1.401395356e-18 lub = 5.050419372e-25
+ uc = -7.047233185e-12 luc = 3.257995846e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.435587300e-02 lu0 = -1.653819614e-9
+ a0 = 2.153811616e+00 la0 = -6.003081391e-7
+ keta = -2.627560000e-01 lketa = 1.341632136e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 3.323392852e+00 lags = -1.581278596e-6
+ b0 = 1.127829600e-07 lb0 = -5.758697938e-14
+ b1 = 3.173890360e-08 lb1 = -1.620588418e-14
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.376406321e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 7.563089958e-9
+ nfactor = {1.205144350e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.966533552e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.510600000e-05 lcit = -5.160123600e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -2.637958740e-03 leta0 = 2.730749071e-09 weta0 = -1.550963649e-25 peta0 = -1.232595164e-32
+ etab = 1.276500000e-04 letab = -1.290030900e-10
+ dsub = -4.956880000e-01 ldsub = 7.636982928e-07 pdsub = -5.048709793e-29
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.620019160e-01 lpclm = 8.315023169e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 1.571215528e-02 lpdiblc2 = -4.271963126e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.486711313e-05 lalpha0 = 5.410880632e-11
+ alpha1 = 0.0
+ beta0 = 1.946704422e+01 lbeta0 = 2.459761774e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.400790320e-01 lkt1 = -1.562485426e-8
+ kt2 = -2.762124600e-02 lkt2 = -4.174539992e-9
+ at = 8.876529520e+04 lat = -3.762762129e-3
+ ute = -9.820566400e-01 lute = -7.513139962e-8
+ ua1 = 2.768818520e-09 lua1 = -6.678231963e-16
+ ub1 = -2.513713280e-18 lub1 = 6.237557408e-25
+ uc1 = 8.841616320e-11 luc1 = -5.112237653e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.85 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {5.092823266e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.795022070e-8
+ k1 = 3.398589120e-01 lk1 = 6.792567353e-8
+ k2 = -2.232455539e-03 lk2 = -1.894914030e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.388827547e+05 lvsat = -2.090026456e-2
+ ua = -1.480514959e-09 lua = -1.912462720e-16
+ ub = 2.596290184e-18 lub = -1.050713620e-25
+ uc = 7.232514722e-11 luc = -7.947578976e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.011729432e-02 lu0 = -4.595601340e-9
+ a0 = 4.187890080e-01 la0 = 2.855944045e-7
+ keta = 2.825571761e-02 lketa = -1.442736941e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.625831760e-01 lags = -1.205491757e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.345075300e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.963328048e-9
+ nfactor = {1.817064934e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.420670488e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.120000000e-07 lcit = 2.661247200e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 2.544581982e-03 leta0 = 8.454377845e-11
+ etab = 8.716641908e-03 letab = -4.514542358e-09 wetab = -6.203854594e-25 petab = 1.602373714e-31
+ dsub = 1.678227699e+00 ldsub = -3.463030631e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 8.100136800e-02 lpclm = 1.245091115e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.165497440e-03 lpdiblc2 = 2.644960367e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.188041066e-03 lalpha0 = 6.785257227e-10 walpha0 = -5.169878828e-26 palpha0 = -2.465190329e-32
+ alpha1 = 0.0
+ beta0 = 1.839744226e+01 lbeta0 = 3.005900535e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.701066800e-01 lkt1 = -2.927371920e-10
+ kt2 = -4.758758640e-02 lkt2 = 6.020273416e-9
+ at = 1.108500544e+05 lat = -1.503924018e-2
+ ute = -1.242925840e+00 lute = 5.806841390e-8
+ ua1 = 1.797282480e-09 lua1 = -1.717568943e-16
+ ub1 = -1.743427928e-18 lub1 = 2.304480400e-25
+ uc1 = -3.144029984e-11 luc1 = 1.007633350e-17 puc1 = -7.346839693e-40
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.86 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {3.681378229e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.167963037e-9
+ k1 = 3.534651714e-01 lk1 = 6.437988233e-8
+ k2 = 1.686991157e-02 lk2 = -2.392721717e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 4.937364457e+04 lvsat = 2.848580954e-2
+ ua = -3.315463863e-09 lua = 2.869414123e-16
+ ub = 2.286660094e-18 lub = -2.438176057e-26
+ uc = 1.378339890e-10 luc = -2.501918314e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = -1.580679657e-02 lu0 = 7.372216747e-9
+ a0 = 5.639011714e+00 la0 = -1.074795633e-6
+ keta = -1.009132772e-01 lketa = 1.923407063e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.993509143e+00 lags = 7.801084826e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-8.261519446e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.559814600e-9
+ nfactor = {7.171397426e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.708472098e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.872182252e-01 leta0 = 4.953673133e-08 weta0 = -8.271806126e-24 peta0 = -2.761013168e-30
+ etab = 5.346018086e-02 letab = -1.617470861e-08 petab = 7.888609052e-31
+ dsub = 4.344881727e-01 ldsub = -2.218454253e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.232932200e+00 lpclm = -1.756840633e-7
+ pdiblc1 = 1.345722857e+00 lpdiblc1 = -2.490613766e-7
+ pdiblc2 = 1.223876000e-02 lpdiblc2 = 1.986814400e-11
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.896676555e-03 lalpha0 = -6.465516894e-10
+ alpha1 = 0.0
+ beta0 = 3.356855993e+01 lbeta0 = -9.476927294e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.771386000e-01 lkt1 = 1.539781160e-9
+ kt2 = -9.594694286e-03 lkt2 = -3.880674269e-9
+ at = 7.967800000e+03 lat = 1.177187532e-2
+ ute = 9.447137143e-01 lute = -5.120304539e-7
+ ua1 = 4.461338229e-09 lua1 = -8.660098224e-16 wua1 = -7.888609052e-31
+ ub1 = -3.709906971e-18 lub1 = 7.429124788e-25 wub1 = -3.673419846e-40
+ uc1 = 4.258244457e-11 luc1 = -9.213993695e-18 wuc1 = -3.081487911e-33
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt__model.87 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -5.3e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 5.8175e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.363696e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.363696e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {2.666245949e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.818045821e-08 wvth0 = 1.215707731e-07 pvth0 = -2.317138935e-14
+ k1 = 5.474494667e-01 lk1 = 2.740647565e-8
+ k2 = -1.908607291e-01 lk2 = 1.566624293e-08 wk2 = 3.149886801e-08 pk2 = -6.003684242e-15
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -4.527559666e+04 lvsat = 4.652595492e-02 wvsat = 4.728897020e-02 pvsat = -9.013277720e-9
+ ua = 7.879959843e-11 lua = -3.600052035e-16 wua = 2.847320897e-16 pua = -5.426993629e-23
+ ub = -4.769423026e-18 lub = 1.320507682e-24 wub = 1.854035626e-24 pub = -3.533791902e-31
+ uc = -4.060716821e-10 luc = 7.864923778e-17 wuc = 1.280700919e-16 puc = -2.441015952e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 5.740901945e-02 lu0 = -6.582717787e-09 wu0 = 4.346724492e-09 pu0 = -8.284856881e-16
+ a0 = 0.0
+ keta = -5.173987401e-01 lketa = 9.861619987e-08 wketa = 3.706227627e-07 pketa = -7.064069856e-14
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 3.301260000e-01 lags = 1.466236244e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-3.347005338e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.048765109e-08 wvoff = 4.413854116e-12 pvoff = -8.412805944e-19
+ nfactor = {-4.591715034e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.382714930e-06 wnfactor = 7.783132240e-07 pnfactor = -1.483465005e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 3.055864403e-01 leta0 = -4.439183791e-8
+ etab = -1.884032559e-01 letab = 2.992446244e-8
+ dsub = 6.288891707e-01 ldsub = -5.923737274e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.643546667e-02 lpclm = 5.618021405e-8
+ pdiblc1 = -5.105553333e+00 lpdiblc1 = 9.805518653e-07 wpdiblc1 = 2.646977960e-22 ppdiblc1 = -8.835242138e-29
+ pdiblc2 = 1.567812667e-02 lpdiblc2 = -6.356751427e-10
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.740867895e-03 lalpha0 = -8.074545589e-10 walpha0 = -6.726911048e-10 palpha0 = 1.282149246e-16
+ alpha1 = 0.0
+ beta0 = 1.723718178e+02 lbeta0 = -2.740359367e-05 wbeta0 = -3.998683961e-05 pbeta0 = 7.621491630e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.086873333e-02 lkt1 = -4.921125543e-8
+ kt2 = -8.597228000e-02 lkt2 = 1.067689357e-8
+ at = -1.419322429e+05 lat = 4.034282350e-02 wat = 5.654505002e-02 pat = -1.077748653e-8
+ ute = -1.836454000e+00 lute = 1.806011240e-8
+ ua1 = 2.642099863e-09 lua1 = -5.192629900e-16 wua1 = -5.915323654e-16 pua1 = 1.127460689e-22
+ ub1 = -6.707176000e-19 lub1 = 1.636429846e-25
+ uc1 = -1.383862920e-10 luc1 = 2.527864750e-17 wuc1 = 6.162975822e-33 puc1 = -1.469367939e-39
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.537795114e-10
+ cgso = 2.537795114e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.45065e-11
+ cgdl = 2.45065e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = -2.164e-9
+ dwc = 5.8175e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0014211795
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.79518848e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 2.10922964e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.ends sky130_fd_pr__nfet_01v8_lvt
