magic
tech sky130A
magscale 1 2
timestamp 1624884095
<< checkpaint >>
rect -1353 -1260 2209 2865
<< nwell >>
rect -85 1548 913 1568
rect -93 1266 913 1548
rect -85 800 913 1266
<< pwell >>
rect 67 671 873 728
rect -45 76 873 671
<< mvnmos >>
rect 146 102 266 702
rect 322 102 442 702
rect 498 102 618 702
rect 674 102 794 702
<< mvpmos >>
rect 134 866 234 1466
rect 290 866 390 1466
rect 446 866 546 1466
rect 602 866 702 1466
<< mvndiff >>
rect 93 624 146 702
rect 93 590 101 624
rect 135 590 146 624
rect 93 556 146 590
rect 93 522 101 556
rect 135 522 146 556
rect 93 488 146 522
rect 93 454 101 488
rect 135 454 146 488
rect 93 420 146 454
rect 93 386 101 420
rect 135 386 146 420
rect 93 352 146 386
rect 93 318 101 352
rect 135 318 146 352
rect 93 284 146 318
rect 93 250 101 284
rect 135 250 146 284
rect 93 216 146 250
rect 93 182 101 216
rect 135 182 146 216
rect 93 148 146 182
rect 93 114 101 148
rect 135 114 146 148
rect 93 102 146 114
rect 266 624 322 702
rect 266 590 277 624
rect 311 590 322 624
rect 266 556 322 590
rect 266 522 277 556
rect 311 522 322 556
rect 266 488 322 522
rect 266 454 277 488
rect 311 454 322 488
rect 266 420 322 454
rect 266 386 277 420
rect 311 386 322 420
rect 266 352 322 386
rect 266 318 277 352
rect 311 318 322 352
rect 266 284 322 318
rect 266 250 277 284
rect 311 250 322 284
rect 266 216 322 250
rect 266 182 277 216
rect 311 182 322 216
rect 266 148 322 182
rect 266 114 277 148
rect 311 114 322 148
rect 266 102 322 114
rect 442 624 498 702
rect 442 590 453 624
rect 487 590 498 624
rect 442 556 498 590
rect 442 522 453 556
rect 487 522 498 556
rect 442 488 498 522
rect 442 454 453 488
rect 487 454 498 488
rect 442 420 498 454
rect 442 386 453 420
rect 487 386 498 420
rect 442 352 498 386
rect 442 318 453 352
rect 487 318 498 352
rect 442 284 498 318
rect 442 250 453 284
rect 487 250 498 284
rect 442 216 498 250
rect 442 182 453 216
rect 487 182 498 216
rect 442 148 498 182
rect 442 114 453 148
rect 487 114 498 148
rect 442 102 498 114
rect 618 624 674 702
rect 618 590 629 624
rect 663 590 674 624
rect 618 556 674 590
rect 618 522 629 556
rect 663 522 674 556
rect 618 488 674 522
rect 618 454 629 488
rect 663 454 674 488
rect 618 420 674 454
rect 618 386 629 420
rect 663 386 674 420
rect 618 352 674 386
rect 618 318 629 352
rect 663 318 674 352
rect 618 284 674 318
rect 618 250 629 284
rect 663 250 674 284
rect 618 216 674 250
rect 618 182 629 216
rect 663 182 674 216
rect 618 148 674 182
rect 618 114 629 148
rect 663 114 674 148
rect 618 102 674 114
rect 794 624 847 702
rect 794 590 805 624
rect 839 590 847 624
rect 794 556 847 590
rect 794 522 805 556
rect 839 522 847 556
rect 794 488 847 522
rect 794 454 805 488
rect 839 454 847 488
rect 794 420 847 454
rect 794 386 805 420
rect 839 386 847 420
rect 794 352 847 386
rect 794 318 805 352
rect 839 318 847 352
rect 794 284 847 318
rect 794 250 805 284
rect 839 250 847 284
rect 794 216 847 250
rect 794 182 805 216
rect 839 182 847 216
rect 794 148 847 182
rect 794 114 805 148
rect 839 114 847 148
rect 794 102 847 114
<< mvpdiff >>
rect 81 1454 134 1466
rect 81 1420 89 1454
rect 123 1420 134 1454
rect 81 1386 134 1420
rect 81 1352 89 1386
rect 123 1352 134 1386
rect 81 1318 134 1352
rect 81 1284 89 1318
rect 123 1284 134 1318
rect 81 1250 134 1284
rect 81 1216 89 1250
rect 123 1216 134 1250
rect 81 1182 134 1216
rect 81 1148 89 1182
rect 123 1148 134 1182
rect 81 1114 134 1148
rect 81 1080 89 1114
rect 123 1080 134 1114
rect 81 1046 134 1080
rect 81 1012 89 1046
rect 123 1012 134 1046
rect 81 978 134 1012
rect 81 944 89 978
rect 123 944 134 978
rect 81 866 134 944
rect 234 1454 290 1466
rect 234 1420 245 1454
rect 279 1420 290 1454
rect 234 1386 290 1420
rect 234 1352 245 1386
rect 279 1352 290 1386
rect 234 1318 290 1352
rect 234 1284 245 1318
rect 279 1284 290 1318
rect 234 1250 290 1284
rect 234 1216 245 1250
rect 279 1216 290 1250
rect 234 1182 290 1216
rect 234 1148 245 1182
rect 279 1148 290 1182
rect 234 1114 290 1148
rect 234 1080 245 1114
rect 279 1080 290 1114
rect 234 1046 290 1080
rect 234 1012 245 1046
rect 279 1012 290 1046
rect 234 978 290 1012
rect 234 944 245 978
rect 279 944 290 978
rect 234 866 290 944
rect 390 1454 446 1466
rect 390 1420 401 1454
rect 435 1420 446 1454
rect 390 1386 446 1420
rect 390 1352 401 1386
rect 435 1352 446 1386
rect 390 1318 446 1352
rect 390 1284 401 1318
rect 435 1284 446 1318
rect 390 1250 446 1284
rect 390 1216 401 1250
rect 435 1216 446 1250
rect 390 1182 446 1216
rect 390 1148 401 1182
rect 435 1148 446 1182
rect 390 1114 446 1148
rect 390 1080 401 1114
rect 435 1080 446 1114
rect 390 1046 446 1080
rect 390 1012 401 1046
rect 435 1012 446 1046
rect 390 978 446 1012
rect 390 944 401 978
rect 435 944 446 978
rect 390 866 446 944
rect 546 1454 602 1466
rect 546 1420 557 1454
rect 591 1420 602 1454
rect 546 1386 602 1420
rect 546 1352 557 1386
rect 591 1352 602 1386
rect 546 1318 602 1352
rect 546 1284 557 1318
rect 591 1284 602 1318
rect 546 1250 602 1284
rect 546 1216 557 1250
rect 591 1216 602 1250
rect 546 1182 602 1216
rect 546 1148 557 1182
rect 591 1148 602 1182
rect 546 1114 602 1148
rect 546 1080 557 1114
rect 591 1080 602 1114
rect 546 1046 602 1080
rect 546 1012 557 1046
rect 591 1012 602 1046
rect 546 978 602 1012
rect 546 944 557 978
rect 591 944 602 978
rect 546 866 602 944
rect 702 1454 755 1466
rect 702 1420 713 1454
rect 747 1420 755 1454
rect 702 1386 755 1420
rect 702 1352 713 1386
rect 747 1352 755 1386
rect 702 1318 755 1352
rect 702 1284 713 1318
rect 747 1284 755 1318
rect 702 1250 755 1284
rect 702 1216 713 1250
rect 747 1216 755 1250
rect 702 1182 755 1216
rect 702 1148 713 1182
rect 747 1148 755 1182
rect 702 1114 755 1148
rect 702 1080 713 1114
rect 747 1080 755 1114
rect 702 1046 755 1080
rect 702 1012 713 1046
rect 747 1012 755 1046
rect 702 978 755 1012
rect 702 944 713 978
rect 747 944 755 978
rect 702 866 755 944
<< mvndiffc >>
rect 101 590 135 624
rect 101 522 135 556
rect 101 454 135 488
rect 101 386 135 420
rect 101 318 135 352
rect 101 250 135 284
rect 101 182 135 216
rect 101 114 135 148
rect 277 590 311 624
rect 277 522 311 556
rect 277 454 311 488
rect 277 386 311 420
rect 277 318 311 352
rect 277 250 311 284
rect 277 182 311 216
rect 277 114 311 148
rect 453 590 487 624
rect 453 522 487 556
rect 453 454 487 488
rect 453 386 487 420
rect 453 318 487 352
rect 453 250 487 284
rect 453 182 487 216
rect 453 114 487 148
rect 629 590 663 624
rect 629 522 663 556
rect 629 454 663 488
rect 629 386 663 420
rect 629 318 663 352
rect 629 250 663 284
rect 629 182 663 216
rect 629 114 663 148
rect 805 590 839 624
rect 805 522 839 556
rect 805 454 839 488
rect 805 386 839 420
rect 805 318 839 352
rect 805 250 839 284
rect 805 182 839 216
rect 805 114 839 148
<< mvpdiffc >>
rect 89 1420 123 1454
rect 89 1352 123 1386
rect 89 1284 123 1318
rect 89 1216 123 1250
rect 89 1148 123 1182
rect 89 1080 123 1114
rect 89 1012 123 1046
rect 89 944 123 978
rect 245 1420 279 1454
rect 245 1352 279 1386
rect 245 1284 279 1318
rect 245 1216 279 1250
rect 245 1148 279 1182
rect 245 1080 279 1114
rect 245 1012 279 1046
rect 245 944 279 978
rect 401 1420 435 1454
rect 401 1352 435 1386
rect 401 1284 435 1318
rect 401 1216 435 1250
rect 401 1148 435 1182
rect 401 1080 435 1114
rect 401 1012 435 1046
rect 401 944 435 978
rect 557 1420 591 1454
rect 557 1352 591 1386
rect 557 1284 591 1318
rect 557 1216 591 1250
rect 557 1148 591 1182
rect 557 1080 591 1114
rect 557 1012 591 1046
rect 557 944 591 978
rect 713 1420 747 1454
rect 713 1352 747 1386
rect 713 1284 747 1318
rect 713 1216 747 1250
rect 713 1148 747 1182
rect 713 1080 747 1114
rect 713 1012 747 1046
rect 713 944 747 978
<< mvpsubdiff >>
rect -19 597 19 645
rect -19 563 -17 597
rect 17 563 19 597
rect -19 529 19 563
rect -19 495 -17 529
rect 17 495 19 529
rect -19 461 19 495
rect -19 427 -17 461
rect 17 427 19 461
rect -19 393 19 427
rect -19 359 -17 393
rect 17 359 19 393
rect -19 325 19 359
rect -19 291 -17 325
rect 17 291 19 325
rect -19 257 19 291
rect -19 223 -17 257
rect 17 223 19 257
rect -19 189 19 223
rect -19 155 -17 189
rect 17 155 19 189
rect -19 102 19 155
<< mvnsubdiff >>
rect -27 1458 7 1482
rect -27 1390 7 1424
rect -27 1332 7 1356
rect 809 1413 847 1462
rect 809 1379 811 1413
rect 845 1379 847 1413
rect 809 1345 847 1379
rect 809 1311 811 1345
rect 845 1311 847 1345
rect 809 1277 847 1311
rect 809 1243 811 1277
rect 845 1243 847 1277
rect 809 1209 847 1243
rect 809 1175 811 1209
rect 845 1175 847 1209
rect 809 1134 847 1175
rect 809 1100 811 1134
rect 845 1100 847 1134
rect 809 1066 847 1100
rect 809 1032 811 1066
rect 845 1032 847 1066
rect 809 998 847 1032
rect 809 964 811 998
rect 845 964 847 998
rect 809 930 847 964
rect 809 896 811 930
rect 845 896 847 930
rect 809 866 847 896
<< mvpsubdiffcont >>
rect -17 563 17 597
rect -17 495 17 529
rect -17 427 17 461
rect -17 359 17 393
rect -17 291 17 325
rect -17 223 17 257
rect -17 155 17 189
<< mvnsubdiffcont >>
rect -27 1424 7 1458
rect -27 1356 7 1390
rect 811 1379 845 1413
rect 811 1311 845 1345
rect 811 1243 845 1277
rect 811 1175 845 1209
rect 811 1100 845 1134
rect 811 1032 845 1066
rect 811 964 845 998
rect 811 896 845 930
<< poly >>
rect 290 1548 702 1564
rect 290 1514 342 1548
rect 376 1514 410 1548
rect 444 1514 478 1548
rect 512 1514 546 1548
rect 580 1514 614 1548
rect 648 1514 702 1548
rect 290 1492 702 1514
rect 134 1466 234 1492
rect 290 1466 390 1492
rect 446 1466 546 1492
rect 602 1466 702 1492
rect 134 840 234 866
rect 290 840 390 866
rect 446 840 546 866
rect 602 840 702 866
rect 92 796 234 840
rect 92 782 442 796
rect 92 748 112 782
rect 146 748 180 782
rect 214 778 442 782
rect 214 748 317 778
rect 92 744 317 748
rect 351 744 442 778
rect 92 728 442 744
rect 146 702 266 728
rect 322 702 442 728
rect 498 785 794 840
rect 498 751 527 785
rect 561 751 595 785
rect 629 751 663 785
rect 697 751 731 785
rect 765 751 794 785
rect 498 728 794 751
rect 498 702 618 728
rect 674 702 794 728
rect 146 76 266 102
rect 322 76 442 102
rect 146 54 442 76
rect 146 20 175 54
rect 209 20 243 54
rect 277 20 311 54
rect 345 20 379 54
rect 413 20 442 54
rect 146 0 442 20
rect 498 76 618 102
rect 674 76 794 102
rect 498 54 794 76
rect 498 20 527 54
rect 561 20 595 54
rect 629 20 663 54
rect 697 20 731 54
rect 765 20 794 54
rect 498 0 794 20
<< polycont >>
rect 342 1514 376 1548
rect 410 1514 444 1548
rect 478 1514 512 1548
rect 546 1514 580 1548
rect 614 1514 648 1548
rect 112 748 146 782
rect 180 748 214 782
rect 317 744 351 778
rect 527 751 561 785
rect 595 751 629 785
rect 663 751 697 785
rect 731 751 765 785
rect 175 20 209 54
rect 243 20 277 54
rect 311 20 345 54
rect 379 20 413 54
rect 527 20 561 54
rect 595 20 629 54
rect 663 20 697 54
rect 731 20 765 54
<< locali >>
rect 292 1593 931 1605
rect 292 1559 309 1593
rect 343 1559 381 1593
rect 415 1559 453 1593
rect 487 1559 526 1593
rect 560 1559 599 1593
rect 633 1559 672 1593
rect 706 1559 745 1593
rect 779 1559 818 1593
rect 852 1559 891 1593
rect 925 1559 931 1593
rect 292 1548 931 1559
rect 292 1514 342 1548
rect 376 1514 410 1548
rect 444 1514 478 1548
rect 512 1514 546 1548
rect 580 1514 614 1548
rect 648 1514 931 1548
rect 292 1512 931 1514
rect -27 1458 48 1482
rect 7 1424 48 1458
rect -27 1390 48 1424
rect 7 1356 48 1390
rect -27 1332 48 1356
rect -23 1268 48 1332
rect -23 1234 14 1268
rect -23 1189 48 1234
rect -23 1155 14 1189
rect -23 1110 48 1155
rect -23 1076 14 1110
rect -23 1031 48 1076
rect -23 997 14 1031
rect -23 952 48 997
rect -23 918 14 952
rect 89 1454 123 1470
rect 89 1386 123 1420
rect 89 1332 123 1352
rect 245 1454 279 1470
rect 245 1386 279 1420
rect 89 1318 101 1332
rect 135 1298 173 1332
rect 245 1318 279 1352
rect 401 1454 435 1470
rect 401 1386 435 1420
rect 401 1332 435 1352
rect 557 1454 591 1470
rect 557 1386 591 1420
rect 89 1250 123 1284
rect 89 1182 123 1216
rect 89 1114 123 1148
rect 89 1046 123 1080
rect 89 978 123 1012
rect 89 928 123 944
rect 409 1318 447 1332
rect 435 1298 447 1318
rect 557 1318 591 1352
rect 713 1454 747 1470
rect 713 1386 747 1420
rect 713 1332 747 1352
rect 245 1250 279 1284
rect 245 1182 279 1216
rect 245 1114 279 1148
rect 245 1046 279 1068
rect 245 978 279 996
rect 401 1250 435 1284
rect 401 1182 435 1216
rect 401 1114 435 1148
rect 401 1046 435 1080
rect 401 978 435 1012
rect 37 782 367 796
rect 37 748 112 782
rect 146 748 180 782
rect 214 778 367 782
rect 214 748 317 778
rect 37 744 317 748
rect 351 744 367 778
rect 37 703 367 744
rect 401 717 435 944
rect 675 1298 713 1332
rect 557 1250 591 1284
rect 557 1182 591 1216
rect 557 1114 591 1148
rect 557 1046 591 1068
rect 557 978 591 996
rect 713 1250 747 1284
rect 713 1182 747 1216
rect 713 1114 747 1148
rect 713 1046 747 1080
rect 713 978 747 1012
rect 713 928 747 944
rect 811 1413 845 1454
rect 811 1345 845 1379
rect 811 1277 845 1311
rect 811 1209 845 1243
rect 811 1134 845 1175
rect 811 1066 845 1068
rect 811 1030 845 1032
rect 811 958 845 964
rect 811 874 845 896
rect 511 751 527 785
rect 561 751 595 785
rect 629 751 663 785
rect 697 751 731 785
rect 765 751 781 785
rect 401 674 663 717
rect -17 597 17 637
rect -17 529 17 542
rect -17 461 17 470
rect -17 393 17 398
rect -17 325 17 359
rect -17 257 17 291
rect -17 189 17 223
rect -17 110 17 155
rect 101 624 135 640
rect 101 556 135 590
rect 101 488 135 522
rect 101 420 135 454
rect 101 352 135 386
rect 277 624 311 640
rect 277 576 311 590
rect 277 504 311 522
rect 277 432 311 454
rect 277 352 311 386
rect 101 284 135 318
rect 169 295 207 329
rect 453 624 487 640
rect 453 556 487 590
rect 453 488 487 522
rect 453 420 487 454
rect 453 352 487 386
rect 101 216 135 250
rect 101 148 135 182
rect 101 98 135 114
rect 277 284 311 318
rect 449 318 453 329
rect 629 624 663 674
rect 629 556 663 590
rect 629 488 663 522
rect 629 420 663 454
rect 629 352 663 386
rect 449 295 487 318
rect 805 624 839 640
rect 805 556 839 590
rect 805 488 839 522
rect 805 420 839 454
rect 805 352 839 386
rect 277 216 311 250
rect 277 148 311 182
rect 277 98 311 114
rect 453 284 487 295
rect 453 216 487 250
rect 453 148 487 182
rect 453 98 487 114
rect 629 284 663 318
rect 733 295 771 329
rect 629 216 663 250
rect 629 148 663 182
rect 629 98 663 114
rect 805 284 839 318
rect 805 216 839 250
rect 805 148 839 182
rect 805 98 839 114
rect 159 20 175 54
rect 209 20 243 54
rect 277 20 311 54
rect 345 20 379 54
rect 413 20 429 54
rect 511 20 527 54
rect 561 20 595 54
rect 629 20 663 54
rect 697 20 731 54
rect 765 20 781 54
<< viali >>
rect 309 1559 343 1593
rect 381 1559 415 1593
rect 453 1559 487 1593
rect 526 1559 560 1593
rect 599 1559 633 1593
rect 672 1559 706 1593
rect 745 1559 779 1593
rect 818 1559 852 1593
rect 891 1559 925 1593
rect 14 1234 48 1268
rect 14 1155 48 1189
rect 14 1076 48 1110
rect 14 997 48 1031
rect 14 918 48 952
rect 101 1318 135 1332
rect 101 1298 123 1318
rect 123 1298 135 1318
rect 173 1298 207 1332
rect 375 1318 409 1332
rect 375 1298 401 1318
rect 401 1298 409 1318
rect 447 1298 481 1332
rect 245 1080 279 1102
rect 245 1068 279 1080
rect 245 1012 279 1030
rect 245 996 279 1012
rect 245 944 279 958
rect 245 924 279 944
rect 641 1298 675 1332
rect 713 1318 747 1332
rect 713 1298 747 1318
rect 557 1080 591 1102
rect 557 1068 591 1080
rect 557 1012 591 1030
rect 557 996 591 1012
rect 557 944 591 958
rect 557 924 591 944
rect 811 1100 845 1102
rect 811 1068 845 1100
rect 811 998 845 1030
rect 811 996 845 998
rect 811 930 845 958
rect 811 924 845 930
rect -17 563 17 576
rect -17 542 17 563
rect -17 495 17 504
rect -17 470 17 495
rect -17 427 17 432
rect -17 398 17 427
rect 277 556 311 576
rect 277 542 311 556
rect 277 488 311 504
rect 277 470 311 488
rect 277 420 311 432
rect 277 398 311 420
rect 135 295 169 329
rect 207 295 241 329
rect 415 295 449 329
rect 487 295 521 329
rect 699 295 733 329
rect 771 295 805 329
<< metal1 >>
tri 815 1599 821 1605 se
rect 821 1599 827 1605
rect 297 1593 827 1599
rect 297 1559 309 1593
rect 343 1559 381 1593
rect 415 1559 453 1593
rect 487 1559 526 1593
rect 560 1559 599 1593
rect 633 1559 672 1593
rect 706 1559 745 1593
rect 779 1559 818 1593
rect 297 1553 827 1559
rect 879 1553 891 1605
rect 943 1553 949 1605
rect 89 1332 759 1338
rect 89 1298 101 1332
rect 135 1298 173 1332
rect 207 1298 375 1332
rect 409 1298 447 1332
rect 481 1298 641 1332
rect 675 1298 713 1332
rect 747 1298 759 1332
rect 89 1292 759 1298
rect 8 1268 54 1280
rect 8 1234 14 1268
rect 48 1234 54 1268
rect 8 1189 54 1234
rect 8 1155 14 1189
rect 48 1155 54 1189
tri -26 1110 8 1144 se
rect 8 1110 54 1155
tri -28 1108 -26 1110 se
rect -26 1108 14 1110
rect -29 1076 14 1108
rect 48 1108 54 1110
tri 54 1108 90 1144 sw
rect 48 1102 857 1108
rect 48 1076 245 1102
rect -29 1068 245 1076
rect 279 1068 557 1102
rect 591 1068 811 1102
rect 845 1068 857 1102
rect -29 1031 857 1068
rect -29 997 14 1031
rect 48 1030 857 1031
rect 48 997 245 1030
rect -29 996 245 997
rect 279 996 557 1030
rect 591 996 811 1030
rect 845 996 857 1030
rect -29 958 857 996
rect -29 952 245 958
rect -29 918 14 952
rect 48 924 245 952
rect 279 924 557 958
rect 591 924 811 958
rect 845 924 857 958
rect 48 918 857 924
rect -29 906 857 918
tri 784 826 790 832 ne
rect 790 826 796 878
rect 848 826 860 878
rect 912 826 918 878
tri 918 826 924 832 nw
rect -29 576 857 582
rect -29 542 -17 576
rect 17 542 277 576
rect 311 542 857 576
rect -29 504 857 542
rect -29 470 -17 504
rect 17 470 277 504
rect 311 470 857 504
rect -29 432 857 470
rect -29 398 -17 432
rect 17 398 277 432
rect 311 398 857 432
rect -29 380 857 398
rect 129 329 811 341
rect 129 295 135 329
rect 169 295 207 329
rect 241 295 415 329
rect 449 295 487 329
rect 521 295 699 329
rect 733 295 771 329
rect 805 295 811 329
rect 129 283 811 295
<< via1 >>
rect 827 1593 879 1605
rect 827 1559 852 1593
rect 852 1559 879 1593
rect 827 1553 879 1559
rect 891 1593 943 1605
rect 891 1559 925 1593
rect 925 1559 943 1593
rect 891 1553 943 1559
rect 796 826 848 878
rect 860 826 912 878
<< metal2 >>
rect 821 1553 827 1605
rect 879 1553 891 1605
rect 943 1553 949 1605
tri 866 1524 895 1553 ne
tri 867 1019 895 1047 se
rect 895 1025 949 1553
rect 895 1019 943 1025
tri 943 1019 949 1025 nw
tri 790 878 867 955 se
rect 867 878 918 1019
tri 918 994 943 1019 nw
rect 790 826 796 878
rect 848 826 860 878
rect 912 826 918 878
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_0
timestamp 1624884095
transform 0 -1 230 -1 0 798
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180854  sky130_fd_pr__via_pol1__example_5595914180854_0
timestamp 1624884095
transform 0 1 326 1 0 1498
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808298  sky130_fd_pr__via_pol1__example_55959141808298_0
timestamp 1624884095
transform 0 -1 781 -1 0 801
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808298  sky130_fd_pr__via_pol1__example_55959141808298_1
timestamp 1624884095
transform 0 1 511 1 0 4
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808298  sky130_fd_pr__via_pol1__example_55959141808298_2
timestamp 1624884095
transform 0 1 159 1 0 4
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1624884095
transform -1 0 481 0 -1 1332
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1624884095
transform -1 0 747 0 -1 1332
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1624884095
transform -1 0 207 0 -1 1332
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_0
timestamp 1624884095
transform 1 0 -17 0 1 398
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_1
timestamp 1624884095
transform 1 0 811 0 -1 1102
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_2
timestamp 1624884095
transform 1 0 557 0 -1 1102
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_3
timestamp 1624884095
transform 1 0 245 0 -1 1102
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808128  sky130_fd_pr__via_l1m1__example_55959141808128_4
timestamp 1624884095
transform 1 0 277 0 1 398
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_0
timestamp 1624884095
transform 0 -1 805 1 0 295
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_1
timestamp 1624884095
transform 0 -1 521 1 0 295
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_2
timestamp 1624884095
transform 0 -1 241 1 0 295
box 0 0 1 1
use sky130_fd_pr__pfet_01v8__example_55959141808314  sky130_fd_pr__pfet_01v8__example_55959141808314_0
timestamp 1624884095
transform -1 0 234 0 -1 1466
box -28 0 128 267
use sky130_fd_pr__pfet_01v8__example_55959141808363  sky130_fd_pr__pfet_01v8__example_55959141808363_0
timestamp 1624884095
transform 1 0 290 0 -1 1466
box -28 0 440 267
use sky130_fd_pr__nfet_01v8__example_55959141808362  sky130_fd_pr__nfet_01v8__example_55959141808362_0
timestamp 1624884095
transform 1 0 498 0 1 102
box -28 0 324 267
use sky130_fd_pr__nfet_01v8__example_55959141808362  sky130_fd_pr__nfet_01v8__example_55959141808362_1
timestamp 1624884095
transform 1 0 146 0 1 102
box -28 0 324 267
<< labels >>
flabel locali s 96 748 130 782 8 FreeSans 300 0 0 0 PUEN_H
port 1 nsew
flabel locali s 747 751 781 785 7 FreeSans 300 0 0 0 DRVHI_H
port 2 nsew
flabel metal1 s 107 1292 147 1338 3 FreeSans 300 180 0 0 PU_H_N
port 3 nsew
flabel metal1 s -29 380 5 582 7 FreeSans 300 0 0 0 VGND_IO
port 4 nsew
flabel metal1 s -29 906 8 1108 7 FreeSans 300 0 0 0 VCC_IO
port 5 nsew
flabel metal1 s 823 380 857 582 7 FreeSans 300 180 0 0 VGND_IO
port 4 nsew
flabel metal1 s 719 1292 759 1338 3 FreeSans 300 0 0 0 PU_H_N
port 3 nsew
flabel metal1 s 820 906 857 1108 6 FreeSans 300 180 0 0 VCC_IO
port 5 nsew
flabel comment s 389 312 389 312 0 FreeSans 200 0 0 0 INT
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 11928220
string GDS_START 11919692
<< end >>
