magic
tech sky130A
magscale 1 2
timestamp 1624883981
<< checkpaint >>
rect -1250 -1349 1894 1561
<< pwell >>
rect 10 10 634 230
<< nmoslvt >>
rect 92 36 122 204
rect 178 36 208 204
rect 264 36 294 204
rect 350 36 380 204
rect 436 36 466 204
rect 522 36 552 204
<< ndiff >>
rect 36 173 92 204
rect 36 139 47 173
rect 81 139 92 173
rect 36 101 92 139
rect 36 67 47 101
rect 81 67 92 101
rect 36 36 92 67
rect 122 173 178 204
rect 122 139 133 173
rect 167 139 178 173
rect 122 101 178 139
rect 122 67 133 101
rect 167 67 178 101
rect 122 36 178 67
rect 208 173 264 204
rect 208 139 219 173
rect 253 139 264 173
rect 208 101 264 139
rect 208 67 219 101
rect 253 67 264 101
rect 208 36 264 67
rect 294 173 350 204
rect 294 139 305 173
rect 339 139 350 173
rect 294 101 350 139
rect 294 67 305 101
rect 339 67 350 101
rect 294 36 350 67
rect 380 173 436 204
rect 380 139 391 173
rect 425 139 436 173
rect 380 101 436 139
rect 380 67 391 101
rect 425 67 436 101
rect 380 36 436 67
rect 466 173 522 204
rect 466 139 477 173
rect 511 139 522 173
rect 466 101 522 139
rect 466 67 477 101
rect 511 67 522 101
rect 466 36 522 67
rect 552 173 608 204
rect 552 139 563 173
rect 597 139 608 173
rect 552 101 608 139
rect 552 67 563 101
rect 597 67 608 101
rect 552 36 608 67
<< ndiffc >>
rect 47 139 81 173
rect 47 67 81 101
rect 133 139 167 173
rect 133 67 167 101
rect 219 139 253 173
rect 219 67 253 101
rect 305 139 339 173
rect 305 67 339 101
rect 391 139 425 173
rect 391 67 425 101
rect 477 139 511 173
rect 477 67 511 101
rect 563 139 597 173
rect 563 67 597 101
<< poly >>
rect 92 285 552 301
rect 92 251 135 285
rect 169 251 203 285
rect 237 251 271 285
rect 305 251 339 285
rect 373 251 407 285
rect 441 251 475 285
rect 509 251 552 285
rect 92 230 552 251
rect 92 204 122 230
rect 178 204 208 230
rect 264 204 294 230
rect 350 204 380 230
rect 436 204 466 230
rect 522 204 552 230
rect 92 10 122 36
rect 178 10 208 36
rect 264 10 294 36
rect 350 10 380 36
rect 436 10 466 36
rect 522 10 552 36
<< polycont >>
rect 135 251 169 285
rect 203 251 237 285
rect 271 251 305 285
rect 339 251 373 285
rect 407 251 441 285
rect 475 251 509 285
<< locali >>
rect 119 285 525 301
rect 119 251 125 285
rect 169 251 197 285
rect 237 251 269 285
rect 305 251 339 285
rect 375 251 407 285
rect 447 251 475 285
rect 519 251 525 285
rect 119 235 525 251
rect 47 173 81 189
rect 47 101 81 139
rect 47 51 81 67
rect 133 173 167 189
rect 133 101 167 139
rect 133 51 167 67
rect 219 173 253 189
rect 219 101 253 139
rect 219 51 253 67
rect 305 173 339 189
rect 305 101 339 139
rect 305 51 339 67
rect 391 173 425 189
rect 391 101 425 139
rect 391 51 425 67
rect 477 173 511 189
rect 477 101 511 139
rect 477 51 511 67
rect 563 173 597 189
rect 563 101 597 139
rect 563 51 597 67
<< viali >>
rect 125 251 135 285
rect 135 251 159 285
rect 197 251 203 285
rect 203 251 231 285
rect 269 251 271 285
rect 271 251 303 285
rect 341 251 373 285
rect 373 251 375 285
rect 413 251 441 285
rect 441 251 447 285
rect 485 251 509 285
rect 509 251 519 285
rect 47 139 81 173
rect 47 67 81 101
rect 133 139 167 173
rect 133 67 167 101
rect 219 139 253 173
rect 219 67 253 101
rect 305 139 339 173
rect 305 67 339 101
rect 391 139 425 173
rect 391 67 425 101
rect 477 139 511 173
rect 477 67 511 101
rect 563 139 597 173
rect 563 67 597 101
<< metal1 >>
rect 113 285 531 297
rect 113 251 125 285
rect 159 251 197 285
rect 231 251 269 285
rect 303 251 341 285
rect 375 251 413 285
rect 447 251 485 285
rect 519 251 531 285
rect 113 239 531 251
rect 41 173 87 189
rect 41 139 47 173
rect 81 139 87 173
rect 41 101 87 139
rect 41 67 47 101
rect 81 67 87 101
rect 41 -29 87 67
rect 124 176 176 189
rect 124 112 176 124
rect 124 51 176 60
rect 213 173 259 189
rect 213 139 219 173
rect 253 139 259 173
rect 213 101 259 139
rect 213 67 219 101
rect 253 67 259 101
rect 213 -29 259 67
rect 296 176 348 189
rect 296 112 348 124
rect 296 51 348 60
rect 385 173 431 189
rect 385 139 391 173
rect 425 139 431 173
rect 385 101 431 139
rect 385 67 391 101
rect 425 67 431 101
rect 385 -29 431 67
rect 468 176 520 189
rect 468 112 520 124
rect 468 51 520 60
rect 557 173 603 189
rect 557 139 563 173
rect 597 139 603 173
rect 557 101 603 139
rect 557 67 563 101
rect 597 67 603 101
rect 557 -29 603 67
rect 41 -89 603 -29
<< via1 >>
rect 124 173 176 176
rect 124 139 133 173
rect 133 139 167 173
rect 167 139 176 173
rect 124 124 176 139
rect 124 101 176 112
rect 124 67 133 101
rect 133 67 167 101
rect 167 67 176 101
rect 124 60 176 67
rect 296 173 348 176
rect 296 139 305 173
rect 305 139 339 173
rect 339 139 348 173
rect 296 124 348 139
rect 296 101 348 112
rect 296 67 305 101
rect 305 67 339 101
rect 339 67 348 101
rect 296 60 348 67
rect 468 173 520 176
rect 468 139 477 173
rect 477 139 511 173
rect 511 139 520 173
rect 468 124 520 139
rect 468 101 520 112
rect 468 67 477 101
rect 477 67 511 101
rect 511 67 520 101
rect 468 60 520 67
<< metal2 >>
rect 117 186 183 195
rect 117 130 122 186
rect 178 130 183 186
rect 117 124 124 130
rect 176 124 183 130
rect 117 112 183 124
rect 117 106 124 112
rect 176 106 183 112
rect 117 50 122 106
rect 178 50 183 106
rect 117 41 183 50
rect 289 186 355 195
rect 289 130 294 186
rect 350 130 355 186
rect 289 124 296 130
rect 348 124 355 130
rect 289 112 355 124
rect 289 106 296 112
rect 348 106 355 112
rect 289 50 294 106
rect 350 50 355 106
rect 289 41 355 50
rect 461 186 527 195
rect 461 130 466 186
rect 522 130 527 186
rect 461 124 468 130
rect 520 124 527 130
rect 461 112 527 124
rect 461 106 468 112
rect 520 106 527 112
rect 461 50 466 106
rect 522 50 527 106
rect 461 41 527 50
<< via2 >>
rect 122 176 178 186
rect 122 130 124 176
rect 124 130 176 176
rect 176 130 178 176
rect 122 60 124 106
rect 124 60 176 106
rect 176 60 178 106
rect 122 50 178 60
rect 294 176 350 186
rect 294 130 296 176
rect 296 130 348 176
rect 348 130 350 176
rect 294 60 296 106
rect 296 60 348 106
rect 348 60 350 106
rect 294 50 350 60
rect 466 176 522 186
rect 466 130 468 176
rect 468 130 520 176
rect 520 130 522 176
rect 466 60 468 106
rect 468 60 520 106
rect 520 60 522 106
rect 466 50 522 60
<< metal3 >>
rect 117 186 527 195
rect 117 130 122 186
rect 178 130 294 186
rect 350 130 466 186
rect 522 130 527 186
rect 117 129 527 130
rect 117 106 183 129
rect 117 50 122 106
rect 178 50 183 106
rect 117 41 183 50
rect 289 106 355 129
rect 289 50 294 106
rect 350 50 355 106
rect 289 41 355 50
rect 461 106 527 129
rect 461 50 466 106
rect 522 50 527 106
rect 461 41 527 50
<< labels >>
flabel metal3 s 117 129 527 195 0 FreeSans 400 0 0 0 DRAIN
port 1 nsew
flabel metal1 s 41 -89 603 -29 0 FreeSans 400 0 0 0 SOURCE
port 2 nsew
flabel metal1 s 113 239 531 297 0 FreeSans 400 0 0 0 GATE
port 3 nsew
flabel pwell s 73 210 89 225 0 FreeSans 200 0 0 0 SUBSTRATE
port 4 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 5909170
string GDS_START 5899892
string path 1.600 4.725 1.600 -2.225 
<< end >>
