magic
tech sky130A
magscale 1 2
timestamp 1624884095
<< checkpaint >>
rect -1525 -1260 9355 1760
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_0
timestamp 1624884095
transform -1 0 -165 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_1
timestamp 1624884095
transform 1 0 471 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_2
timestamp 1624884095
transform 1 0 1307 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_3
timestamp 1624884095
transform 1 0 2143 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_4
timestamp 1624884095
transform 1 0 2979 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_5
timestamp 1624884095
transform 1 0 3815 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_6
timestamp 1624884095
transform 1 0 4651 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_7
timestamp 1624884095
transform 1 0 5487 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_8
timestamp 1624884095
transform 1 0 6323 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_9
timestamp 1624884095
transform 1 0 7159 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_10
timestamp 1624884095
transform 1 0 7995 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 8095 471 8095 471 0 FreeSans 300 0 0 0 S
flabel comment s 7677 500 7677 500 0 FreeSans 300 0 0 0 D
flabel comment s 7259 471 7259 471 0 FreeSans 300 0 0 0 S
flabel comment s 6841 500 6841 500 0 FreeSans 300 0 0 0 D
flabel comment s 6423 471 6423 471 0 FreeSans 300 0 0 0 S
flabel comment s 6005 500 6005 500 0 FreeSans 300 0 0 0 D
flabel comment s 5587 471 5587 471 0 FreeSans 300 0 0 0 S
flabel comment s 5169 500 5169 500 0 FreeSans 300 0 0 0 D
flabel comment s 4751 471 4751 471 0 FreeSans 300 0 0 0 S
flabel comment s 4333 500 4333 500 0 FreeSans 300 0 0 0 D
flabel comment s 3915 471 3915 471 0 FreeSans 300 0 0 0 S
flabel comment s 3497 500 3497 500 0 FreeSans 300 0 0 0 D
flabel comment s 3079 471 3079 471 0 FreeSans 300 0 0 0 S
flabel comment s 2661 500 2661 500 0 FreeSans 300 0 0 0 D
flabel comment s 2243 471 2243 471 0 FreeSans 300 0 0 0 S
flabel comment s 1825 500 1825 500 0 FreeSans 300 0 0 0 D
flabel comment s 1407 471 1407 471 0 FreeSans 300 0 0 0 S
flabel comment s 989 500 989 500 0 FreeSans 300 0 0 0 D
flabel comment s 571 471 571 471 0 FreeSans 300 0 0 0 S
flabel comment s 153 500 153 500 0 FreeSans 300 0 0 0 D
flabel comment s -265 471 -265 471 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 17335378
string GDS_START 17324772
<< end >>
