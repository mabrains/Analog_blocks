magic
tech sky130A
magscale 1 2
timestamp 1624884095
<< checkpaint >>
rect -1430 -1857 4690 1781
<< pwell >>
rect -170 444 -84 521
rect -170 -120 3430 444
rect -170 -597 -84 -120
<< mvnmos >>
rect 92 334 1692 418
rect 1748 334 3348 418
rect 92 120 1692 204
rect 1748 120 3348 204
rect 92 -94 1692 -10
rect 1748 -94 3348 -10
<< mvndiff >>
rect 36 406 92 418
rect 36 372 47 406
rect 81 372 92 406
rect 36 334 92 372
rect 1692 406 1748 418
rect 1692 372 1703 406
rect 1737 372 1748 406
rect 1692 334 1748 372
rect 3348 406 3404 418
rect 3348 372 3359 406
rect 3393 372 3404 406
rect 3348 334 3404 372
rect 36 192 92 204
rect 36 158 47 192
rect 81 158 92 192
rect 36 120 92 158
rect 1692 192 1748 204
rect 1692 158 1703 192
rect 1737 158 1748 192
rect 1692 120 1748 158
rect 3348 192 3404 204
rect 3348 158 3359 192
rect 3393 158 3404 192
rect 3348 120 3404 158
rect 36 -48 92 -10
rect 36 -82 47 -48
rect 81 -82 92 -48
rect 36 -94 92 -82
rect 1692 -48 1748 -10
rect 1692 -82 1703 -48
rect 1737 -82 1748 -48
rect 1692 -94 1748 -82
rect 3348 -48 3404 -10
rect 3348 -82 3359 -48
rect 3393 -82 3404 -48
rect 3348 -94 3404 -82
<< mvndiffc >>
rect 47 372 81 406
rect 1703 372 1737 406
rect 3359 372 3393 406
rect 47 158 81 192
rect 1703 158 1737 192
rect 3359 158 3393 192
rect 47 -82 81 -48
rect 1703 -82 1737 -48
rect 3359 -82 3393 -48
<< psubdiff >>
rect -144 461 -110 495
rect -144 392 -110 427
rect -144 323 -110 358
rect -144 254 -110 289
rect -144 185 -110 220
rect -144 116 -110 151
rect -144 47 -110 82
rect -144 -22 -110 13
rect -144 -91 -110 -56
rect -144 -160 -110 -125
rect -144 -229 -110 -194
rect -144 -298 -110 -263
rect -144 -367 -110 -332
rect -144 -435 -110 -401
rect -144 -503 -110 -469
rect -144 -571 -110 -537
<< psubdiffcont >>
rect -144 427 -110 461
rect -144 358 -110 392
rect -144 289 -110 323
rect -144 220 -110 254
rect -144 151 -110 185
rect -144 82 -110 116
rect -144 13 -110 47
rect -144 -56 -110 -22
rect -144 -125 -110 -91
rect -144 -194 -110 -160
rect -144 -263 -110 -229
rect -144 -332 -110 -298
rect -144 -401 -110 -367
rect -144 -469 -110 -435
rect -144 -537 -110 -503
<< poly >>
rect 92 418 1692 450
rect 1748 418 3348 450
rect 92 302 1692 334
rect 1748 302 3348 334
rect 92 286 3348 302
rect 92 252 108 286
rect 142 252 178 286
rect 212 252 248 286
rect 282 252 318 286
rect 352 252 388 286
rect 422 252 458 286
rect 492 252 528 286
rect 562 252 598 286
rect 632 252 668 286
rect 702 252 738 286
rect 772 252 808 286
rect 842 252 878 286
rect 912 252 948 286
rect 982 252 1018 286
rect 1052 252 1088 286
rect 1122 252 1158 286
rect 1192 252 1228 286
rect 1262 252 1297 286
rect 1331 252 1366 286
rect 1400 252 1435 286
rect 1469 252 1504 286
rect 1538 252 1573 286
rect 1607 252 1642 286
rect 1676 252 1711 286
rect 1745 252 1780 286
rect 1814 252 1849 286
rect 1883 252 1918 286
rect 1952 252 1987 286
rect 2021 252 2056 286
rect 2090 252 2125 286
rect 2159 252 2194 286
rect 2228 252 2263 286
rect 2297 252 2332 286
rect 2366 252 2401 286
rect 2435 252 2470 286
rect 2504 252 2539 286
rect 2573 252 2608 286
rect 2642 252 2677 286
rect 2711 252 2746 286
rect 2780 252 2815 286
rect 2849 252 2884 286
rect 2918 252 2953 286
rect 2987 252 3022 286
rect 3056 252 3091 286
rect 3125 252 3160 286
rect 3194 252 3229 286
rect 3263 252 3298 286
rect 3332 252 3348 286
rect 92 236 3348 252
rect 92 204 1692 236
rect 1748 204 3348 236
rect 92 88 1692 120
rect 1748 88 3348 120
rect 92 72 3348 88
rect 92 38 108 72
rect 142 38 178 72
rect 212 38 248 72
rect 282 38 318 72
rect 352 38 388 72
rect 422 38 458 72
rect 492 38 528 72
rect 562 38 598 72
rect 632 38 668 72
rect 702 38 738 72
rect 772 38 808 72
rect 842 38 878 72
rect 912 38 948 72
rect 982 38 1018 72
rect 1052 38 1088 72
rect 1122 38 1158 72
rect 1192 38 1228 72
rect 1262 38 1297 72
rect 1331 38 1366 72
rect 1400 38 1435 72
rect 1469 38 1504 72
rect 1538 38 1573 72
rect 1607 38 1642 72
rect 1676 38 1711 72
rect 1745 38 1780 72
rect 1814 38 1849 72
rect 1883 38 1918 72
rect 1952 38 1987 72
rect 2021 38 2056 72
rect 2090 38 2125 72
rect 2159 38 2194 72
rect 2228 38 2263 72
rect 2297 38 2332 72
rect 2366 38 2401 72
rect 2435 38 2470 72
rect 2504 38 2539 72
rect 2573 38 2608 72
rect 2642 38 2677 72
rect 2711 38 2746 72
rect 2780 38 2815 72
rect 2849 38 2884 72
rect 2918 38 2953 72
rect 2987 38 3022 72
rect 3056 38 3091 72
rect 3125 38 3160 72
rect 3194 38 3229 72
rect 3263 38 3298 72
rect 3332 38 3348 72
rect 92 22 3348 38
rect 92 -10 1692 22
rect 1748 -10 3348 22
rect 92 -126 1692 -94
rect 1748 -126 3348 -94
<< polycont >>
rect 108 252 142 286
rect 178 252 212 286
rect 248 252 282 286
rect 318 252 352 286
rect 388 252 422 286
rect 458 252 492 286
rect 528 252 562 286
rect 598 252 632 286
rect 668 252 702 286
rect 738 252 772 286
rect 808 252 842 286
rect 878 252 912 286
rect 948 252 982 286
rect 1018 252 1052 286
rect 1088 252 1122 286
rect 1158 252 1192 286
rect 1228 252 1262 286
rect 1297 252 1331 286
rect 1366 252 1400 286
rect 1435 252 1469 286
rect 1504 252 1538 286
rect 1573 252 1607 286
rect 1642 252 1676 286
rect 1711 252 1745 286
rect 1780 252 1814 286
rect 1849 252 1883 286
rect 1918 252 1952 286
rect 1987 252 2021 286
rect 2056 252 2090 286
rect 2125 252 2159 286
rect 2194 252 2228 286
rect 2263 252 2297 286
rect 2332 252 2366 286
rect 2401 252 2435 286
rect 2470 252 2504 286
rect 2539 252 2573 286
rect 2608 252 2642 286
rect 2677 252 2711 286
rect 2746 252 2780 286
rect 2815 252 2849 286
rect 2884 252 2918 286
rect 2953 252 2987 286
rect 3022 252 3056 286
rect 3091 252 3125 286
rect 3160 252 3194 286
rect 3229 252 3263 286
rect 3298 252 3332 286
rect 108 38 142 72
rect 178 38 212 72
rect 248 38 282 72
rect 318 38 352 72
rect 388 38 422 72
rect 458 38 492 72
rect 528 38 562 72
rect 598 38 632 72
rect 668 38 702 72
rect 738 38 772 72
rect 808 38 842 72
rect 878 38 912 72
rect 948 38 982 72
rect 1018 38 1052 72
rect 1088 38 1122 72
rect 1158 38 1192 72
rect 1228 38 1262 72
rect 1297 38 1331 72
rect 1366 38 1400 72
rect 1435 38 1469 72
rect 1504 38 1538 72
rect 1573 38 1607 72
rect 1642 38 1676 72
rect 1711 38 1745 72
rect 1780 38 1814 72
rect 1849 38 1883 72
rect 1918 38 1952 72
rect 1987 38 2021 72
rect 2056 38 2090 72
rect 2125 38 2159 72
rect 2194 38 2228 72
rect 2263 38 2297 72
rect 2332 38 2366 72
rect 2401 38 2435 72
rect 2470 38 2504 72
rect 2539 38 2573 72
rect 2608 38 2642 72
rect 2677 38 2711 72
rect 2746 38 2780 72
rect 2815 38 2849 72
rect 2884 38 2918 72
rect 2953 38 2987 72
rect 3022 38 3056 72
rect 3091 38 3125 72
rect 3160 38 3194 72
rect 3229 38 3263 72
rect 3298 38 3332 72
<< locali >>
rect -144 461 -110 495
rect -144 421 -110 427
rect -144 344 -110 358
rect 81 388 119 422
rect 1737 388 1775 422
rect 3321 388 3359 422
rect 47 356 81 372
rect 1703 356 1737 372
rect 3359 356 3393 372
rect -144 267 -110 289
rect 92 252 108 286
rect 142 252 178 286
rect 212 252 248 286
rect 282 252 318 286
rect 352 252 388 286
rect 422 252 458 286
rect 492 252 528 286
rect 562 252 598 286
rect 632 252 668 286
rect 702 252 738 286
rect 772 252 808 286
rect 842 252 878 286
rect 912 252 948 286
rect 982 252 1018 286
rect 1052 252 1088 286
rect 1122 252 1158 286
rect 1192 252 1228 286
rect 1262 252 1297 286
rect 1331 252 1366 286
rect 1400 252 1435 286
rect 1469 252 1504 286
rect 1538 252 1573 286
rect 1607 252 1642 286
rect 1676 252 1711 286
rect 1745 252 1780 286
rect 1814 252 1849 286
rect 1883 252 1918 286
rect 1952 252 1987 286
rect 2021 252 2056 286
rect 2090 252 2125 286
rect 2159 252 2194 286
rect 2228 252 2263 286
rect 2297 252 2332 286
rect 2366 252 2401 286
rect 2435 252 2470 286
rect 2504 252 2539 286
rect 2573 252 2608 286
rect 2642 252 2677 286
rect 2711 252 2746 286
rect 2780 252 2815 286
rect 2849 252 2884 286
rect 2918 252 2953 286
rect 2987 252 3022 286
rect 3056 252 3091 286
rect 3125 252 3160 286
rect 3194 252 3229 286
rect 3263 252 3298 286
rect 3332 252 3348 286
rect -144 190 -110 220
rect -144 116 -110 151
rect 81 174 119 208
rect 47 142 81 158
rect -144 47 -110 80
rect 339 72 1534 252
rect 1665 174 1703 208
rect 1703 142 1737 158
rect 1837 72 3125 252
rect 3321 174 3359 208
rect 3359 142 3393 158
rect 92 38 108 72
rect 142 38 178 72
rect 212 38 248 72
rect 282 38 318 72
rect 352 38 388 72
rect 422 38 458 72
rect 492 38 528 72
rect 562 38 598 72
rect 632 38 668 72
rect 702 38 738 72
rect 772 38 808 72
rect 842 38 878 72
rect 912 38 948 72
rect 982 38 1018 72
rect 1052 38 1088 72
rect 1122 38 1158 72
rect 1192 38 1228 72
rect 1262 38 1297 72
rect 1331 38 1366 72
rect 1400 38 1435 72
rect 1469 38 1504 72
rect 1538 38 1573 72
rect 1607 38 1642 72
rect 1676 38 1711 72
rect 1745 38 1780 72
rect 1814 38 1849 72
rect 1883 38 1918 72
rect 1952 38 1987 72
rect 2021 38 2056 72
rect 2090 38 2125 72
rect 2159 38 2194 72
rect 2228 38 2263 72
rect 2297 38 2332 72
rect 2366 38 2401 72
rect 2435 38 2470 72
rect 2504 38 2539 72
rect 2573 38 2608 72
rect 2642 38 2677 72
rect 2711 38 2746 72
rect 2780 38 2815 72
rect 2849 38 2884 72
rect 2918 38 2953 72
rect 2987 38 3022 72
rect 3056 38 3091 72
rect 3125 38 3160 72
rect 3194 38 3229 72
rect 3263 38 3298 72
rect 3332 38 3348 72
rect -144 -22 -110 4
rect -144 -91 -110 -72
rect 47 -48 81 -32
rect 1703 -48 1737 -32
rect 3359 -48 3393 -32
rect 81 -98 119 -64
rect 1737 -98 1775 -64
rect 3321 -98 3359 -64
rect -144 -160 -110 -148
rect -144 -229 -110 -224
rect -144 -266 -110 -263
rect -144 -342 -110 -332
rect -144 -418 -110 -401
rect -144 -494 -110 -469
rect -144 -571 -110 -537
<< viali >>
rect -144 392 -110 421
rect -144 387 -110 392
rect 47 406 81 422
rect 47 388 81 406
rect 119 388 153 422
rect 1703 406 1737 422
rect 1703 388 1737 406
rect 1775 388 1809 422
rect 3287 388 3321 422
rect 3359 406 3393 422
rect 3359 388 3393 406
rect -144 323 -110 344
rect -144 310 -110 323
rect -144 254 -110 267
rect -144 233 -110 254
rect -144 185 -110 190
rect -144 156 -110 185
rect 47 192 81 208
rect 47 174 81 192
rect 119 174 153 208
rect -144 82 -110 114
rect -144 80 -110 82
rect 1631 174 1665 208
rect 1703 192 1737 208
rect 1703 174 1737 192
rect 3287 174 3321 208
rect 3359 192 3393 208
rect 3359 174 3393 192
rect -144 13 -110 38
rect -144 4 -110 13
rect -144 -56 -110 -38
rect -144 -72 -110 -56
rect 47 -82 81 -64
rect 47 -98 81 -82
rect 119 -98 153 -64
rect 1703 -82 1737 -64
rect 1703 -98 1737 -82
rect 1775 -98 1809 -64
rect 3287 -98 3321 -64
rect 3359 -82 3393 -64
rect 3359 -98 3393 -82
rect -144 -125 -110 -114
rect -144 -148 -110 -125
rect -144 -194 -110 -190
rect -144 -224 -110 -194
rect -144 -298 -110 -266
rect -144 -300 -110 -298
rect -144 -367 -110 -342
rect -144 -376 -110 -367
rect -144 -435 -110 -418
rect -144 -452 -110 -435
rect -144 -503 -110 -494
rect -144 -528 -110 -503
<< metal1 >>
rect -104 433 726 434
rect -150 422 726 433
rect -150 421 47 422
rect -150 387 -144 421
rect -110 388 47 421
rect 81 388 119 422
rect 153 388 726 422
rect -110 387 726 388
rect -150 376 726 387
rect 727 377 728 433
rect 768 377 769 433
rect 770 422 2382 434
rect 770 388 1703 422
rect 1737 388 1775 422
rect 1809 388 2382 422
rect 770 376 2382 388
rect 2383 377 2384 433
rect 2424 377 2425 433
rect 2426 428 3399 434
rect 2426 422 3405 428
rect 2426 388 3287 422
rect 3321 388 3359 422
rect 3393 388 3405 422
rect 2426 376 3405 388
rect -150 344 -104 376
rect -150 310 -144 344
rect -110 310 -104 344
rect -150 267 -104 310
rect -150 233 -144 267
rect -110 233 -104 267
rect -150 190 -104 233
rect 3353 220 3405 376
rect -150 156 -144 190
rect -110 156 -104 190
rect -150 114 -104 156
rect -150 80 -144 114
rect -110 80 -104 114
rect -150 38 -104 80
rect -150 4 -144 38
rect -110 4 -104 38
rect -150 -38 -104 4
rect -150 -72 -144 -38
rect -110 -72 -104 -38
rect -150 -114 -104 -72
rect 35 208 726 220
rect 35 174 47 208
rect 81 174 119 208
rect 153 174 726 208
rect 35 162 726 174
rect 727 163 728 219
rect 768 163 769 219
rect 770 208 2382 220
rect 770 174 1631 208
rect 1665 174 1703 208
rect 1737 174 2382 208
rect 770 162 2382 174
rect 2383 163 2384 219
rect 2424 163 2425 219
rect 2426 208 3405 220
rect 2426 174 3287 208
rect 3321 174 3359 208
rect 3393 174 3405 208
rect 2426 162 3405 174
rect 35 -52 87 162
tri 1029 -52 1079 -2 se
rect 1079 -52 1532 -2
tri 1532 -52 1582 -2 sw
rect 35 -64 726 -52
rect 35 -98 47 -64
rect 81 -98 119 -64
rect 153 -98 726 -64
rect 35 -104 726 -98
rect 41 -110 726 -104
rect 727 -109 728 -53
rect 768 -109 769 -53
rect 770 -60 2382 -52
rect 770 -64 1099 -60
tri 1099 -64 1103 -60 nw
tri 1508 -64 1512 -60 ne
rect 1512 -64 2382 -60
rect 770 -98 1065 -64
tri 1065 -98 1099 -64 nw
tri 1512 -98 1546 -64 ne
rect 1546 -98 1703 -64
rect 1737 -98 1775 -64
rect 1809 -98 2382 -64
rect 770 -110 1053 -98
tri 1053 -110 1065 -98 nw
tri 1546 -110 1558 -98 ne
rect 1558 -110 2382 -98
rect 2383 -109 2384 -53
rect 2424 -109 2425 -53
rect 2426 -64 3405 -52
rect 2426 -98 3287 -64
rect 3321 -98 3359 -64
rect 3393 -98 3405 -64
rect 2426 -110 3405 -98
rect -150 -148 -144 -114
rect -110 -148 -104 -114
rect -150 -190 -104 -148
rect -150 -224 -144 -190
rect -110 -224 -104 -190
rect -150 -266 -104 -224
rect -150 -300 -144 -266
rect -110 -300 -104 -266
rect -150 -342 -104 -300
rect -150 -376 -144 -342
rect -110 -376 -104 -342
rect -150 -418 -104 -376
rect -150 -452 -144 -418
rect -110 -452 -104 -418
rect -150 -494 -104 -452
rect -150 -528 -144 -494
rect -110 -528 -104 -494
rect -150 -540 -104 -528
<< rmetal1 >>
rect 726 433 728 434
rect 726 377 727 433
rect 726 376 728 377
rect 768 433 770 434
rect 769 377 770 433
rect 2382 433 2384 434
rect 768 376 770 377
rect 2382 377 2383 433
rect 2382 376 2384 377
rect 2424 433 2426 434
rect 2425 377 2426 433
rect 2424 376 2426 377
rect 726 219 728 220
rect 726 163 727 219
rect 726 162 728 163
rect 768 219 770 220
rect 769 163 770 219
rect 2382 219 2384 220
rect 768 162 770 163
rect 2382 163 2383 219
rect 2382 162 2384 163
rect 2424 219 2426 220
rect 2425 163 2426 219
rect 2424 162 2426 163
rect 726 -53 728 -52
rect 726 -109 727 -53
rect 726 -110 728 -109
rect 768 -53 770 -52
rect 769 -109 770 -53
rect 2382 -53 2384 -52
rect 768 -110 770 -109
rect 2382 -109 2383 -53
rect 2382 -110 2384 -109
rect 2424 -53 2426 -52
rect 2425 -109 2426 -53
rect 2424 -110 2426 -109
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1624884095
transform 1 0 47 0 1 -98
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1624884095
transform 1 0 47 0 1 174
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1624884095
transform 1 0 1703 0 1 -98
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1624884095
transform 1 0 1631 0 1 174
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_4
timestamp 1624884095
transform 1 0 3287 0 1 -98
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_5
timestamp 1624884095
transform 1 0 3287 0 1 174
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_6
timestamp 1624884095
transform 1 0 3287 0 1 388
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_7
timestamp 1624884095
transform 1 0 1703 0 1 388
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_8
timestamp 1624884095
transform 1 0 47 0 1 388
box 0 0 1 1
use sky130_fd_io__tk_em1o_cdns_5595914180891  sky130_fd_io__tk_em1o_cdns_5595914180891_0
timestamp 1624884095
transform 1 0 2330 0 1 376
box 0 24 148 28
use sky130_fd_io__tk_em1o_cdns_5595914180891  sky130_fd_io__tk_em1o_cdns_5595914180891_1
timestamp 1624884095
transform 1 0 2330 0 1 162
box 0 24 148 28
use sky130_fd_io__tk_em1o_cdns_5595914180891  sky130_fd_io__tk_em1o_cdns_5595914180891_2
timestamp 1624884095
transform 1 0 674 0 1 162
box 0 24 148 28
use sky130_fd_io__tk_em1o_cdns_5595914180891  sky130_fd_io__tk_em1o_cdns_5595914180891_3
timestamp 1624884095
transform 1 0 2330 0 1 -110
box 0 24 148 28
use sky130_fd_io__tk_em1o_cdns_5595914180891  sky130_fd_io__tk_em1o_cdns_5595914180891_4
timestamp 1624884095
transform 1 0 674 0 1 -110
box 0 24 148 28
use sky130_fd_io__tk_em1o_cdns_5595914180891  sky130_fd_io__tk_em1o_cdns_5595914180891_5
timestamp 1624884095
transform 1 0 674 0 1 376
box 0 24 148 28
use sky130_fd_pr__nfet_01v8__example_5595914180889  sky130_fd_pr__nfet_01v8__example_5595914180889_0
timestamp 1624884095
transform 1 0 92 0 -1 418
box -28 0 3284 13
use sky130_fd_pr__nfet_01v8__example_5595914180889  sky130_fd_pr__nfet_01v8__example_5595914180889_1
timestamp 1624884095
transform 1 0 92 0 -1 204
box -28 0 3284 13
use sky130_fd_pr__nfet_01v8__example_5595914180889  sky130_fd_pr__nfet_01v8__example_5595914180889_2
timestamp 1624884095
transform 1 0 92 0 1 -94
box -28 0 3284 13
<< labels >>
flabel metal1 s 3318 -107 3382 -56 3 FreeSans 520 0 0 0 OUT
port 1 nsew
flabel metal1 s 57 380 151 426 3 FreeSans 520 0 0 0 VGND
port 2 nsew
flabel locali s 722 85 907 204 3 FreeSans 520 0 0 0 E_N
port 3 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 40016964
string GDS_START 40005438
<< end >>
