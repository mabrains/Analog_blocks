magic
tech sky130A
magscale 1 2
timestamp 1624884095
<< checkpaint >>
rect -1302 -1236 1970 2376
<< nwell >>
rect -42 415 710 1116
<< pwell >>
rect 40 118 494 310
<< mvnmos >>
rect 119 144 239 284
rect 295 144 415 284
<< mvpmos >>
rect 119 750 239 950
rect 295 750 415 950
rect 471 750 591 950
rect 119 482 239 682
rect 295 482 415 682
rect 471 482 591 682
<< mvndiff >>
rect 66 272 119 284
rect 66 238 74 272
rect 108 238 119 272
rect 66 204 119 238
rect 66 170 74 204
rect 108 170 119 204
rect 66 144 119 170
rect 239 144 295 284
rect 415 272 468 284
rect 415 238 426 272
rect 460 238 468 272
rect 415 204 468 238
rect 415 170 426 204
rect 460 170 468 204
rect 415 144 468 170
<< mvpdiff >>
rect 66 932 119 950
rect 66 898 74 932
rect 108 898 119 932
rect 66 864 119 898
rect 66 830 74 864
rect 108 830 119 864
rect 66 796 119 830
rect 66 762 74 796
rect 108 762 119 796
rect 66 750 119 762
rect 239 932 295 950
rect 239 898 250 932
rect 284 898 295 932
rect 239 864 295 898
rect 239 830 250 864
rect 284 830 295 864
rect 239 796 295 830
rect 239 762 250 796
rect 284 762 295 796
rect 239 750 295 762
rect 415 932 471 950
rect 415 898 426 932
rect 460 898 471 932
rect 415 864 471 898
rect 415 830 426 864
rect 460 830 471 864
rect 415 796 471 830
rect 415 762 426 796
rect 460 762 471 796
rect 415 750 471 762
rect 591 932 644 950
rect 591 898 602 932
rect 636 898 644 932
rect 591 864 644 898
rect 591 830 602 864
rect 636 830 644 864
rect 591 796 644 830
rect 591 762 602 796
rect 636 762 644 796
rect 591 750 644 762
rect 66 664 119 682
rect 66 630 74 664
rect 108 630 119 664
rect 66 596 119 630
rect 66 562 74 596
rect 108 562 119 596
rect 66 528 119 562
rect 66 494 74 528
rect 108 494 119 528
rect 66 482 119 494
rect 239 664 295 682
rect 239 630 250 664
rect 284 630 295 664
rect 239 596 295 630
rect 239 562 250 596
rect 284 562 295 596
rect 239 528 295 562
rect 239 494 250 528
rect 284 494 295 528
rect 239 482 295 494
rect 415 664 471 682
rect 415 630 426 664
rect 460 630 471 664
rect 415 596 471 630
rect 415 562 426 596
rect 460 562 471 596
rect 415 528 471 562
rect 415 494 426 528
rect 460 494 471 528
rect 415 482 471 494
rect 591 664 644 682
rect 591 630 602 664
rect 636 630 644 664
rect 591 596 644 630
rect 591 562 602 596
rect 636 562 644 596
rect 591 528 644 562
rect 591 494 602 528
rect 636 494 644 528
rect 591 482 644 494
<< mvndiffc >>
rect 74 238 108 272
rect 74 170 108 204
rect 426 238 460 272
rect 426 170 460 204
<< mvpdiffc >>
rect 74 898 108 932
rect 74 830 108 864
rect 74 762 108 796
rect 250 898 284 932
rect 250 830 284 864
rect 250 762 284 796
rect 426 898 460 932
rect 426 830 460 864
rect 426 762 460 796
rect 602 898 636 932
rect 602 830 636 864
rect 602 762 636 796
rect 74 630 108 664
rect 74 562 108 596
rect 74 494 108 528
rect 250 630 284 664
rect 250 562 284 596
rect 250 494 284 528
rect 426 630 460 664
rect 426 562 460 596
rect 426 494 460 528
rect 602 630 636 664
rect 602 562 636 596
rect 602 494 636 528
<< poly >>
rect 119 950 239 976
rect 295 950 415 976
rect 471 950 591 976
rect 119 724 239 750
rect 295 724 415 750
rect 471 724 591 750
rect 119 682 239 708
rect 295 682 415 708
rect 471 682 591 708
rect 119 456 239 482
rect 295 456 415 482
rect 471 456 591 482
rect 119 432 591 456
rect 119 398 165 432
rect 199 398 336 432
rect 370 398 591 432
rect 119 364 591 398
rect 119 330 165 364
rect 199 330 336 364
rect 370 330 591 364
rect 119 310 591 330
rect 119 284 239 310
rect 295 284 415 310
rect 119 118 239 144
rect 295 118 415 144
<< polycont >>
rect 165 398 199 432
rect 336 398 370 432
rect 165 330 199 364
rect 336 330 370 364
<< locali >>
rect 74 932 108 944
rect 74 864 108 872
rect 74 796 108 830
rect 74 664 108 762
rect 74 596 108 630
rect 74 528 108 562
rect 74 478 108 494
rect 250 932 284 950
rect 250 864 284 898
rect 250 796 284 830
rect 250 664 284 762
rect 250 596 284 630
rect 250 528 284 562
rect 149 398 165 432
rect 199 398 215 432
rect 149 364 215 398
rect 149 330 165 364
rect 199 330 215 364
rect 74 272 108 288
rect 74 227 108 238
rect 250 261 284 494
rect 426 932 460 944
rect 426 864 460 872
rect 426 796 460 830
rect 426 664 460 762
rect 426 596 460 630
rect 426 528 460 562
rect 426 478 460 494
rect 602 932 636 948
rect 602 864 636 898
rect 602 796 636 830
rect 602 664 636 762
rect 602 596 636 630
rect 602 528 636 562
rect 320 398 336 432
rect 370 398 386 432
rect 320 364 386 398
rect 320 330 336 364
rect 370 330 386 364
rect 426 272 460 288
rect 250 238 426 261
rect 602 238 636 494
rect 250 227 636 238
rect 74 155 108 170
rect 421 204 636 227
rect 421 170 426 204
rect 421 154 460 170
<< viali >>
rect 74 944 108 978
rect 74 898 108 906
rect 74 872 108 898
rect 426 944 460 978
rect 426 898 460 906
rect 426 872 460 898
rect 74 204 108 227
rect 74 193 108 204
rect 74 121 108 155
<< metal1 >>
rect 25 978 644 1062
rect 25 944 74 978
rect 108 944 426 978
rect 460 944 644 978
rect 25 906 644 944
rect 25 872 74 906
rect 108 872 426 906
rect 460 872 644 906
rect 25 859 644 872
rect 24 227 503 239
rect 24 193 74 227
rect 108 193 503 227
rect 24 155 503 193
rect 24 121 74 155
rect 108 121 503 155
rect 24 24 503 121
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1624884095
transform 0 -1 108 1 0 872
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1624884095
transform 0 -1 460 1 0 872
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1624884095
transform 0 -1 108 -1 0 227
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_0
timestamp 1624884095
transform 0 1 149 -1 0 448
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_1
timestamp 1624884095
transform 0 1 320 -1 0 448
box 0 0 1 1
use sky130_fd_pr__nfet_01v8__example_559591418089  sky130_fd_pr__nfet_01v8__example_559591418089_0
timestamp 1624884095
transform 1 0 119 0 -1 284
box -28 0 145 70
use sky130_fd_pr__nfet_01v8__example_559591418087  sky130_fd_pr__nfet_01v8__example_559591418087_0
timestamp 1624884095
transform 1 0 295 0 -1 284
box -25 0 148 70
use sky130_fd_pr__pfet_01v8__example_559591418085  sky130_fd_pr__pfet_01v8__example_559591418085_0
timestamp 1624884095
transform 1 0 119 0 1 750
box -28 0 148 97
use sky130_fd_pr__pfet_01v8__example_559591418085  sky130_fd_pr__pfet_01v8__example_559591418085_1
timestamp 1624884095
transform 1 0 295 0 1 750
box -28 0 148 97
use sky130_fd_pr__pfet_01v8__example_559591418085  sky130_fd_pr__pfet_01v8__example_559591418085_2
timestamp 1624884095
transform 1 0 119 0 1 482
box -28 0 148 97
use sky130_fd_pr__pfet_01v8__example_559591418085  sky130_fd_pr__pfet_01v8__example_559591418085_3
timestamp 1624884095
transform 1 0 471 0 1 482
box -28 0 148 97
use sky130_fd_pr__pfet_01v8__example_559591418085  sky130_fd_pr__pfet_01v8__example_559591418085_4
timestamp 1624884095
transform 1 0 471 0 1 750
box -28 0 148 97
use sky130_fd_pr__pfet_01v8__example_559591418085  sky130_fd_pr__pfet_01v8__example_559591418085_5
timestamp 1624884095
transform 1 0 295 0 1 482
box -28 0 148 97
<< labels >>
flabel locali s 321 352 383 391 0 FreeSans 400 0 0 0 IN1
port 1 nsew
flabel locali s 156 353 207 394 0 FreeSans 400 0 0 0 IN0
port 2 nsew
flabel locali s 250 256 284 532 0 FreeSans 200 0 0 0 OUT
port 3 nsew
flabel metal1 s 24 24 107 238 0 FreeSans 320 0 0 0 VGND
port 4 nsew
flabel metal1 s 561 859 644 1062 0 FreeSans 320 0 0 0 VPWR
port 5 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 35752958
string GDS_START 35750400
<< end >>
