magic
tech sky130A
magscale 1 2
timestamp 1624884095
<< checkpaint >>
rect -1310 -1333 11639 3689
<< dnwell >>
rect 3713 109 10299 2399
rect 3713 7 6890 109
<< nwell >>
rect 170 294 1560 2158
rect 1985 224 3349 2174
rect 3633 2311 10329 2429
rect 3633 2193 10379 2311
rect 3633 213 3919 2193
rect 6776 315 7010 2193
rect 10093 315 10379 2193
rect 6775 213 10379 315
rect 3633 79 10379 213
rect 3633 29 8312 79
rect 3633 -73 7011 29
<< pwell >>
rect -50 2234 3563 2388
rect -50 164 104 2234
rect 1621 164 1925 2234
rect 3409 164 3563 2234
rect -50 10 3563 164
rect 3979 307 6715 2099
rect 7071 409 10023 2133
<< mvnmos >>
rect 4176 475 4276 1875
rect 4346 475 4446 1875
rect 4502 475 4602 1875
rect 4672 475 4772 1875
rect 4828 475 4928 1875
rect 4998 475 5098 1875
rect 5154 475 5254 1875
rect 5447 475 5547 1875
rect 5603 475 5703 1875
rect 5773 475 5873 1875
rect 5929 475 6029 1875
rect 6099 475 6199 1875
rect 6255 475 6355 1875
rect 6425 475 6525 1875
rect 7261 543 7361 1943
rect 7431 543 7531 1943
rect 7587 543 7687 1943
rect 7757 543 7857 1943
rect 7913 543 8013 1943
rect 8083 543 8183 1943
rect 8239 543 8339 1943
rect 8532 543 8632 1943
rect 8688 543 8788 1943
rect 8858 543 8958 1943
rect 9014 543 9114 1943
rect 9184 543 9284 1943
rect 9340 543 9440 1943
rect 9510 543 9610 1943
rect 9666 543 9766 1943
<< mvpmos >>
rect 414 475 514 1875
rect 570 475 670 1875
rect 740 475 840 1875
rect 896 475 996 1875
rect 1066 475 1166 1875
rect 1222 475 1322 1875
rect 2291 475 2391 1875
rect 2461 475 2561 1875
rect 2617 475 2717 1875
rect 2787 475 2887 1875
rect 2943 475 3043 1875
<< mvndiff >>
rect 4120 1813 4176 1875
rect 4120 1779 4131 1813
rect 4165 1779 4176 1813
rect 4120 1745 4176 1779
rect 4120 1711 4131 1745
rect 4165 1711 4176 1745
rect 4120 1677 4176 1711
rect 4120 1643 4131 1677
rect 4165 1643 4176 1677
rect 4120 1609 4176 1643
rect 4120 1575 4131 1609
rect 4165 1575 4176 1609
rect 4120 1541 4176 1575
rect 4120 1507 4131 1541
rect 4165 1507 4176 1541
rect 4120 1473 4176 1507
rect 4120 1439 4131 1473
rect 4165 1439 4176 1473
rect 4120 1405 4176 1439
rect 4120 1371 4131 1405
rect 4165 1371 4176 1405
rect 4120 1337 4176 1371
rect 4120 1303 4131 1337
rect 4165 1303 4176 1337
rect 4120 1269 4176 1303
rect 4120 1235 4131 1269
rect 4165 1235 4176 1269
rect 4120 1201 4176 1235
rect 4120 1167 4131 1201
rect 4165 1167 4176 1201
rect 4120 1133 4176 1167
rect 4120 1099 4131 1133
rect 4165 1099 4176 1133
rect 4120 1065 4176 1099
rect 4120 1031 4131 1065
rect 4165 1031 4176 1065
rect 4120 997 4176 1031
rect 4120 963 4131 997
rect 4165 963 4176 997
rect 4120 929 4176 963
rect 4120 895 4131 929
rect 4165 895 4176 929
rect 4120 861 4176 895
rect 4120 827 4131 861
rect 4165 827 4176 861
rect 4120 793 4176 827
rect 4120 759 4131 793
rect 4165 759 4176 793
rect 4120 725 4176 759
rect 4120 691 4131 725
rect 4165 691 4176 725
rect 4120 657 4176 691
rect 4120 623 4131 657
rect 4165 623 4176 657
rect 4120 589 4176 623
rect 4120 555 4131 589
rect 4165 555 4176 589
rect 4120 521 4176 555
rect 4120 487 4131 521
rect 4165 487 4176 521
rect 4120 475 4176 487
rect 4276 1813 4346 1875
rect 4276 1779 4294 1813
rect 4328 1779 4346 1813
rect 4276 1745 4346 1779
rect 4276 1711 4294 1745
rect 4328 1711 4346 1745
rect 4276 1677 4346 1711
rect 4276 1643 4294 1677
rect 4328 1643 4346 1677
rect 4276 1609 4346 1643
rect 4276 1575 4294 1609
rect 4328 1575 4346 1609
rect 4276 1541 4346 1575
rect 4276 1507 4294 1541
rect 4328 1507 4346 1541
rect 4276 1473 4346 1507
rect 4276 1439 4294 1473
rect 4328 1439 4346 1473
rect 4276 1405 4346 1439
rect 4276 1371 4294 1405
rect 4328 1371 4346 1405
rect 4276 1337 4346 1371
rect 4276 1303 4294 1337
rect 4328 1303 4346 1337
rect 4276 1269 4346 1303
rect 4276 1235 4294 1269
rect 4328 1235 4346 1269
rect 4276 1201 4346 1235
rect 4276 1167 4294 1201
rect 4328 1167 4346 1201
rect 4276 1133 4346 1167
rect 4276 1099 4294 1133
rect 4328 1099 4346 1133
rect 4276 1065 4346 1099
rect 4276 1031 4294 1065
rect 4328 1031 4346 1065
rect 4276 997 4346 1031
rect 4276 963 4294 997
rect 4328 963 4346 997
rect 4276 929 4346 963
rect 4276 895 4294 929
rect 4328 895 4346 929
rect 4276 861 4346 895
rect 4276 827 4294 861
rect 4328 827 4346 861
rect 4276 793 4346 827
rect 4276 759 4294 793
rect 4328 759 4346 793
rect 4276 725 4346 759
rect 4276 691 4294 725
rect 4328 691 4346 725
rect 4276 657 4346 691
rect 4276 623 4294 657
rect 4328 623 4346 657
rect 4276 589 4346 623
rect 4276 555 4294 589
rect 4328 555 4346 589
rect 4276 521 4346 555
rect 4276 487 4294 521
rect 4328 487 4346 521
rect 4276 475 4346 487
rect 4446 1813 4502 1875
rect 4446 1779 4457 1813
rect 4491 1779 4502 1813
rect 4446 1745 4502 1779
rect 4446 1711 4457 1745
rect 4491 1711 4502 1745
rect 4446 1677 4502 1711
rect 4446 1643 4457 1677
rect 4491 1643 4502 1677
rect 4446 1609 4502 1643
rect 4446 1575 4457 1609
rect 4491 1575 4502 1609
rect 4446 1541 4502 1575
rect 4446 1507 4457 1541
rect 4491 1507 4502 1541
rect 4446 1473 4502 1507
rect 4446 1439 4457 1473
rect 4491 1439 4502 1473
rect 4446 1405 4502 1439
rect 4446 1371 4457 1405
rect 4491 1371 4502 1405
rect 4446 1337 4502 1371
rect 4446 1303 4457 1337
rect 4491 1303 4502 1337
rect 4446 1269 4502 1303
rect 4446 1235 4457 1269
rect 4491 1235 4502 1269
rect 4446 1201 4502 1235
rect 4446 1167 4457 1201
rect 4491 1167 4502 1201
rect 4446 1133 4502 1167
rect 4446 1099 4457 1133
rect 4491 1099 4502 1133
rect 4446 1065 4502 1099
rect 4446 1031 4457 1065
rect 4491 1031 4502 1065
rect 4446 997 4502 1031
rect 4446 963 4457 997
rect 4491 963 4502 997
rect 4446 929 4502 963
rect 4446 895 4457 929
rect 4491 895 4502 929
rect 4446 861 4502 895
rect 4446 827 4457 861
rect 4491 827 4502 861
rect 4446 793 4502 827
rect 4446 759 4457 793
rect 4491 759 4502 793
rect 4446 725 4502 759
rect 4446 691 4457 725
rect 4491 691 4502 725
rect 4446 657 4502 691
rect 4446 623 4457 657
rect 4491 623 4502 657
rect 4446 589 4502 623
rect 4446 555 4457 589
rect 4491 555 4502 589
rect 4446 521 4502 555
rect 4446 487 4457 521
rect 4491 487 4502 521
rect 4446 475 4502 487
rect 4602 1813 4672 1875
rect 4602 1779 4620 1813
rect 4654 1779 4672 1813
rect 4602 1745 4672 1779
rect 4602 1711 4620 1745
rect 4654 1711 4672 1745
rect 4602 1677 4672 1711
rect 4602 1643 4620 1677
rect 4654 1643 4672 1677
rect 4602 1609 4672 1643
rect 4602 1575 4620 1609
rect 4654 1575 4672 1609
rect 4602 1541 4672 1575
rect 4602 1507 4620 1541
rect 4654 1507 4672 1541
rect 4602 1473 4672 1507
rect 4602 1439 4620 1473
rect 4654 1439 4672 1473
rect 4602 1405 4672 1439
rect 4602 1371 4620 1405
rect 4654 1371 4672 1405
rect 4602 1337 4672 1371
rect 4602 1303 4620 1337
rect 4654 1303 4672 1337
rect 4602 1269 4672 1303
rect 4602 1235 4620 1269
rect 4654 1235 4672 1269
rect 4602 1201 4672 1235
rect 4602 1167 4620 1201
rect 4654 1167 4672 1201
rect 4602 1133 4672 1167
rect 4602 1099 4620 1133
rect 4654 1099 4672 1133
rect 4602 1065 4672 1099
rect 4602 1031 4620 1065
rect 4654 1031 4672 1065
rect 4602 997 4672 1031
rect 4602 963 4620 997
rect 4654 963 4672 997
rect 4602 929 4672 963
rect 4602 895 4620 929
rect 4654 895 4672 929
rect 4602 861 4672 895
rect 4602 827 4620 861
rect 4654 827 4672 861
rect 4602 793 4672 827
rect 4602 759 4620 793
rect 4654 759 4672 793
rect 4602 725 4672 759
rect 4602 691 4620 725
rect 4654 691 4672 725
rect 4602 657 4672 691
rect 4602 623 4620 657
rect 4654 623 4672 657
rect 4602 589 4672 623
rect 4602 555 4620 589
rect 4654 555 4672 589
rect 4602 521 4672 555
rect 4602 487 4620 521
rect 4654 487 4672 521
rect 4602 475 4672 487
rect 4772 1813 4828 1875
rect 4772 1779 4783 1813
rect 4817 1779 4828 1813
rect 4772 1745 4828 1779
rect 4772 1711 4783 1745
rect 4817 1711 4828 1745
rect 4772 1677 4828 1711
rect 4772 1643 4783 1677
rect 4817 1643 4828 1677
rect 4772 1609 4828 1643
rect 4772 1575 4783 1609
rect 4817 1575 4828 1609
rect 4772 1541 4828 1575
rect 4772 1507 4783 1541
rect 4817 1507 4828 1541
rect 4772 1473 4828 1507
rect 4772 1439 4783 1473
rect 4817 1439 4828 1473
rect 4772 1405 4828 1439
rect 4772 1371 4783 1405
rect 4817 1371 4828 1405
rect 4772 1337 4828 1371
rect 4772 1303 4783 1337
rect 4817 1303 4828 1337
rect 4772 1269 4828 1303
rect 4772 1235 4783 1269
rect 4817 1235 4828 1269
rect 4772 1201 4828 1235
rect 4772 1167 4783 1201
rect 4817 1167 4828 1201
rect 4772 1133 4828 1167
rect 4772 1099 4783 1133
rect 4817 1099 4828 1133
rect 4772 1065 4828 1099
rect 4772 1031 4783 1065
rect 4817 1031 4828 1065
rect 4772 997 4828 1031
rect 4772 963 4783 997
rect 4817 963 4828 997
rect 4772 929 4828 963
rect 4772 895 4783 929
rect 4817 895 4828 929
rect 4772 861 4828 895
rect 4772 827 4783 861
rect 4817 827 4828 861
rect 4772 793 4828 827
rect 4772 759 4783 793
rect 4817 759 4828 793
rect 4772 725 4828 759
rect 4772 691 4783 725
rect 4817 691 4828 725
rect 4772 657 4828 691
rect 4772 623 4783 657
rect 4817 623 4828 657
rect 4772 589 4828 623
rect 4772 555 4783 589
rect 4817 555 4828 589
rect 4772 521 4828 555
rect 4772 487 4783 521
rect 4817 487 4828 521
rect 4772 475 4828 487
rect 4928 1813 4998 1875
rect 4928 1779 4946 1813
rect 4980 1779 4998 1813
rect 4928 1745 4998 1779
rect 4928 1711 4946 1745
rect 4980 1711 4998 1745
rect 4928 1677 4998 1711
rect 4928 1643 4946 1677
rect 4980 1643 4998 1677
rect 4928 1609 4998 1643
rect 4928 1575 4946 1609
rect 4980 1575 4998 1609
rect 4928 1541 4998 1575
rect 4928 1507 4946 1541
rect 4980 1507 4998 1541
rect 4928 1473 4998 1507
rect 4928 1439 4946 1473
rect 4980 1439 4998 1473
rect 4928 1405 4998 1439
rect 4928 1371 4946 1405
rect 4980 1371 4998 1405
rect 4928 1337 4998 1371
rect 4928 1303 4946 1337
rect 4980 1303 4998 1337
rect 4928 1269 4998 1303
rect 4928 1235 4946 1269
rect 4980 1235 4998 1269
rect 4928 1201 4998 1235
rect 4928 1167 4946 1201
rect 4980 1167 4998 1201
rect 4928 1133 4998 1167
rect 4928 1099 4946 1133
rect 4980 1099 4998 1133
rect 4928 1065 4998 1099
rect 4928 1031 4946 1065
rect 4980 1031 4998 1065
rect 4928 997 4998 1031
rect 4928 963 4946 997
rect 4980 963 4998 997
rect 4928 929 4998 963
rect 4928 895 4946 929
rect 4980 895 4998 929
rect 4928 861 4998 895
rect 4928 827 4946 861
rect 4980 827 4998 861
rect 4928 793 4998 827
rect 4928 759 4946 793
rect 4980 759 4998 793
rect 4928 725 4998 759
rect 4928 691 4946 725
rect 4980 691 4998 725
rect 4928 657 4998 691
rect 4928 623 4946 657
rect 4980 623 4998 657
rect 4928 589 4998 623
rect 4928 555 4946 589
rect 4980 555 4998 589
rect 4928 521 4998 555
rect 4928 487 4946 521
rect 4980 487 4998 521
rect 4928 475 4998 487
rect 5098 1813 5154 1875
rect 5098 1779 5109 1813
rect 5143 1779 5154 1813
rect 5098 1745 5154 1779
rect 5098 1711 5109 1745
rect 5143 1711 5154 1745
rect 5098 1677 5154 1711
rect 5098 1643 5109 1677
rect 5143 1643 5154 1677
rect 5098 1609 5154 1643
rect 5098 1575 5109 1609
rect 5143 1575 5154 1609
rect 5098 1541 5154 1575
rect 5098 1507 5109 1541
rect 5143 1507 5154 1541
rect 5098 1473 5154 1507
rect 5098 1439 5109 1473
rect 5143 1439 5154 1473
rect 5098 1405 5154 1439
rect 5098 1371 5109 1405
rect 5143 1371 5154 1405
rect 5098 1337 5154 1371
rect 5098 1303 5109 1337
rect 5143 1303 5154 1337
rect 5098 1269 5154 1303
rect 5098 1235 5109 1269
rect 5143 1235 5154 1269
rect 5098 1201 5154 1235
rect 5098 1167 5109 1201
rect 5143 1167 5154 1201
rect 5098 1133 5154 1167
rect 5098 1099 5109 1133
rect 5143 1099 5154 1133
rect 5098 1065 5154 1099
rect 5098 1031 5109 1065
rect 5143 1031 5154 1065
rect 5098 997 5154 1031
rect 5098 963 5109 997
rect 5143 963 5154 997
rect 5098 929 5154 963
rect 5098 895 5109 929
rect 5143 895 5154 929
rect 5098 861 5154 895
rect 5098 827 5109 861
rect 5143 827 5154 861
rect 5098 793 5154 827
rect 5098 759 5109 793
rect 5143 759 5154 793
rect 5098 725 5154 759
rect 5098 691 5109 725
rect 5143 691 5154 725
rect 5098 657 5154 691
rect 5098 623 5109 657
rect 5143 623 5154 657
rect 5098 589 5154 623
rect 5098 555 5109 589
rect 5143 555 5154 589
rect 5098 521 5154 555
rect 5098 487 5109 521
rect 5143 487 5154 521
rect 5098 475 5154 487
rect 5254 1813 5317 1875
rect 5254 1779 5272 1813
rect 5306 1779 5317 1813
rect 5254 1745 5317 1779
rect 5254 1711 5272 1745
rect 5306 1711 5317 1745
rect 5254 1677 5317 1711
rect 5254 1643 5272 1677
rect 5306 1643 5317 1677
rect 5254 1609 5317 1643
rect 5254 1575 5272 1609
rect 5306 1575 5317 1609
rect 5254 1541 5317 1575
rect 5254 1507 5272 1541
rect 5306 1507 5317 1541
rect 5254 1473 5317 1507
rect 5254 1439 5272 1473
rect 5306 1439 5317 1473
rect 5254 1405 5317 1439
rect 5254 1371 5272 1405
rect 5306 1371 5317 1405
rect 5254 1337 5317 1371
rect 5254 1303 5272 1337
rect 5306 1303 5317 1337
rect 5254 1269 5317 1303
rect 5254 1235 5272 1269
rect 5306 1235 5317 1269
rect 5254 1201 5317 1235
rect 5254 1167 5272 1201
rect 5306 1167 5317 1201
rect 5254 1133 5317 1167
rect 5254 1099 5272 1133
rect 5306 1099 5317 1133
rect 5254 1065 5317 1099
rect 5254 1031 5272 1065
rect 5306 1031 5317 1065
rect 5254 997 5317 1031
rect 5254 963 5272 997
rect 5306 963 5317 997
rect 5254 929 5317 963
rect 5254 895 5272 929
rect 5306 895 5317 929
rect 5254 861 5317 895
rect 5254 827 5272 861
rect 5306 827 5317 861
rect 5254 793 5317 827
rect 5254 759 5272 793
rect 5306 759 5317 793
rect 5254 725 5317 759
rect 5254 691 5272 725
rect 5306 691 5317 725
rect 5254 657 5317 691
rect 5254 623 5272 657
rect 5306 623 5317 657
rect 5254 589 5317 623
rect 5254 555 5272 589
rect 5306 555 5317 589
rect 5254 521 5317 555
rect 5254 487 5272 521
rect 5306 487 5317 521
rect 5254 475 5317 487
rect 5384 1813 5447 1875
rect 5384 1779 5395 1813
rect 5429 1779 5447 1813
rect 5384 1745 5447 1779
rect 5384 1711 5395 1745
rect 5429 1711 5447 1745
rect 5384 1677 5447 1711
rect 5384 1643 5395 1677
rect 5429 1643 5447 1677
rect 5384 1609 5447 1643
rect 5384 1575 5395 1609
rect 5429 1575 5447 1609
rect 5384 1541 5447 1575
rect 5384 1507 5395 1541
rect 5429 1507 5447 1541
rect 5384 1473 5447 1507
rect 5384 1439 5395 1473
rect 5429 1439 5447 1473
rect 5384 1405 5447 1439
rect 5384 1371 5395 1405
rect 5429 1371 5447 1405
rect 5384 1337 5447 1371
rect 5384 1303 5395 1337
rect 5429 1303 5447 1337
rect 5384 1269 5447 1303
rect 5384 1235 5395 1269
rect 5429 1235 5447 1269
rect 5384 1201 5447 1235
rect 5384 1167 5395 1201
rect 5429 1167 5447 1201
rect 5384 1133 5447 1167
rect 5384 1099 5395 1133
rect 5429 1099 5447 1133
rect 5384 1065 5447 1099
rect 5384 1031 5395 1065
rect 5429 1031 5447 1065
rect 5384 997 5447 1031
rect 5384 963 5395 997
rect 5429 963 5447 997
rect 5384 929 5447 963
rect 5384 895 5395 929
rect 5429 895 5447 929
rect 5384 861 5447 895
rect 5384 827 5395 861
rect 5429 827 5447 861
rect 5384 793 5447 827
rect 5384 759 5395 793
rect 5429 759 5447 793
rect 5384 725 5447 759
rect 5384 691 5395 725
rect 5429 691 5447 725
rect 5384 657 5447 691
rect 5384 623 5395 657
rect 5429 623 5447 657
rect 5384 589 5447 623
rect 5384 555 5395 589
rect 5429 555 5447 589
rect 5384 521 5447 555
rect 5384 487 5395 521
rect 5429 487 5447 521
rect 5384 475 5447 487
rect 5547 1813 5603 1875
rect 5547 1779 5558 1813
rect 5592 1779 5603 1813
rect 5547 1745 5603 1779
rect 5547 1711 5558 1745
rect 5592 1711 5603 1745
rect 5547 1677 5603 1711
rect 5547 1643 5558 1677
rect 5592 1643 5603 1677
rect 5547 1609 5603 1643
rect 5547 1575 5558 1609
rect 5592 1575 5603 1609
rect 5547 1541 5603 1575
rect 5547 1507 5558 1541
rect 5592 1507 5603 1541
rect 5547 1473 5603 1507
rect 5547 1439 5558 1473
rect 5592 1439 5603 1473
rect 5547 1405 5603 1439
rect 5547 1371 5558 1405
rect 5592 1371 5603 1405
rect 5547 1337 5603 1371
rect 5547 1303 5558 1337
rect 5592 1303 5603 1337
rect 5547 1269 5603 1303
rect 5547 1235 5558 1269
rect 5592 1235 5603 1269
rect 5547 1201 5603 1235
rect 5547 1167 5558 1201
rect 5592 1167 5603 1201
rect 5547 1133 5603 1167
rect 5547 1099 5558 1133
rect 5592 1099 5603 1133
rect 5547 1065 5603 1099
rect 5547 1031 5558 1065
rect 5592 1031 5603 1065
rect 5547 997 5603 1031
rect 5547 963 5558 997
rect 5592 963 5603 997
rect 5547 929 5603 963
rect 5547 895 5558 929
rect 5592 895 5603 929
rect 5547 861 5603 895
rect 5547 827 5558 861
rect 5592 827 5603 861
rect 5547 793 5603 827
rect 5547 759 5558 793
rect 5592 759 5603 793
rect 5547 725 5603 759
rect 5547 691 5558 725
rect 5592 691 5603 725
rect 5547 657 5603 691
rect 5547 623 5558 657
rect 5592 623 5603 657
rect 5547 589 5603 623
rect 5547 555 5558 589
rect 5592 555 5603 589
rect 5547 521 5603 555
rect 5547 487 5558 521
rect 5592 487 5603 521
rect 5547 475 5603 487
rect 5703 1813 5773 1875
rect 5703 1779 5721 1813
rect 5755 1779 5773 1813
rect 5703 1745 5773 1779
rect 5703 1711 5721 1745
rect 5755 1711 5773 1745
rect 5703 1677 5773 1711
rect 5703 1643 5721 1677
rect 5755 1643 5773 1677
rect 5703 1609 5773 1643
rect 5703 1575 5721 1609
rect 5755 1575 5773 1609
rect 5703 1541 5773 1575
rect 5703 1507 5721 1541
rect 5755 1507 5773 1541
rect 5703 1473 5773 1507
rect 5703 1439 5721 1473
rect 5755 1439 5773 1473
rect 5703 1405 5773 1439
rect 5703 1371 5721 1405
rect 5755 1371 5773 1405
rect 5703 1337 5773 1371
rect 5703 1303 5721 1337
rect 5755 1303 5773 1337
rect 5703 1269 5773 1303
rect 5703 1235 5721 1269
rect 5755 1235 5773 1269
rect 5703 1201 5773 1235
rect 5703 1167 5721 1201
rect 5755 1167 5773 1201
rect 5703 1133 5773 1167
rect 5703 1099 5721 1133
rect 5755 1099 5773 1133
rect 5703 1065 5773 1099
rect 5703 1031 5721 1065
rect 5755 1031 5773 1065
rect 5703 997 5773 1031
rect 5703 963 5721 997
rect 5755 963 5773 997
rect 5703 929 5773 963
rect 5703 895 5721 929
rect 5755 895 5773 929
rect 5703 861 5773 895
rect 5703 827 5721 861
rect 5755 827 5773 861
rect 5703 793 5773 827
rect 5703 759 5721 793
rect 5755 759 5773 793
rect 5703 725 5773 759
rect 5703 691 5721 725
rect 5755 691 5773 725
rect 5703 657 5773 691
rect 5703 623 5721 657
rect 5755 623 5773 657
rect 5703 589 5773 623
rect 5703 555 5721 589
rect 5755 555 5773 589
rect 5703 521 5773 555
rect 5703 487 5721 521
rect 5755 487 5773 521
rect 5703 475 5773 487
rect 5873 1813 5929 1875
rect 5873 1779 5884 1813
rect 5918 1779 5929 1813
rect 5873 1745 5929 1779
rect 5873 1711 5884 1745
rect 5918 1711 5929 1745
rect 5873 1677 5929 1711
rect 5873 1643 5884 1677
rect 5918 1643 5929 1677
rect 5873 1609 5929 1643
rect 5873 1575 5884 1609
rect 5918 1575 5929 1609
rect 5873 1541 5929 1575
rect 5873 1507 5884 1541
rect 5918 1507 5929 1541
rect 5873 1473 5929 1507
rect 5873 1439 5884 1473
rect 5918 1439 5929 1473
rect 5873 1405 5929 1439
rect 5873 1371 5884 1405
rect 5918 1371 5929 1405
rect 5873 1337 5929 1371
rect 5873 1303 5884 1337
rect 5918 1303 5929 1337
rect 5873 1269 5929 1303
rect 5873 1235 5884 1269
rect 5918 1235 5929 1269
rect 5873 1201 5929 1235
rect 5873 1167 5884 1201
rect 5918 1167 5929 1201
rect 5873 1133 5929 1167
rect 5873 1099 5884 1133
rect 5918 1099 5929 1133
rect 5873 1065 5929 1099
rect 5873 1031 5884 1065
rect 5918 1031 5929 1065
rect 5873 997 5929 1031
rect 5873 963 5884 997
rect 5918 963 5929 997
rect 5873 929 5929 963
rect 5873 895 5884 929
rect 5918 895 5929 929
rect 5873 861 5929 895
rect 5873 827 5884 861
rect 5918 827 5929 861
rect 5873 793 5929 827
rect 5873 759 5884 793
rect 5918 759 5929 793
rect 5873 725 5929 759
rect 5873 691 5884 725
rect 5918 691 5929 725
rect 5873 657 5929 691
rect 5873 623 5884 657
rect 5918 623 5929 657
rect 5873 589 5929 623
rect 5873 555 5884 589
rect 5918 555 5929 589
rect 5873 521 5929 555
rect 5873 487 5884 521
rect 5918 487 5929 521
rect 5873 475 5929 487
rect 6029 1813 6099 1875
rect 6029 1779 6047 1813
rect 6081 1779 6099 1813
rect 6029 1745 6099 1779
rect 6029 1711 6047 1745
rect 6081 1711 6099 1745
rect 6029 1677 6099 1711
rect 6029 1643 6047 1677
rect 6081 1643 6099 1677
rect 6029 1609 6099 1643
rect 6029 1575 6047 1609
rect 6081 1575 6099 1609
rect 6029 1541 6099 1575
rect 6029 1507 6047 1541
rect 6081 1507 6099 1541
rect 6029 1473 6099 1507
rect 6029 1439 6047 1473
rect 6081 1439 6099 1473
rect 6029 1405 6099 1439
rect 6029 1371 6047 1405
rect 6081 1371 6099 1405
rect 6029 1337 6099 1371
rect 6029 1303 6047 1337
rect 6081 1303 6099 1337
rect 6029 1269 6099 1303
rect 6029 1235 6047 1269
rect 6081 1235 6099 1269
rect 6029 1201 6099 1235
rect 6029 1167 6047 1201
rect 6081 1167 6099 1201
rect 6029 1133 6099 1167
rect 6029 1099 6047 1133
rect 6081 1099 6099 1133
rect 6029 1065 6099 1099
rect 6029 1031 6047 1065
rect 6081 1031 6099 1065
rect 6029 997 6099 1031
rect 6029 963 6047 997
rect 6081 963 6099 997
rect 6029 929 6099 963
rect 6029 895 6047 929
rect 6081 895 6099 929
rect 6029 861 6099 895
rect 6029 827 6047 861
rect 6081 827 6099 861
rect 6029 793 6099 827
rect 6029 759 6047 793
rect 6081 759 6099 793
rect 6029 725 6099 759
rect 6029 691 6047 725
rect 6081 691 6099 725
rect 6029 657 6099 691
rect 6029 623 6047 657
rect 6081 623 6099 657
rect 6029 589 6099 623
rect 6029 555 6047 589
rect 6081 555 6099 589
rect 6029 521 6099 555
rect 6029 487 6047 521
rect 6081 487 6099 521
rect 6029 475 6099 487
rect 6199 1813 6255 1875
rect 6199 1779 6210 1813
rect 6244 1779 6255 1813
rect 6199 1745 6255 1779
rect 6199 1711 6210 1745
rect 6244 1711 6255 1745
rect 6199 1677 6255 1711
rect 6199 1643 6210 1677
rect 6244 1643 6255 1677
rect 6199 1609 6255 1643
rect 6199 1575 6210 1609
rect 6244 1575 6255 1609
rect 6199 1541 6255 1575
rect 6199 1507 6210 1541
rect 6244 1507 6255 1541
rect 6199 1473 6255 1507
rect 6199 1439 6210 1473
rect 6244 1439 6255 1473
rect 6199 1405 6255 1439
rect 6199 1371 6210 1405
rect 6244 1371 6255 1405
rect 6199 1337 6255 1371
rect 6199 1303 6210 1337
rect 6244 1303 6255 1337
rect 6199 1269 6255 1303
rect 6199 1235 6210 1269
rect 6244 1235 6255 1269
rect 6199 1201 6255 1235
rect 6199 1167 6210 1201
rect 6244 1167 6255 1201
rect 6199 1133 6255 1167
rect 6199 1099 6210 1133
rect 6244 1099 6255 1133
rect 6199 1065 6255 1099
rect 6199 1031 6210 1065
rect 6244 1031 6255 1065
rect 6199 997 6255 1031
rect 6199 963 6210 997
rect 6244 963 6255 997
rect 6199 929 6255 963
rect 6199 895 6210 929
rect 6244 895 6255 929
rect 6199 861 6255 895
rect 6199 827 6210 861
rect 6244 827 6255 861
rect 6199 793 6255 827
rect 6199 759 6210 793
rect 6244 759 6255 793
rect 6199 725 6255 759
rect 6199 691 6210 725
rect 6244 691 6255 725
rect 6199 657 6255 691
rect 6199 623 6210 657
rect 6244 623 6255 657
rect 6199 589 6255 623
rect 6199 555 6210 589
rect 6244 555 6255 589
rect 6199 521 6255 555
rect 6199 487 6210 521
rect 6244 487 6255 521
rect 6199 475 6255 487
rect 6355 1813 6425 1875
rect 6355 1779 6373 1813
rect 6407 1779 6425 1813
rect 6355 1745 6425 1779
rect 6355 1711 6373 1745
rect 6407 1711 6425 1745
rect 6355 1677 6425 1711
rect 6355 1643 6373 1677
rect 6407 1643 6425 1677
rect 6355 1609 6425 1643
rect 6355 1575 6373 1609
rect 6407 1575 6425 1609
rect 6355 1541 6425 1575
rect 6355 1507 6373 1541
rect 6407 1507 6425 1541
rect 6355 1473 6425 1507
rect 6355 1439 6373 1473
rect 6407 1439 6425 1473
rect 6355 1405 6425 1439
rect 6355 1371 6373 1405
rect 6407 1371 6425 1405
rect 6355 1337 6425 1371
rect 6355 1303 6373 1337
rect 6407 1303 6425 1337
rect 6355 1269 6425 1303
rect 6355 1235 6373 1269
rect 6407 1235 6425 1269
rect 6355 1201 6425 1235
rect 6355 1167 6373 1201
rect 6407 1167 6425 1201
rect 6355 1133 6425 1167
rect 6355 1099 6373 1133
rect 6407 1099 6425 1133
rect 6355 1065 6425 1099
rect 6355 1031 6373 1065
rect 6407 1031 6425 1065
rect 6355 997 6425 1031
rect 6355 963 6373 997
rect 6407 963 6425 997
rect 6355 929 6425 963
rect 6355 895 6373 929
rect 6407 895 6425 929
rect 6355 861 6425 895
rect 6355 827 6373 861
rect 6407 827 6425 861
rect 6355 793 6425 827
rect 6355 759 6373 793
rect 6407 759 6425 793
rect 6355 725 6425 759
rect 6355 691 6373 725
rect 6407 691 6425 725
rect 6355 657 6425 691
rect 6355 623 6373 657
rect 6407 623 6425 657
rect 6355 589 6425 623
rect 6355 555 6373 589
rect 6407 555 6425 589
rect 6355 521 6425 555
rect 6355 487 6373 521
rect 6407 487 6425 521
rect 6355 475 6425 487
rect 6525 1813 6581 1875
rect 6525 1779 6536 1813
rect 6570 1779 6581 1813
rect 6525 1745 6581 1779
rect 6525 1711 6536 1745
rect 6570 1711 6581 1745
rect 6525 1677 6581 1711
rect 6525 1643 6536 1677
rect 6570 1643 6581 1677
rect 6525 1609 6581 1643
rect 6525 1575 6536 1609
rect 6570 1575 6581 1609
rect 6525 1541 6581 1575
rect 6525 1507 6536 1541
rect 6570 1507 6581 1541
rect 6525 1473 6581 1507
rect 6525 1439 6536 1473
rect 6570 1439 6581 1473
rect 6525 1405 6581 1439
rect 6525 1371 6536 1405
rect 6570 1371 6581 1405
rect 6525 1337 6581 1371
rect 6525 1303 6536 1337
rect 6570 1303 6581 1337
rect 6525 1269 6581 1303
rect 6525 1235 6536 1269
rect 6570 1235 6581 1269
rect 6525 1201 6581 1235
rect 6525 1167 6536 1201
rect 6570 1167 6581 1201
rect 6525 1133 6581 1167
rect 6525 1099 6536 1133
rect 6570 1099 6581 1133
rect 6525 1065 6581 1099
rect 6525 1031 6536 1065
rect 6570 1031 6581 1065
rect 6525 997 6581 1031
rect 6525 963 6536 997
rect 6570 963 6581 997
rect 6525 929 6581 963
rect 6525 895 6536 929
rect 6570 895 6581 929
rect 6525 861 6581 895
rect 6525 827 6536 861
rect 6570 827 6581 861
rect 6525 793 6581 827
rect 6525 759 6536 793
rect 6570 759 6581 793
rect 6525 725 6581 759
rect 6525 691 6536 725
rect 6570 691 6581 725
rect 6525 657 6581 691
rect 6525 623 6536 657
rect 6570 623 6581 657
rect 6525 589 6581 623
rect 6525 555 6536 589
rect 6570 555 6581 589
rect 6525 521 6581 555
rect 6525 487 6536 521
rect 6570 487 6581 521
rect 6525 475 6581 487
rect 7205 1881 7261 1943
rect 7205 1847 7216 1881
rect 7250 1847 7261 1881
rect 7205 1813 7261 1847
rect 7205 1779 7216 1813
rect 7250 1779 7261 1813
rect 7205 1745 7261 1779
rect 7205 1711 7216 1745
rect 7250 1711 7261 1745
rect 7205 1677 7261 1711
rect 7205 1643 7216 1677
rect 7250 1643 7261 1677
rect 7205 1609 7261 1643
rect 7205 1575 7216 1609
rect 7250 1575 7261 1609
rect 7205 1541 7261 1575
rect 7205 1507 7216 1541
rect 7250 1507 7261 1541
rect 7205 1473 7261 1507
rect 7205 1439 7216 1473
rect 7250 1439 7261 1473
rect 7205 1405 7261 1439
rect 7205 1371 7216 1405
rect 7250 1371 7261 1405
rect 7205 1337 7261 1371
rect 7205 1303 7216 1337
rect 7250 1303 7261 1337
rect 7205 1269 7261 1303
rect 7205 1235 7216 1269
rect 7250 1235 7261 1269
rect 7205 1201 7261 1235
rect 7205 1167 7216 1201
rect 7250 1167 7261 1201
rect 7205 1133 7261 1167
rect 7205 1099 7216 1133
rect 7250 1099 7261 1133
rect 7205 1065 7261 1099
rect 7205 1031 7216 1065
rect 7250 1031 7261 1065
rect 7205 997 7261 1031
rect 7205 963 7216 997
rect 7250 963 7261 997
rect 7205 929 7261 963
rect 7205 895 7216 929
rect 7250 895 7261 929
rect 7205 861 7261 895
rect 7205 827 7216 861
rect 7250 827 7261 861
rect 7205 793 7261 827
rect 7205 759 7216 793
rect 7250 759 7261 793
rect 7205 725 7261 759
rect 7205 691 7216 725
rect 7250 691 7261 725
rect 7205 657 7261 691
rect 7205 623 7216 657
rect 7250 623 7261 657
rect 7205 589 7261 623
rect 7205 555 7216 589
rect 7250 555 7261 589
rect 7205 543 7261 555
rect 7361 1881 7431 1943
rect 7361 1847 7379 1881
rect 7413 1847 7431 1881
rect 7361 1813 7431 1847
rect 7361 1779 7379 1813
rect 7413 1779 7431 1813
rect 7361 1745 7431 1779
rect 7361 1711 7379 1745
rect 7413 1711 7431 1745
rect 7361 1677 7431 1711
rect 7361 1643 7379 1677
rect 7413 1643 7431 1677
rect 7361 1609 7431 1643
rect 7361 1575 7379 1609
rect 7413 1575 7431 1609
rect 7361 1541 7431 1575
rect 7361 1507 7379 1541
rect 7413 1507 7431 1541
rect 7361 1473 7431 1507
rect 7361 1439 7379 1473
rect 7413 1439 7431 1473
rect 7361 1405 7431 1439
rect 7361 1371 7379 1405
rect 7413 1371 7431 1405
rect 7361 1337 7431 1371
rect 7361 1303 7379 1337
rect 7413 1303 7431 1337
rect 7361 1269 7431 1303
rect 7361 1235 7379 1269
rect 7413 1235 7431 1269
rect 7361 1201 7431 1235
rect 7361 1167 7379 1201
rect 7413 1167 7431 1201
rect 7361 1133 7431 1167
rect 7361 1099 7379 1133
rect 7413 1099 7431 1133
rect 7361 1065 7431 1099
rect 7361 1031 7379 1065
rect 7413 1031 7431 1065
rect 7361 997 7431 1031
rect 7361 963 7379 997
rect 7413 963 7431 997
rect 7361 929 7431 963
rect 7361 895 7379 929
rect 7413 895 7431 929
rect 7361 861 7431 895
rect 7361 827 7379 861
rect 7413 827 7431 861
rect 7361 793 7431 827
rect 7361 759 7379 793
rect 7413 759 7431 793
rect 7361 725 7431 759
rect 7361 691 7379 725
rect 7413 691 7431 725
rect 7361 657 7431 691
rect 7361 623 7379 657
rect 7413 623 7431 657
rect 7361 589 7431 623
rect 7361 555 7379 589
rect 7413 555 7431 589
rect 7361 543 7431 555
rect 7531 1881 7587 1943
rect 7531 1847 7542 1881
rect 7576 1847 7587 1881
rect 7531 1813 7587 1847
rect 7531 1779 7542 1813
rect 7576 1779 7587 1813
rect 7531 1745 7587 1779
rect 7531 1711 7542 1745
rect 7576 1711 7587 1745
rect 7531 1677 7587 1711
rect 7531 1643 7542 1677
rect 7576 1643 7587 1677
rect 7531 1609 7587 1643
rect 7531 1575 7542 1609
rect 7576 1575 7587 1609
rect 7531 1541 7587 1575
rect 7531 1507 7542 1541
rect 7576 1507 7587 1541
rect 7531 1473 7587 1507
rect 7531 1439 7542 1473
rect 7576 1439 7587 1473
rect 7531 1405 7587 1439
rect 7531 1371 7542 1405
rect 7576 1371 7587 1405
rect 7531 1337 7587 1371
rect 7531 1303 7542 1337
rect 7576 1303 7587 1337
rect 7531 1269 7587 1303
rect 7531 1235 7542 1269
rect 7576 1235 7587 1269
rect 7531 1201 7587 1235
rect 7531 1167 7542 1201
rect 7576 1167 7587 1201
rect 7531 1133 7587 1167
rect 7531 1099 7542 1133
rect 7576 1099 7587 1133
rect 7531 1065 7587 1099
rect 7531 1031 7542 1065
rect 7576 1031 7587 1065
rect 7531 997 7587 1031
rect 7531 963 7542 997
rect 7576 963 7587 997
rect 7531 929 7587 963
rect 7531 895 7542 929
rect 7576 895 7587 929
rect 7531 861 7587 895
rect 7531 827 7542 861
rect 7576 827 7587 861
rect 7531 793 7587 827
rect 7531 759 7542 793
rect 7576 759 7587 793
rect 7531 725 7587 759
rect 7531 691 7542 725
rect 7576 691 7587 725
rect 7531 657 7587 691
rect 7531 623 7542 657
rect 7576 623 7587 657
rect 7531 589 7587 623
rect 7531 555 7542 589
rect 7576 555 7587 589
rect 7531 543 7587 555
rect 7687 1881 7757 1943
rect 7687 1847 7705 1881
rect 7739 1847 7757 1881
rect 7687 1813 7757 1847
rect 7687 1779 7705 1813
rect 7739 1779 7757 1813
rect 7687 1745 7757 1779
rect 7687 1711 7705 1745
rect 7739 1711 7757 1745
rect 7687 1677 7757 1711
rect 7687 1643 7705 1677
rect 7739 1643 7757 1677
rect 7687 1609 7757 1643
rect 7687 1575 7705 1609
rect 7739 1575 7757 1609
rect 7687 1541 7757 1575
rect 7687 1507 7705 1541
rect 7739 1507 7757 1541
rect 7687 1473 7757 1507
rect 7687 1439 7705 1473
rect 7739 1439 7757 1473
rect 7687 1405 7757 1439
rect 7687 1371 7705 1405
rect 7739 1371 7757 1405
rect 7687 1337 7757 1371
rect 7687 1303 7705 1337
rect 7739 1303 7757 1337
rect 7687 1269 7757 1303
rect 7687 1235 7705 1269
rect 7739 1235 7757 1269
rect 7687 1201 7757 1235
rect 7687 1167 7705 1201
rect 7739 1167 7757 1201
rect 7687 1133 7757 1167
rect 7687 1099 7705 1133
rect 7739 1099 7757 1133
rect 7687 1065 7757 1099
rect 7687 1031 7705 1065
rect 7739 1031 7757 1065
rect 7687 997 7757 1031
rect 7687 963 7705 997
rect 7739 963 7757 997
rect 7687 929 7757 963
rect 7687 895 7705 929
rect 7739 895 7757 929
rect 7687 861 7757 895
rect 7687 827 7705 861
rect 7739 827 7757 861
rect 7687 793 7757 827
rect 7687 759 7705 793
rect 7739 759 7757 793
rect 7687 725 7757 759
rect 7687 691 7705 725
rect 7739 691 7757 725
rect 7687 657 7757 691
rect 7687 623 7705 657
rect 7739 623 7757 657
rect 7687 589 7757 623
rect 7687 555 7705 589
rect 7739 555 7757 589
rect 7687 543 7757 555
rect 7857 1881 7913 1943
rect 7857 1847 7868 1881
rect 7902 1847 7913 1881
rect 7857 1813 7913 1847
rect 7857 1779 7868 1813
rect 7902 1779 7913 1813
rect 7857 1745 7913 1779
rect 7857 1711 7868 1745
rect 7902 1711 7913 1745
rect 7857 1677 7913 1711
rect 7857 1643 7868 1677
rect 7902 1643 7913 1677
rect 7857 1609 7913 1643
rect 7857 1575 7868 1609
rect 7902 1575 7913 1609
rect 7857 1541 7913 1575
rect 7857 1507 7868 1541
rect 7902 1507 7913 1541
rect 7857 1473 7913 1507
rect 7857 1439 7868 1473
rect 7902 1439 7913 1473
rect 7857 1405 7913 1439
rect 7857 1371 7868 1405
rect 7902 1371 7913 1405
rect 7857 1337 7913 1371
rect 7857 1303 7868 1337
rect 7902 1303 7913 1337
rect 7857 1269 7913 1303
rect 7857 1235 7868 1269
rect 7902 1235 7913 1269
rect 7857 1201 7913 1235
rect 7857 1167 7868 1201
rect 7902 1167 7913 1201
rect 7857 1133 7913 1167
rect 7857 1099 7868 1133
rect 7902 1099 7913 1133
rect 7857 1065 7913 1099
rect 7857 1031 7868 1065
rect 7902 1031 7913 1065
rect 7857 997 7913 1031
rect 7857 963 7868 997
rect 7902 963 7913 997
rect 7857 929 7913 963
rect 7857 895 7868 929
rect 7902 895 7913 929
rect 7857 861 7913 895
rect 7857 827 7868 861
rect 7902 827 7913 861
rect 7857 793 7913 827
rect 7857 759 7868 793
rect 7902 759 7913 793
rect 7857 725 7913 759
rect 7857 691 7868 725
rect 7902 691 7913 725
rect 7857 657 7913 691
rect 7857 623 7868 657
rect 7902 623 7913 657
rect 7857 589 7913 623
rect 7857 555 7868 589
rect 7902 555 7913 589
rect 7857 543 7913 555
rect 8013 1881 8083 1943
rect 8013 1847 8031 1881
rect 8065 1847 8083 1881
rect 8013 1813 8083 1847
rect 8013 1779 8031 1813
rect 8065 1779 8083 1813
rect 8013 1745 8083 1779
rect 8013 1711 8031 1745
rect 8065 1711 8083 1745
rect 8013 1677 8083 1711
rect 8013 1643 8031 1677
rect 8065 1643 8083 1677
rect 8013 1609 8083 1643
rect 8013 1575 8031 1609
rect 8065 1575 8083 1609
rect 8013 1541 8083 1575
rect 8013 1507 8031 1541
rect 8065 1507 8083 1541
rect 8013 1473 8083 1507
rect 8013 1439 8031 1473
rect 8065 1439 8083 1473
rect 8013 1405 8083 1439
rect 8013 1371 8031 1405
rect 8065 1371 8083 1405
rect 8013 1337 8083 1371
rect 8013 1303 8031 1337
rect 8065 1303 8083 1337
rect 8013 1269 8083 1303
rect 8013 1235 8031 1269
rect 8065 1235 8083 1269
rect 8013 1201 8083 1235
rect 8013 1167 8031 1201
rect 8065 1167 8083 1201
rect 8013 1133 8083 1167
rect 8013 1099 8031 1133
rect 8065 1099 8083 1133
rect 8013 1065 8083 1099
rect 8013 1031 8031 1065
rect 8065 1031 8083 1065
rect 8013 997 8083 1031
rect 8013 963 8031 997
rect 8065 963 8083 997
rect 8013 929 8083 963
rect 8013 895 8031 929
rect 8065 895 8083 929
rect 8013 861 8083 895
rect 8013 827 8031 861
rect 8065 827 8083 861
rect 8013 793 8083 827
rect 8013 759 8031 793
rect 8065 759 8083 793
rect 8013 725 8083 759
rect 8013 691 8031 725
rect 8065 691 8083 725
rect 8013 657 8083 691
rect 8013 623 8031 657
rect 8065 623 8083 657
rect 8013 589 8083 623
rect 8013 555 8031 589
rect 8065 555 8083 589
rect 8013 543 8083 555
rect 8183 1881 8239 1943
rect 8183 1847 8194 1881
rect 8228 1847 8239 1881
rect 8183 1813 8239 1847
rect 8183 1779 8194 1813
rect 8228 1779 8239 1813
rect 8183 1745 8239 1779
rect 8183 1711 8194 1745
rect 8228 1711 8239 1745
rect 8183 1677 8239 1711
rect 8183 1643 8194 1677
rect 8228 1643 8239 1677
rect 8183 1609 8239 1643
rect 8183 1575 8194 1609
rect 8228 1575 8239 1609
rect 8183 1541 8239 1575
rect 8183 1507 8194 1541
rect 8228 1507 8239 1541
rect 8183 1473 8239 1507
rect 8183 1439 8194 1473
rect 8228 1439 8239 1473
rect 8183 1405 8239 1439
rect 8183 1371 8194 1405
rect 8228 1371 8239 1405
rect 8183 1337 8239 1371
rect 8183 1303 8194 1337
rect 8228 1303 8239 1337
rect 8183 1269 8239 1303
rect 8183 1235 8194 1269
rect 8228 1235 8239 1269
rect 8183 1201 8239 1235
rect 8183 1167 8194 1201
rect 8228 1167 8239 1201
rect 8183 1133 8239 1167
rect 8183 1099 8194 1133
rect 8228 1099 8239 1133
rect 8183 1065 8239 1099
rect 8183 1031 8194 1065
rect 8228 1031 8239 1065
rect 8183 997 8239 1031
rect 8183 963 8194 997
rect 8228 963 8239 997
rect 8183 929 8239 963
rect 8183 895 8194 929
rect 8228 895 8239 929
rect 8183 861 8239 895
rect 8183 827 8194 861
rect 8228 827 8239 861
rect 8183 793 8239 827
rect 8183 759 8194 793
rect 8228 759 8239 793
rect 8183 725 8239 759
rect 8183 691 8194 725
rect 8228 691 8239 725
rect 8183 657 8239 691
rect 8183 623 8194 657
rect 8228 623 8239 657
rect 8183 589 8239 623
rect 8183 555 8194 589
rect 8228 555 8239 589
rect 8183 543 8239 555
rect 8339 1881 8402 1943
rect 8339 1847 8357 1881
rect 8391 1847 8402 1881
rect 8339 1813 8402 1847
rect 8339 1779 8357 1813
rect 8391 1779 8402 1813
rect 8339 1745 8402 1779
rect 8339 1711 8357 1745
rect 8391 1711 8402 1745
rect 8339 1677 8402 1711
rect 8339 1643 8357 1677
rect 8391 1643 8402 1677
rect 8339 1609 8402 1643
rect 8339 1575 8357 1609
rect 8391 1575 8402 1609
rect 8339 1541 8402 1575
rect 8339 1507 8357 1541
rect 8391 1507 8402 1541
rect 8339 1473 8402 1507
rect 8339 1439 8357 1473
rect 8391 1439 8402 1473
rect 8339 1405 8402 1439
rect 8339 1371 8357 1405
rect 8391 1371 8402 1405
rect 8339 1337 8402 1371
rect 8339 1303 8357 1337
rect 8391 1303 8402 1337
rect 8339 1269 8402 1303
rect 8339 1235 8357 1269
rect 8391 1235 8402 1269
rect 8339 1201 8402 1235
rect 8339 1167 8357 1201
rect 8391 1167 8402 1201
rect 8339 1133 8402 1167
rect 8339 1099 8357 1133
rect 8391 1099 8402 1133
rect 8339 1065 8402 1099
rect 8339 1031 8357 1065
rect 8391 1031 8402 1065
rect 8339 997 8402 1031
rect 8339 963 8357 997
rect 8391 963 8402 997
rect 8339 929 8402 963
rect 8339 895 8357 929
rect 8391 895 8402 929
rect 8339 861 8402 895
rect 8339 827 8357 861
rect 8391 827 8402 861
rect 8339 793 8402 827
rect 8339 759 8357 793
rect 8391 759 8402 793
rect 8339 725 8402 759
rect 8339 691 8357 725
rect 8391 691 8402 725
rect 8339 657 8402 691
rect 8339 623 8357 657
rect 8391 623 8402 657
rect 8339 589 8402 623
rect 8339 555 8357 589
rect 8391 555 8402 589
rect 8339 543 8402 555
rect 8469 1881 8532 1943
rect 8469 1847 8480 1881
rect 8514 1847 8532 1881
rect 8469 1813 8532 1847
rect 8469 1779 8480 1813
rect 8514 1779 8532 1813
rect 8469 1745 8532 1779
rect 8469 1711 8480 1745
rect 8514 1711 8532 1745
rect 8469 1677 8532 1711
rect 8469 1643 8480 1677
rect 8514 1643 8532 1677
rect 8469 1609 8532 1643
rect 8469 1575 8480 1609
rect 8514 1575 8532 1609
rect 8469 1541 8532 1575
rect 8469 1507 8480 1541
rect 8514 1507 8532 1541
rect 8469 1473 8532 1507
rect 8469 1439 8480 1473
rect 8514 1439 8532 1473
rect 8469 1405 8532 1439
rect 8469 1371 8480 1405
rect 8514 1371 8532 1405
rect 8469 1337 8532 1371
rect 8469 1303 8480 1337
rect 8514 1303 8532 1337
rect 8469 1269 8532 1303
rect 8469 1235 8480 1269
rect 8514 1235 8532 1269
rect 8469 1201 8532 1235
rect 8469 1167 8480 1201
rect 8514 1167 8532 1201
rect 8469 1133 8532 1167
rect 8469 1099 8480 1133
rect 8514 1099 8532 1133
rect 8469 1065 8532 1099
rect 8469 1031 8480 1065
rect 8514 1031 8532 1065
rect 8469 997 8532 1031
rect 8469 963 8480 997
rect 8514 963 8532 997
rect 8469 929 8532 963
rect 8469 895 8480 929
rect 8514 895 8532 929
rect 8469 861 8532 895
rect 8469 827 8480 861
rect 8514 827 8532 861
rect 8469 793 8532 827
rect 8469 759 8480 793
rect 8514 759 8532 793
rect 8469 725 8532 759
rect 8469 691 8480 725
rect 8514 691 8532 725
rect 8469 657 8532 691
rect 8469 623 8480 657
rect 8514 623 8532 657
rect 8469 589 8532 623
rect 8469 555 8480 589
rect 8514 555 8532 589
rect 8469 543 8532 555
rect 8632 1881 8688 1943
rect 8632 1847 8643 1881
rect 8677 1847 8688 1881
rect 8632 1813 8688 1847
rect 8632 1779 8643 1813
rect 8677 1779 8688 1813
rect 8632 1745 8688 1779
rect 8632 1711 8643 1745
rect 8677 1711 8688 1745
rect 8632 1677 8688 1711
rect 8632 1643 8643 1677
rect 8677 1643 8688 1677
rect 8632 1609 8688 1643
rect 8632 1575 8643 1609
rect 8677 1575 8688 1609
rect 8632 1541 8688 1575
rect 8632 1507 8643 1541
rect 8677 1507 8688 1541
rect 8632 1473 8688 1507
rect 8632 1439 8643 1473
rect 8677 1439 8688 1473
rect 8632 1405 8688 1439
rect 8632 1371 8643 1405
rect 8677 1371 8688 1405
rect 8632 1337 8688 1371
rect 8632 1303 8643 1337
rect 8677 1303 8688 1337
rect 8632 1269 8688 1303
rect 8632 1235 8643 1269
rect 8677 1235 8688 1269
rect 8632 1201 8688 1235
rect 8632 1167 8643 1201
rect 8677 1167 8688 1201
rect 8632 1133 8688 1167
rect 8632 1099 8643 1133
rect 8677 1099 8688 1133
rect 8632 1065 8688 1099
rect 8632 1031 8643 1065
rect 8677 1031 8688 1065
rect 8632 997 8688 1031
rect 8632 963 8643 997
rect 8677 963 8688 997
rect 8632 929 8688 963
rect 8632 895 8643 929
rect 8677 895 8688 929
rect 8632 861 8688 895
rect 8632 827 8643 861
rect 8677 827 8688 861
rect 8632 793 8688 827
rect 8632 759 8643 793
rect 8677 759 8688 793
rect 8632 725 8688 759
rect 8632 691 8643 725
rect 8677 691 8688 725
rect 8632 657 8688 691
rect 8632 623 8643 657
rect 8677 623 8688 657
rect 8632 589 8688 623
rect 8632 555 8643 589
rect 8677 555 8688 589
rect 8632 543 8688 555
rect 8788 1881 8858 1943
rect 8788 1847 8806 1881
rect 8840 1847 8858 1881
rect 8788 1813 8858 1847
rect 8788 1779 8806 1813
rect 8840 1779 8858 1813
rect 8788 1745 8858 1779
rect 8788 1711 8806 1745
rect 8840 1711 8858 1745
rect 8788 1677 8858 1711
rect 8788 1643 8806 1677
rect 8840 1643 8858 1677
rect 8788 1609 8858 1643
rect 8788 1575 8806 1609
rect 8840 1575 8858 1609
rect 8788 1541 8858 1575
rect 8788 1507 8806 1541
rect 8840 1507 8858 1541
rect 8788 1473 8858 1507
rect 8788 1439 8806 1473
rect 8840 1439 8858 1473
rect 8788 1405 8858 1439
rect 8788 1371 8806 1405
rect 8840 1371 8858 1405
rect 8788 1337 8858 1371
rect 8788 1303 8806 1337
rect 8840 1303 8858 1337
rect 8788 1269 8858 1303
rect 8788 1235 8806 1269
rect 8840 1235 8858 1269
rect 8788 1201 8858 1235
rect 8788 1167 8806 1201
rect 8840 1167 8858 1201
rect 8788 1133 8858 1167
rect 8788 1099 8806 1133
rect 8840 1099 8858 1133
rect 8788 1065 8858 1099
rect 8788 1031 8806 1065
rect 8840 1031 8858 1065
rect 8788 997 8858 1031
rect 8788 963 8806 997
rect 8840 963 8858 997
rect 8788 929 8858 963
rect 8788 895 8806 929
rect 8840 895 8858 929
rect 8788 861 8858 895
rect 8788 827 8806 861
rect 8840 827 8858 861
rect 8788 793 8858 827
rect 8788 759 8806 793
rect 8840 759 8858 793
rect 8788 725 8858 759
rect 8788 691 8806 725
rect 8840 691 8858 725
rect 8788 657 8858 691
rect 8788 623 8806 657
rect 8840 623 8858 657
rect 8788 589 8858 623
rect 8788 555 8806 589
rect 8840 555 8858 589
rect 8788 543 8858 555
rect 8958 1881 9014 1943
rect 8958 1847 8969 1881
rect 9003 1847 9014 1881
rect 8958 1813 9014 1847
rect 8958 1779 8969 1813
rect 9003 1779 9014 1813
rect 8958 1745 9014 1779
rect 8958 1711 8969 1745
rect 9003 1711 9014 1745
rect 8958 1677 9014 1711
rect 8958 1643 8969 1677
rect 9003 1643 9014 1677
rect 8958 1609 9014 1643
rect 8958 1575 8969 1609
rect 9003 1575 9014 1609
rect 8958 1541 9014 1575
rect 8958 1507 8969 1541
rect 9003 1507 9014 1541
rect 8958 1473 9014 1507
rect 8958 1439 8969 1473
rect 9003 1439 9014 1473
rect 8958 1405 9014 1439
rect 8958 1371 8969 1405
rect 9003 1371 9014 1405
rect 8958 1337 9014 1371
rect 8958 1303 8969 1337
rect 9003 1303 9014 1337
rect 8958 1269 9014 1303
rect 8958 1235 8969 1269
rect 9003 1235 9014 1269
rect 8958 1201 9014 1235
rect 8958 1167 8969 1201
rect 9003 1167 9014 1201
rect 8958 1133 9014 1167
rect 8958 1099 8969 1133
rect 9003 1099 9014 1133
rect 8958 1065 9014 1099
rect 8958 1031 8969 1065
rect 9003 1031 9014 1065
rect 8958 997 9014 1031
rect 8958 963 8969 997
rect 9003 963 9014 997
rect 8958 929 9014 963
rect 8958 895 8969 929
rect 9003 895 9014 929
rect 8958 861 9014 895
rect 8958 827 8969 861
rect 9003 827 9014 861
rect 8958 793 9014 827
rect 8958 759 8969 793
rect 9003 759 9014 793
rect 8958 725 9014 759
rect 8958 691 8969 725
rect 9003 691 9014 725
rect 8958 657 9014 691
rect 8958 623 8969 657
rect 9003 623 9014 657
rect 8958 589 9014 623
rect 8958 555 8969 589
rect 9003 555 9014 589
rect 8958 543 9014 555
rect 9114 1881 9184 1943
rect 9114 1847 9132 1881
rect 9166 1847 9184 1881
rect 9114 1813 9184 1847
rect 9114 1779 9132 1813
rect 9166 1779 9184 1813
rect 9114 1745 9184 1779
rect 9114 1711 9132 1745
rect 9166 1711 9184 1745
rect 9114 1677 9184 1711
rect 9114 1643 9132 1677
rect 9166 1643 9184 1677
rect 9114 1609 9184 1643
rect 9114 1575 9132 1609
rect 9166 1575 9184 1609
rect 9114 1541 9184 1575
rect 9114 1507 9132 1541
rect 9166 1507 9184 1541
rect 9114 1473 9184 1507
rect 9114 1439 9132 1473
rect 9166 1439 9184 1473
rect 9114 1405 9184 1439
rect 9114 1371 9132 1405
rect 9166 1371 9184 1405
rect 9114 1337 9184 1371
rect 9114 1303 9132 1337
rect 9166 1303 9184 1337
rect 9114 1269 9184 1303
rect 9114 1235 9132 1269
rect 9166 1235 9184 1269
rect 9114 1201 9184 1235
rect 9114 1167 9132 1201
rect 9166 1167 9184 1201
rect 9114 1133 9184 1167
rect 9114 1099 9132 1133
rect 9166 1099 9184 1133
rect 9114 1065 9184 1099
rect 9114 1031 9132 1065
rect 9166 1031 9184 1065
rect 9114 997 9184 1031
rect 9114 963 9132 997
rect 9166 963 9184 997
rect 9114 929 9184 963
rect 9114 895 9132 929
rect 9166 895 9184 929
rect 9114 861 9184 895
rect 9114 827 9132 861
rect 9166 827 9184 861
rect 9114 793 9184 827
rect 9114 759 9132 793
rect 9166 759 9184 793
rect 9114 725 9184 759
rect 9114 691 9132 725
rect 9166 691 9184 725
rect 9114 657 9184 691
rect 9114 623 9132 657
rect 9166 623 9184 657
rect 9114 589 9184 623
rect 9114 555 9132 589
rect 9166 555 9184 589
rect 9114 543 9184 555
rect 9284 1881 9340 1943
rect 9284 1847 9295 1881
rect 9329 1847 9340 1881
rect 9284 1813 9340 1847
rect 9284 1779 9295 1813
rect 9329 1779 9340 1813
rect 9284 1745 9340 1779
rect 9284 1711 9295 1745
rect 9329 1711 9340 1745
rect 9284 1677 9340 1711
rect 9284 1643 9295 1677
rect 9329 1643 9340 1677
rect 9284 1609 9340 1643
rect 9284 1575 9295 1609
rect 9329 1575 9340 1609
rect 9284 1541 9340 1575
rect 9284 1507 9295 1541
rect 9329 1507 9340 1541
rect 9284 1473 9340 1507
rect 9284 1439 9295 1473
rect 9329 1439 9340 1473
rect 9284 1405 9340 1439
rect 9284 1371 9295 1405
rect 9329 1371 9340 1405
rect 9284 1337 9340 1371
rect 9284 1303 9295 1337
rect 9329 1303 9340 1337
rect 9284 1269 9340 1303
rect 9284 1235 9295 1269
rect 9329 1235 9340 1269
rect 9284 1201 9340 1235
rect 9284 1167 9295 1201
rect 9329 1167 9340 1201
rect 9284 1133 9340 1167
rect 9284 1099 9295 1133
rect 9329 1099 9340 1133
rect 9284 1065 9340 1099
rect 9284 1031 9295 1065
rect 9329 1031 9340 1065
rect 9284 997 9340 1031
rect 9284 963 9295 997
rect 9329 963 9340 997
rect 9284 929 9340 963
rect 9284 895 9295 929
rect 9329 895 9340 929
rect 9284 861 9340 895
rect 9284 827 9295 861
rect 9329 827 9340 861
rect 9284 793 9340 827
rect 9284 759 9295 793
rect 9329 759 9340 793
rect 9284 725 9340 759
rect 9284 691 9295 725
rect 9329 691 9340 725
rect 9284 657 9340 691
rect 9284 623 9295 657
rect 9329 623 9340 657
rect 9284 589 9340 623
rect 9284 555 9295 589
rect 9329 555 9340 589
rect 9284 543 9340 555
rect 9440 1881 9510 1943
rect 9440 1847 9458 1881
rect 9492 1847 9510 1881
rect 9440 1813 9510 1847
rect 9440 1779 9458 1813
rect 9492 1779 9510 1813
rect 9440 1745 9510 1779
rect 9440 1711 9458 1745
rect 9492 1711 9510 1745
rect 9440 1677 9510 1711
rect 9440 1643 9458 1677
rect 9492 1643 9510 1677
rect 9440 1609 9510 1643
rect 9440 1575 9458 1609
rect 9492 1575 9510 1609
rect 9440 1541 9510 1575
rect 9440 1507 9458 1541
rect 9492 1507 9510 1541
rect 9440 1473 9510 1507
rect 9440 1439 9458 1473
rect 9492 1439 9510 1473
rect 9440 1405 9510 1439
rect 9440 1371 9458 1405
rect 9492 1371 9510 1405
rect 9440 1337 9510 1371
rect 9440 1303 9458 1337
rect 9492 1303 9510 1337
rect 9440 1269 9510 1303
rect 9440 1235 9458 1269
rect 9492 1235 9510 1269
rect 9440 1201 9510 1235
rect 9440 1167 9458 1201
rect 9492 1167 9510 1201
rect 9440 1133 9510 1167
rect 9440 1099 9458 1133
rect 9492 1099 9510 1133
rect 9440 1065 9510 1099
rect 9440 1031 9458 1065
rect 9492 1031 9510 1065
rect 9440 997 9510 1031
rect 9440 963 9458 997
rect 9492 963 9510 997
rect 9440 929 9510 963
rect 9440 895 9458 929
rect 9492 895 9510 929
rect 9440 861 9510 895
rect 9440 827 9458 861
rect 9492 827 9510 861
rect 9440 793 9510 827
rect 9440 759 9458 793
rect 9492 759 9510 793
rect 9440 725 9510 759
rect 9440 691 9458 725
rect 9492 691 9510 725
rect 9440 657 9510 691
rect 9440 623 9458 657
rect 9492 623 9510 657
rect 9440 589 9510 623
rect 9440 555 9458 589
rect 9492 555 9510 589
rect 9440 543 9510 555
rect 9610 1881 9666 1943
rect 9610 1847 9621 1881
rect 9655 1847 9666 1881
rect 9610 1813 9666 1847
rect 9610 1779 9621 1813
rect 9655 1779 9666 1813
rect 9610 1745 9666 1779
rect 9610 1711 9621 1745
rect 9655 1711 9666 1745
rect 9610 1677 9666 1711
rect 9610 1643 9621 1677
rect 9655 1643 9666 1677
rect 9610 1609 9666 1643
rect 9610 1575 9621 1609
rect 9655 1575 9666 1609
rect 9610 1541 9666 1575
rect 9610 1507 9621 1541
rect 9655 1507 9666 1541
rect 9610 1473 9666 1507
rect 9610 1439 9621 1473
rect 9655 1439 9666 1473
rect 9610 1405 9666 1439
rect 9610 1371 9621 1405
rect 9655 1371 9666 1405
rect 9610 1337 9666 1371
rect 9610 1303 9621 1337
rect 9655 1303 9666 1337
rect 9610 1269 9666 1303
rect 9610 1235 9621 1269
rect 9655 1235 9666 1269
rect 9610 1201 9666 1235
rect 9610 1167 9621 1201
rect 9655 1167 9666 1201
rect 9610 1133 9666 1167
rect 9610 1099 9621 1133
rect 9655 1099 9666 1133
rect 9610 1065 9666 1099
rect 9610 1031 9621 1065
rect 9655 1031 9666 1065
rect 9610 997 9666 1031
rect 9610 963 9621 997
rect 9655 963 9666 997
rect 9610 929 9666 963
rect 9610 895 9621 929
rect 9655 895 9666 929
rect 9610 861 9666 895
rect 9610 827 9621 861
rect 9655 827 9666 861
rect 9610 793 9666 827
rect 9610 759 9621 793
rect 9655 759 9666 793
rect 9610 725 9666 759
rect 9610 691 9621 725
rect 9655 691 9666 725
rect 9610 657 9666 691
rect 9610 623 9621 657
rect 9655 623 9666 657
rect 9610 589 9666 623
rect 9610 555 9621 589
rect 9655 555 9666 589
rect 9610 543 9666 555
rect 9766 1881 9829 1943
rect 9766 1847 9784 1881
rect 9818 1847 9829 1881
rect 9766 1813 9829 1847
rect 9766 1779 9784 1813
rect 9818 1779 9829 1813
rect 9766 1745 9829 1779
rect 9766 1711 9784 1745
rect 9818 1711 9829 1745
rect 9766 1677 9829 1711
rect 9766 1643 9784 1677
rect 9818 1643 9829 1677
rect 9766 1609 9829 1643
rect 9766 1575 9784 1609
rect 9818 1575 9829 1609
rect 9766 1541 9829 1575
rect 9766 1507 9784 1541
rect 9818 1507 9829 1541
rect 9766 1473 9829 1507
rect 9766 1439 9784 1473
rect 9818 1439 9829 1473
rect 9766 1405 9829 1439
rect 9766 1371 9784 1405
rect 9818 1371 9829 1405
rect 9766 1337 9829 1371
rect 9766 1303 9784 1337
rect 9818 1303 9829 1337
rect 9766 1269 9829 1303
rect 9766 1235 9784 1269
rect 9818 1235 9829 1269
rect 9766 1201 9829 1235
rect 9766 1167 9784 1201
rect 9818 1167 9829 1201
rect 9766 1133 9829 1167
rect 9766 1099 9784 1133
rect 9818 1099 9829 1133
rect 9766 1065 9829 1099
rect 9766 1031 9784 1065
rect 9818 1031 9829 1065
rect 9766 997 9829 1031
rect 9766 963 9784 997
rect 9818 963 9829 997
rect 9766 929 9829 963
rect 9766 895 9784 929
rect 9818 895 9829 929
rect 9766 861 9829 895
rect 9766 827 9784 861
rect 9818 827 9829 861
rect 9766 793 9829 827
rect 9766 759 9784 793
rect 9818 759 9829 793
rect 9766 725 9829 759
rect 9766 691 9784 725
rect 9818 691 9829 725
rect 9766 657 9829 691
rect 9766 623 9784 657
rect 9818 623 9829 657
rect 9766 589 9829 623
rect 9766 555 9784 589
rect 9818 555 9829 589
rect 9766 543 9829 555
<< mvpdiff >>
rect 351 1813 414 1875
rect 351 1779 362 1813
rect 396 1779 414 1813
rect 351 1745 414 1779
rect 351 1711 362 1745
rect 396 1711 414 1745
rect 351 1677 414 1711
rect 351 1643 362 1677
rect 396 1643 414 1677
rect 351 1609 414 1643
rect 351 1575 362 1609
rect 396 1575 414 1609
rect 351 1541 414 1575
rect 351 1507 362 1541
rect 396 1507 414 1541
rect 351 1473 414 1507
rect 351 1439 362 1473
rect 396 1439 414 1473
rect 351 1405 414 1439
rect 351 1371 362 1405
rect 396 1371 414 1405
rect 351 1337 414 1371
rect 351 1303 362 1337
rect 396 1303 414 1337
rect 351 1269 414 1303
rect 351 1235 362 1269
rect 396 1235 414 1269
rect 351 1201 414 1235
rect 351 1167 362 1201
rect 396 1167 414 1201
rect 351 1133 414 1167
rect 351 1099 362 1133
rect 396 1099 414 1133
rect 351 1065 414 1099
rect 351 1031 362 1065
rect 396 1031 414 1065
rect 351 997 414 1031
rect 351 963 362 997
rect 396 963 414 997
rect 351 929 414 963
rect 351 895 362 929
rect 396 895 414 929
rect 351 861 414 895
rect 351 827 362 861
rect 396 827 414 861
rect 351 793 414 827
rect 351 759 362 793
rect 396 759 414 793
rect 351 725 414 759
rect 351 691 362 725
rect 396 691 414 725
rect 351 657 414 691
rect 351 623 362 657
rect 396 623 414 657
rect 351 589 414 623
rect 351 555 362 589
rect 396 555 414 589
rect 351 521 414 555
rect 351 487 362 521
rect 396 487 414 521
rect 351 475 414 487
rect 514 1813 570 1875
rect 514 1779 525 1813
rect 559 1779 570 1813
rect 514 1745 570 1779
rect 514 1711 525 1745
rect 559 1711 570 1745
rect 514 1677 570 1711
rect 514 1643 525 1677
rect 559 1643 570 1677
rect 514 1609 570 1643
rect 514 1575 525 1609
rect 559 1575 570 1609
rect 514 1541 570 1575
rect 514 1507 525 1541
rect 559 1507 570 1541
rect 514 1473 570 1507
rect 514 1439 525 1473
rect 559 1439 570 1473
rect 514 1405 570 1439
rect 514 1371 525 1405
rect 559 1371 570 1405
rect 514 1337 570 1371
rect 514 1303 525 1337
rect 559 1303 570 1337
rect 514 1269 570 1303
rect 514 1235 525 1269
rect 559 1235 570 1269
rect 514 1201 570 1235
rect 514 1167 525 1201
rect 559 1167 570 1201
rect 514 1133 570 1167
rect 514 1099 525 1133
rect 559 1099 570 1133
rect 514 1065 570 1099
rect 514 1031 525 1065
rect 559 1031 570 1065
rect 514 997 570 1031
rect 514 963 525 997
rect 559 963 570 997
rect 514 929 570 963
rect 514 895 525 929
rect 559 895 570 929
rect 514 861 570 895
rect 514 827 525 861
rect 559 827 570 861
rect 514 793 570 827
rect 514 759 525 793
rect 559 759 570 793
rect 514 725 570 759
rect 514 691 525 725
rect 559 691 570 725
rect 514 657 570 691
rect 514 623 525 657
rect 559 623 570 657
rect 514 589 570 623
rect 514 555 525 589
rect 559 555 570 589
rect 514 521 570 555
rect 514 487 525 521
rect 559 487 570 521
rect 514 475 570 487
rect 670 1813 740 1875
rect 670 1779 688 1813
rect 722 1779 740 1813
rect 670 1745 740 1779
rect 670 1711 688 1745
rect 722 1711 740 1745
rect 670 1677 740 1711
rect 670 1643 688 1677
rect 722 1643 740 1677
rect 670 1609 740 1643
rect 670 1575 688 1609
rect 722 1575 740 1609
rect 670 1541 740 1575
rect 670 1507 688 1541
rect 722 1507 740 1541
rect 670 1473 740 1507
rect 670 1439 688 1473
rect 722 1439 740 1473
rect 670 1405 740 1439
rect 670 1371 688 1405
rect 722 1371 740 1405
rect 670 1337 740 1371
rect 670 1303 688 1337
rect 722 1303 740 1337
rect 670 1269 740 1303
rect 670 1235 688 1269
rect 722 1235 740 1269
rect 670 1201 740 1235
rect 670 1167 688 1201
rect 722 1167 740 1201
rect 670 1133 740 1167
rect 670 1099 688 1133
rect 722 1099 740 1133
rect 670 1065 740 1099
rect 670 1031 688 1065
rect 722 1031 740 1065
rect 670 997 740 1031
rect 670 963 688 997
rect 722 963 740 997
rect 670 929 740 963
rect 670 895 688 929
rect 722 895 740 929
rect 670 861 740 895
rect 670 827 688 861
rect 722 827 740 861
rect 670 793 740 827
rect 670 759 688 793
rect 722 759 740 793
rect 670 725 740 759
rect 670 691 688 725
rect 722 691 740 725
rect 670 657 740 691
rect 670 623 688 657
rect 722 623 740 657
rect 670 589 740 623
rect 670 555 688 589
rect 722 555 740 589
rect 670 521 740 555
rect 670 487 688 521
rect 722 487 740 521
rect 670 475 740 487
rect 840 1813 896 1875
rect 840 1779 851 1813
rect 885 1779 896 1813
rect 840 1745 896 1779
rect 840 1711 851 1745
rect 885 1711 896 1745
rect 840 1677 896 1711
rect 840 1643 851 1677
rect 885 1643 896 1677
rect 840 1609 896 1643
rect 840 1575 851 1609
rect 885 1575 896 1609
rect 840 1541 896 1575
rect 840 1507 851 1541
rect 885 1507 896 1541
rect 840 1473 896 1507
rect 840 1439 851 1473
rect 885 1439 896 1473
rect 840 1405 896 1439
rect 840 1371 851 1405
rect 885 1371 896 1405
rect 840 1337 896 1371
rect 840 1303 851 1337
rect 885 1303 896 1337
rect 840 1269 896 1303
rect 840 1235 851 1269
rect 885 1235 896 1269
rect 840 1201 896 1235
rect 840 1167 851 1201
rect 885 1167 896 1201
rect 840 1133 896 1167
rect 840 1099 851 1133
rect 885 1099 896 1133
rect 840 1065 896 1099
rect 840 1031 851 1065
rect 885 1031 896 1065
rect 840 997 896 1031
rect 840 963 851 997
rect 885 963 896 997
rect 840 929 896 963
rect 840 895 851 929
rect 885 895 896 929
rect 840 861 896 895
rect 840 827 851 861
rect 885 827 896 861
rect 840 793 896 827
rect 840 759 851 793
rect 885 759 896 793
rect 840 725 896 759
rect 840 691 851 725
rect 885 691 896 725
rect 840 657 896 691
rect 840 623 851 657
rect 885 623 896 657
rect 840 589 896 623
rect 840 555 851 589
rect 885 555 896 589
rect 840 521 896 555
rect 840 487 851 521
rect 885 487 896 521
rect 840 475 896 487
rect 996 1813 1066 1875
rect 996 1779 1014 1813
rect 1048 1779 1066 1813
rect 996 1745 1066 1779
rect 996 1711 1014 1745
rect 1048 1711 1066 1745
rect 996 1677 1066 1711
rect 996 1643 1014 1677
rect 1048 1643 1066 1677
rect 996 1609 1066 1643
rect 996 1575 1014 1609
rect 1048 1575 1066 1609
rect 996 1541 1066 1575
rect 996 1507 1014 1541
rect 1048 1507 1066 1541
rect 996 1473 1066 1507
rect 996 1439 1014 1473
rect 1048 1439 1066 1473
rect 996 1405 1066 1439
rect 996 1371 1014 1405
rect 1048 1371 1066 1405
rect 996 1337 1066 1371
rect 996 1303 1014 1337
rect 1048 1303 1066 1337
rect 996 1269 1066 1303
rect 996 1235 1014 1269
rect 1048 1235 1066 1269
rect 996 1201 1066 1235
rect 996 1167 1014 1201
rect 1048 1167 1066 1201
rect 996 1133 1066 1167
rect 996 1099 1014 1133
rect 1048 1099 1066 1133
rect 996 1065 1066 1099
rect 996 1031 1014 1065
rect 1048 1031 1066 1065
rect 996 997 1066 1031
rect 996 963 1014 997
rect 1048 963 1066 997
rect 996 929 1066 963
rect 996 895 1014 929
rect 1048 895 1066 929
rect 996 861 1066 895
rect 996 827 1014 861
rect 1048 827 1066 861
rect 996 793 1066 827
rect 996 759 1014 793
rect 1048 759 1066 793
rect 996 725 1066 759
rect 996 691 1014 725
rect 1048 691 1066 725
rect 996 657 1066 691
rect 996 623 1014 657
rect 1048 623 1066 657
rect 996 589 1066 623
rect 996 555 1014 589
rect 1048 555 1066 589
rect 996 521 1066 555
rect 996 487 1014 521
rect 1048 487 1066 521
rect 996 475 1066 487
rect 1166 1813 1222 1875
rect 1166 1779 1177 1813
rect 1211 1779 1222 1813
rect 1166 1745 1222 1779
rect 1166 1711 1177 1745
rect 1211 1711 1222 1745
rect 1166 1677 1222 1711
rect 1166 1643 1177 1677
rect 1211 1643 1222 1677
rect 1166 1609 1222 1643
rect 1166 1575 1177 1609
rect 1211 1575 1222 1609
rect 1166 1541 1222 1575
rect 1166 1507 1177 1541
rect 1211 1507 1222 1541
rect 1166 1473 1222 1507
rect 1166 1439 1177 1473
rect 1211 1439 1222 1473
rect 1166 1405 1222 1439
rect 1166 1371 1177 1405
rect 1211 1371 1222 1405
rect 1166 1337 1222 1371
rect 1166 1303 1177 1337
rect 1211 1303 1222 1337
rect 1166 1269 1222 1303
rect 1166 1235 1177 1269
rect 1211 1235 1222 1269
rect 1166 1201 1222 1235
rect 1166 1167 1177 1201
rect 1211 1167 1222 1201
rect 1166 1133 1222 1167
rect 1166 1099 1177 1133
rect 1211 1099 1222 1133
rect 1166 1065 1222 1099
rect 1166 1031 1177 1065
rect 1211 1031 1222 1065
rect 1166 997 1222 1031
rect 1166 963 1177 997
rect 1211 963 1222 997
rect 1166 929 1222 963
rect 1166 895 1177 929
rect 1211 895 1222 929
rect 1166 861 1222 895
rect 1166 827 1177 861
rect 1211 827 1222 861
rect 1166 793 1222 827
rect 1166 759 1177 793
rect 1211 759 1222 793
rect 1166 725 1222 759
rect 1166 691 1177 725
rect 1211 691 1222 725
rect 1166 657 1222 691
rect 1166 623 1177 657
rect 1211 623 1222 657
rect 1166 589 1222 623
rect 1166 555 1177 589
rect 1211 555 1222 589
rect 1166 521 1222 555
rect 1166 487 1177 521
rect 1211 487 1222 521
rect 1166 475 1222 487
rect 1322 1813 1385 1875
rect 1322 1779 1340 1813
rect 1374 1779 1385 1813
rect 1322 1745 1385 1779
rect 1322 1711 1340 1745
rect 1374 1711 1385 1745
rect 1322 1677 1385 1711
rect 1322 1643 1340 1677
rect 1374 1643 1385 1677
rect 1322 1609 1385 1643
rect 1322 1575 1340 1609
rect 1374 1575 1385 1609
rect 1322 1541 1385 1575
rect 1322 1507 1340 1541
rect 1374 1507 1385 1541
rect 1322 1473 1385 1507
rect 1322 1439 1340 1473
rect 1374 1439 1385 1473
rect 1322 1405 1385 1439
rect 1322 1371 1340 1405
rect 1374 1371 1385 1405
rect 1322 1337 1385 1371
rect 1322 1303 1340 1337
rect 1374 1303 1385 1337
rect 1322 1269 1385 1303
rect 1322 1235 1340 1269
rect 1374 1235 1385 1269
rect 1322 1201 1385 1235
rect 1322 1167 1340 1201
rect 1374 1167 1385 1201
rect 1322 1133 1385 1167
rect 1322 1099 1340 1133
rect 1374 1099 1385 1133
rect 1322 1065 1385 1099
rect 1322 1031 1340 1065
rect 1374 1031 1385 1065
rect 1322 997 1385 1031
rect 1322 963 1340 997
rect 1374 963 1385 997
rect 1322 929 1385 963
rect 1322 895 1340 929
rect 1374 895 1385 929
rect 1322 861 1385 895
rect 1322 827 1340 861
rect 1374 827 1385 861
rect 1322 793 1385 827
rect 1322 759 1340 793
rect 1374 759 1385 793
rect 1322 725 1385 759
rect 1322 691 1340 725
rect 1374 691 1385 725
rect 1322 657 1385 691
rect 1322 623 1340 657
rect 1374 623 1385 657
rect 1322 589 1385 623
rect 1322 555 1340 589
rect 1374 555 1385 589
rect 1322 521 1385 555
rect 1322 487 1340 521
rect 1374 487 1385 521
rect 1322 475 1385 487
rect 2235 1813 2291 1875
rect 2235 1779 2246 1813
rect 2280 1779 2291 1813
rect 2235 1745 2291 1779
rect 2235 1711 2246 1745
rect 2280 1711 2291 1745
rect 2235 1677 2291 1711
rect 2235 1643 2246 1677
rect 2280 1643 2291 1677
rect 2235 1609 2291 1643
rect 2235 1575 2246 1609
rect 2280 1575 2291 1609
rect 2235 1541 2291 1575
rect 2235 1507 2246 1541
rect 2280 1507 2291 1541
rect 2235 1473 2291 1507
rect 2235 1439 2246 1473
rect 2280 1439 2291 1473
rect 2235 1405 2291 1439
rect 2235 1371 2246 1405
rect 2280 1371 2291 1405
rect 2235 1337 2291 1371
rect 2235 1303 2246 1337
rect 2280 1303 2291 1337
rect 2235 1269 2291 1303
rect 2235 1235 2246 1269
rect 2280 1235 2291 1269
rect 2235 1201 2291 1235
rect 2235 1167 2246 1201
rect 2280 1167 2291 1201
rect 2235 1133 2291 1167
rect 2235 1099 2246 1133
rect 2280 1099 2291 1133
rect 2235 1065 2291 1099
rect 2235 1031 2246 1065
rect 2280 1031 2291 1065
rect 2235 997 2291 1031
rect 2235 963 2246 997
rect 2280 963 2291 997
rect 2235 929 2291 963
rect 2235 895 2246 929
rect 2280 895 2291 929
rect 2235 861 2291 895
rect 2235 827 2246 861
rect 2280 827 2291 861
rect 2235 793 2291 827
rect 2235 759 2246 793
rect 2280 759 2291 793
rect 2235 725 2291 759
rect 2235 691 2246 725
rect 2280 691 2291 725
rect 2235 657 2291 691
rect 2235 623 2246 657
rect 2280 623 2291 657
rect 2235 589 2291 623
rect 2235 555 2246 589
rect 2280 555 2291 589
rect 2235 521 2291 555
rect 2235 487 2246 521
rect 2280 487 2291 521
rect 2235 475 2291 487
rect 2391 1813 2461 1875
rect 2391 1779 2409 1813
rect 2443 1779 2461 1813
rect 2391 1745 2461 1779
rect 2391 1711 2409 1745
rect 2443 1711 2461 1745
rect 2391 1677 2461 1711
rect 2391 1643 2409 1677
rect 2443 1643 2461 1677
rect 2391 1609 2461 1643
rect 2391 1575 2409 1609
rect 2443 1575 2461 1609
rect 2391 1541 2461 1575
rect 2391 1507 2409 1541
rect 2443 1507 2461 1541
rect 2391 1473 2461 1507
rect 2391 1439 2409 1473
rect 2443 1439 2461 1473
rect 2391 1405 2461 1439
rect 2391 1371 2409 1405
rect 2443 1371 2461 1405
rect 2391 1337 2461 1371
rect 2391 1303 2409 1337
rect 2443 1303 2461 1337
rect 2391 1269 2461 1303
rect 2391 1235 2409 1269
rect 2443 1235 2461 1269
rect 2391 1201 2461 1235
rect 2391 1167 2409 1201
rect 2443 1167 2461 1201
rect 2391 1133 2461 1167
rect 2391 1099 2409 1133
rect 2443 1099 2461 1133
rect 2391 1065 2461 1099
rect 2391 1031 2409 1065
rect 2443 1031 2461 1065
rect 2391 997 2461 1031
rect 2391 963 2409 997
rect 2443 963 2461 997
rect 2391 929 2461 963
rect 2391 895 2409 929
rect 2443 895 2461 929
rect 2391 861 2461 895
rect 2391 827 2409 861
rect 2443 827 2461 861
rect 2391 793 2461 827
rect 2391 759 2409 793
rect 2443 759 2461 793
rect 2391 725 2461 759
rect 2391 691 2409 725
rect 2443 691 2461 725
rect 2391 657 2461 691
rect 2391 623 2409 657
rect 2443 623 2461 657
rect 2391 589 2461 623
rect 2391 555 2409 589
rect 2443 555 2461 589
rect 2391 521 2461 555
rect 2391 487 2409 521
rect 2443 487 2461 521
rect 2391 475 2461 487
rect 2561 1813 2617 1875
rect 2561 1779 2572 1813
rect 2606 1779 2617 1813
rect 2561 1745 2617 1779
rect 2561 1711 2572 1745
rect 2606 1711 2617 1745
rect 2561 1677 2617 1711
rect 2561 1643 2572 1677
rect 2606 1643 2617 1677
rect 2561 1609 2617 1643
rect 2561 1575 2572 1609
rect 2606 1575 2617 1609
rect 2561 1541 2617 1575
rect 2561 1507 2572 1541
rect 2606 1507 2617 1541
rect 2561 1473 2617 1507
rect 2561 1439 2572 1473
rect 2606 1439 2617 1473
rect 2561 1405 2617 1439
rect 2561 1371 2572 1405
rect 2606 1371 2617 1405
rect 2561 1337 2617 1371
rect 2561 1303 2572 1337
rect 2606 1303 2617 1337
rect 2561 1269 2617 1303
rect 2561 1235 2572 1269
rect 2606 1235 2617 1269
rect 2561 1201 2617 1235
rect 2561 1167 2572 1201
rect 2606 1167 2617 1201
rect 2561 1133 2617 1167
rect 2561 1099 2572 1133
rect 2606 1099 2617 1133
rect 2561 1065 2617 1099
rect 2561 1031 2572 1065
rect 2606 1031 2617 1065
rect 2561 997 2617 1031
rect 2561 963 2572 997
rect 2606 963 2617 997
rect 2561 929 2617 963
rect 2561 895 2572 929
rect 2606 895 2617 929
rect 2561 861 2617 895
rect 2561 827 2572 861
rect 2606 827 2617 861
rect 2561 793 2617 827
rect 2561 759 2572 793
rect 2606 759 2617 793
rect 2561 725 2617 759
rect 2561 691 2572 725
rect 2606 691 2617 725
rect 2561 657 2617 691
rect 2561 623 2572 657
rect 2606 623 2617 657
rect 2561 589 2617 623
rect 2561 555 2572 589
rect 2606 555 2617 589
rect 2561 521 2617 555
rect 2561 487 2572 521
rect 2606 487 2617 521
rect 2561 475 2617 487
rect 2717 1813 2787 1875
rect 2717 1779 2735 1813
rect 2769 1779 2787 1813
rect 2717 1745 2787 1779
rect 2717 1711 2735 1745
rect 2769 1711 2787 1745
rect 2717 1677 2787 1711
rect 2717 1643 2735 1677
rect 2769 1643 2787 1677
rect 2717 1609 2787 1643
rect 2717 1575 2735 1609
rect 2769 1575 2787 1609
rect 2717 1541 2787 1575
rect 2717 1507 2735 1541
rect 2769 1507 2787 1541
rect 2717 1473 2787 1507
rect 2717 1439 2735 1473
rect 2769 1439 2787 1473
rect 2717 1405 2787 1439
rect 2717 1371 2735 1405
rect 2769 1371 2787 1405
rect 2717 1337 2787 1371
rect 2717 1303 2735 1337
rect 2769 1303 2787 1337
rect 2717 1269 2787 1303
rect 2717 1235 2735 1269
rect 2769 1235 2787 1269
rect 2717 1201 2787 1235
rect 2717 1167 2735 1201
rect 2769 1167 2787 1201
rect 2717 1133 2787 1167
rect 2717 1099 2735 1133
rect 2769 1099 2787 1133
rect 2717 1065 2787 1099
rect 2717 1031 2735 1065
rect 2769 1031 2787 1065
rect 2717 997 2787 1031
rect 2717 963 2735 997
rect 2769 963 2787 997
rect 2717 929 2787 963
rect 2717 895 2735 929
rect 2769 895 2787 929
rect 2717 861 2787 895
rect 2717 827 2735 861
rect 2769 827 2787 861
rect 2717 793 2787 827
rect 2717 759 2735 793
rect 2769 759 2787 793
rect 2717 725 2787 759
rect 2717 691 2735 725
rect 2769 691 2787 725
rect 2717 657 2787 691
rect 2717 623 2735 657
rect 2769 623 2787 657
rect 2717 589 2787 623
rect 2717 555 2735 589
rect 2769 555 2787 589
rect 2717 521 2787 555
rect 2717 487 2735 521
rect 2769 487 2787 521
rect 2717 475 2787 487
rect 2887 1813 2943 1875
rect 2887 1779 2898 1813
rect 2932 1779 2943 1813
rect 2887 1745 2943 1779
rect 2887 1711 2898 1745
rect 2932 1711 2943 1745
rect 2887 1677 2943 1711
rect 2887 1643 2898 1677
rect 2932 1643 2943 1677
rect 2887 1609 2943 1643
rect 2887 1575 2898 1609
rect 2932 1575 2943 1609
rect 2887 1541 2943 1575
rect 2887 1507 2898 1541
rect 2932 1507 2943 1541
rect 2887 1473 2943 1507
rect 2887 1439 2898 1473
rect 2932 1439 2943 1473
rect 2887 1405 2943 1439
rect 2887 1371 2898 1405
rect 2932 1371 2943 1405
rect 2887 1337 2943 1371
rect 2887 1303 2898 1337
rect 2932 1303 2943 1337
rect 2887 1269 2943 1303
rect 2887 1235 2898 1269
rect 2932 1235 2943 1269
rect 2887 1201 2943 1235
rect 2887 1167 2898 1201
rect 2932 1167 2943 1201
rect 2887 1133 2943 1167
rect 2887 1099 2898 1133
rect 2932 1099 2943 1133
rect 2887 1065 2943 1099
rect 2887 1031 2898 1065
rect 2932 1031 2943 1065
rect 2887 997 2943 1031
rect 2887 963 2898 997
rect 2932 963 2943 997
rect 2887 929 2943 963
rect 2887 895 2898 929
rect 2932 895 2943 929
rect 2887 861 2943 895
rect 2887 827 2898 861
rect 2932 827 2943 861
rect 2887 793 2943 827
rect 2887 759 2898 793
rect 2932 759 2943 793
rect 2887 725 2943 759
rect 2887 691 2898 725
rect 2932 691 2943 725
rect 2887 657 2943 691
rect 2887 623 2898 657
rect 2932 623 2943 657
rect 2887 589 2943 623
rect 2887 555 2898 589
rect 2932 555 2943 589
rect 2887 521 2943 555
rect 2887 487 2898 521
rect 2932 487 2943 521
rect 2887 475 2943 487
rect 3043 1813 3106 1875
rect 3043 1779 3061 1813
rect 3095 1779 3106 1813
rect 3043 1745 3106 1779
rect 3043 1711 3061 1745
rect 3095 1711 3106 1745
rect 3043 1677 3106 1711
rect 3043 1643 3061 1677
rect 3095 1643 3106 1677
rect 3043 1609 3106 1643
rect 3043 1575 3061 1609
rect 3095 1575 3106 1609
rect 3043 1541 3106 1575
rect 3043 1507 3061 1541
rect 3095 1507 3106 1541
rect 3043 1473 3106 1507
rect 3043 1439 3061 1473
rect 3095 1439 3106 1473
rect 3043 1405 3106 1439
rect 3043 1371 3061 1405
rect 3095 1371 3106 1405
rect 3043 1337 3106 1371
rect 3043 1303 3061 1337
rect 3095 1303 3106 1337
rect 3043 1269 3106 1303
rect 3043 1235 3061 1269
rect 3095 1235 3106 1269
rect 3043 1201 3106 1235
rect 3043 1167 3061 1201
rect 3095 1167 3106 1201
rect 3043 1133 3106 1167
rect 3043 1099 3061 1133
rect 3095 1099 3106 1133
rect 3043 1065 3106 1099
rect 3043 1031 3061 1065
rect 3095 1031 3106 1065
rect 3043 997 3106 1031
rect 3043 963 3061 997
rect 3095 963 3106 997
rect 3043 929 3106 963
rect 3043 895 3061 929
rect 3095 895 3106 929
rect 3043 861 3106 895
rect 3043 827 3061 861
rect 3095 827 3106 861
rect 3043 793 3106 827
rect 3043 759 3061 793
rect 3095 759 3106 793
rect 3043 725 3106 759
rect 3043 691 3061 725
rect 3095 691 3106 725
rect 3043 657 3106 691
rect 3043 623 3061 657
rect 3095 623 3106 657
rect 3043 589 3106 623
rect 3043 555 3061 589
rect 3095 555 3106 589
rect 3043 521 3106 555
rect 3043 487 3061 521
rect 3095 487 3106 521
rect 3043 475 3106 487
<< mvndiffc >>
rect 4131 1779 4165 1813
rect 4131 1711 4165 1745
rect 4131 1643 4165 1677
rect 4131 1575 4165 1609
rect 4131 1507 4165 1541
rect 4131 1439 4165 1473
rect 4131 1371 4165 1405
rect 4131 1303 4165 1337
rect 4131 1235 4165 1269
rect 4131 1167 4165 1201
rect 4131 1099 4165 1133
rect 4131 1031 4165 1065
rect 4131 963 4165 997
rect 4131 895 4165 929
rect 4131 827 4165 861
rect 4131 759 4165 793
rect 4131 691 4165 725
rect 4131 623 4165 657
rect 4131 555 4165 589
rect 4131 487 4165 521
rect 4294 1779 4328 1813
rect 4294 1711 4328 1745
rect 4294 1643 4328 1677
rect 4294 1575 4328 1609
rect 4294 1507 4328 1541
rect 4294 1439 4328 1473
rect 4294 1371 4328 1405
rect 4294 1303 4328 1337
rect 4294 1235 4328 1269
rect 4294 1167 4328 1201
rect 4294 1099 4328 1133
rect 4294 1031 4328 1065
rect 4294 963 4328 997
rect 4294 895 4328 929
rect 4294 827 4328 861
rect 4294 759 4328 793
rect 4294 691 4328 725
rect 4294 623 4328 657
rect 4294 555 4328 589
rect 4294 487 4328 521
rect 4457 1779 4491 1813
rect 4457 1711 4491 1745
rect 4457 1643 4491 1677
rect 4457 1575 4491 1609
rect 4457 1507 4491 1541
rect 4457 1439 4491 1473
rect 4457 1371 4491 1405
rect 4457 1303 4491 1337
rect 4457 1235 4491 1269
rect 4457 1167 4491 1201
rect 4457 1099 4491 1133
rect 4457 1031 4491 1065
rect 4457 963 4491 997
rect 4457 895 4491 929
rect 4457 827 4491 861
rect 4457 759 4491 793
rect 4457 691 4491 725
rect 4457 623 4491 657
rect 4457 555 4491 589
rect 4457 487 4491 521
rect 4620 1779 4654 1813
rect 4620 1711 4654 1745
rect 4620 1643 4654 1677
rect 4620 1575 4654 1609
rect 4620 1507 4654 1541
rect 4620 1439 4654 1473
rect 4620 1371 4654 1405
rect 4620 1303 4654 1337
rect 4620 1235 4654 1269
rect 4620 1167 4654 1201
rect 4620 1099 4654 1133
rect 4620 1031 4654 1065
rect 4620 963 4654 997
rect 4620 895 4654 929
rect 4620 827 4654 861
rect 4620 759 4654 793
rect 4620 691 4654 725
rect 4620 623 4654 657
rect 4620 555 4654 589
rect 4620 487 4654 521
rect 4783 1779 4817 1813
rect 4783 1711 4817 1745
rect 4783 1643 4817 1677
rect 4783 1575 4817 1609
rect 4783 1507 4817 1541
rect 4783 1439 4817 1473
rect 4783 1371 4817 1405
rect 4783 1303 4817 1337
rect 4783 1235 4817 1269
rect 4783 1167 4817 1201
rect 4783 1099 4817 1133
rect 4783 1031 4817 1065
rect 4783 963 4817 997
rect 4783 895 4817 929
rect 4783 827 4817 861
rect 4783 759 4817 793
rect 4783 691 4817 725
rect 4783 623 4817 657
rect 4783 555 4817 589
rect 4783 487 4817 521
rect 4946 1779 4980 1813
rect 4946 1711 4980 1745
rect 4946 1643 4980 1677
rect 4946 1575 4980 1609
rect 4946 1507 4980 1541
rect 4946 1439 4980 1473
rect 4946 1371 4980 1405
rect 4946 1303 4980 1337
rect 4946 1235 4980 1269
rect 4946 1167 4980 1201
rect 4946 1099 4980 1133
rect 4946 1031 4980 1065
rect 4946 963 4980 997
rect 4946 895 4980 929
rect 4946 827 4980 861
rect 4946 759 4980 793
rect 4946 691 4980 725
rect 4946 623 4980 657
rect 4946 555 4980 589
rect 4946 487 4980 521
rect 5109 1779 5143 1813
rect 5109 1711 5143 1745
rect 5109 1643 5143 1677
rect 5109 1575 5143 1609
rect 5109 1507 5143 1541
rect 5109 1439 5143 1473
rect 5109 1371 5143 1405
rect 5109 1303 5143 1337
rect 5109 1235 5143 1269
rect 5109 1167 5143 1201
rect 5109 1099 5143 1133
rect 5109 1031 5143 1065
rect 5109 963 5143 997
rect 5109 895 5143 929
rect 5109 827 5143 861
rect 5109 759 5143 793
rect 5109 691 5143 725
rect 5109 623 5143 657
rect 5109 555 5143 589
rect 5109 487 5143 521
rect 5272 1779 5306 1813
rect 5272 1711 5306 1745
rect 5272 1643 5306 1677
rect 5272 1575 5306 1609
rect 5272 1507 5306 1541
rect 5272 1439 5306 1473
rect 5272 1371 5306 1405
rect 5272 1303 5306 1337
rect 5272 1235 5306 1269
rect 5272 1167 5306 1201
rect 5272 1099 5306 1133
rect 5272 1031 5306 1065
rect 5272 963 5306 997
rect 5272 895 5306 929
rect 5272 827 5306 861
rect 5272 759 5306 793
rect 5272 691 5306 725
rect 5272 623 5306 657
rect 5272 555 5306 589
rect 5272 487 5306 521
rect 5395 1779 5429 1813
rect 5395 1711 5429 1745
rect 5395 1643 5429 1677
rect 5395 1575 5429 1609
rect 5395 1507 5429 1541
rect 5395 1439 5429 1473
rect 5395 1371 5429 1405
rect 5395 1303 5429 1337
rect 5395 1235 5429 1269
rect 5395 1167 5429 1201
rect 5395 1099 5429 1133
rect 5395 1031 5429 1065
rect 5395 963 5429 997
rect 5395 895 5429 929
rect 5395 827 5429 861
rect 5395 759 5429 793
rect 5395 691 5429 725
rect 5395 623 5429 657
rect 5395 555 5429 589
rect 5395 487 5429 521
rect 5558 1779 5592 1813
rect 5558 1711 5592 1745
rect 5558 1643 5592 1677
rect 5558 1575 5592 1609
rect 5558 1507 5592 1541
rect 5558 1439 5592 1473
rect 5558 1371 5592 1405
rect 5558 1303 5592 1337
rect 5558 1235 5592 1269
rect 5558 1167 5592 1201
rect 5558 1099 5592 1133
rect 5558 1031 5592 1065
rect 5558 963 5592 997
rect 5558 895 5592 929
rect 5558 827 5592 861
rect 5558 759 5592 793
rect 5558 691 5592 725
rect 5558 623 5592 657
rect 5558 555 5592 589
rect 5558 487 5592 521
rect 5721 1779 5755 1813
rect 5721 1711 5755 1745
rect 5721 1643 5755 1677
rect 5721 1575 5755 1609
rect 5721 1507 5755 1541
rect 5721 1439 5755 1473
rect 5721 1371 5755 1405
rect 5721 1303 5755 1337
rect 5721 1235 5755 1269
rect 5721 1167 5755 1201
rect 5721 1099 5755 1133
rect 5721 1031 5755 1065
rect 5721 963 5755 997
rect 5721 895 5755 929
rect 5721 827 5755 861
rect 5721 759 5755 793
rect 5721 691 5755 725
rect 5721 623 5755 657
rect 5721 555 5755 589
rect 5721 487 5755 521
rect 5884 1779 5918 1813
rect 5884 1711 5918 1745
rect 5884 1643 5918 1677
rect 5884 1575 5918 1609
rect 5884 1507 5918 1541
rect 5884 1439 5918 1473
rect 5884 1371 5918 1405
rect 5884 1303 5918 1337
rect 5884 1235 5918 1269
rect 5884 1167 5918 1201
rect 5884 1099 5918 1133
rect 5884 1031 5918 1065
rect 5884 963 5918 997
rect 5884 895 5918 929
rect 5884 827 5918 861
rect 5884 759 5918 793
rect 5884 691 5918 725
rect 5884 623 5918 657
rect 5884 555 5918 589
rect 5884 487 5918 521
rect 6047 1779 6081 1813
rect 6047 1711 6081 1745
rect 6047 1643 6081 1677
rect 6047 1575 6081 1609
rect 6047 1507 6081 1541
rect 6047 1439 6081 1473
rect 6047 1371 6081 1405
rect 6047 1303 6081 1337
rect 6047 1235 6081 1269
rect 6047 1167 6081 1201
rect 6047 1099 6081 1133
rect 6047 1031 6081 1065
rect 6047 963 6081 997
rect 6047 895 6081 929
rect 6047 827 6081 861
rect 6047 759 6081 793
rect 6047 691 6081 725
rect 6047 623 6081 657
rect 6047 555 6081 589
rect 6047 487 6081 521
rect 6210 1779 6244 1813
rect 6210 1711 6244 1745
rect 6210 1643 6244 1677
rect 6210 1575 6244 1609
rect 6210 1507 6244 1541
rect 6210 1439 6244 1473
rect 6210 1371 6244 1405
rect 6210 1303 6244 1337
rect 6210 1235 6244 1269
rect 6210 1167 6244 1201
rect 6210 1099 6244 1133
rect 6210 1031 6244 1065
rect 6210 963 6244 997
rect 6210 895 6244 929
rect 6210 827 6244 861
rect 6210 759 6244 793
rect 6210 691 6244 725
rect 6210 623 6244 657
rect 6210 555 6244 589
rect 6210 487 6244 521
rect 6373 1779 6407 1813
rect 6373 1711 6407 1745
rect 6373 1643 6407 1677
rect 6373 1575 6407 1609
rect 6373 1507 6407 1541
rect 6373 1439 6407 1473
rect 6373 1371 6407 1405
rect 6373 1303 6407 1337
rect 6373 1235 6407 1269
rect 6373 1167 6407 1201
rect 6373 1099 6407 1133
rect 6373 1031 6407 1065
rect 6373 963 6407 997
rect 6373 895 6407 929
rect 6373 827 6407 861
rect 6373 759 6407 793
rect 6373 691 6407 725
rect 6373 623 6407 657
rect 6373 555 6407 589
rect 6373 487 6407 521
rect 6536 1779 6570 1813
rect 6536 1711 6570 1745
rect 6536 1643 6570 1677
rect 6536 1575 6570 1609
rect 6536 1507 6570 1541
rect 6536 1439 6570 1473
rect 6536 1371 6570 1405
rect 6536 1303 6570 1337
rect 6536 1235 6570 1269
rect 6536 1167 6570 1201
rect 6536 1099 6570 1133
rect 6536 1031 6570 1065
rect 6536 963 6570 997
rect 6536 895 6570 929
rect 6536 827 6570 861
rect 6536 759 6570 793
rect 6536 691 6570 725
rect 6536 623 6570 657
rect 6536 555 6570 589
rect 6536 487 6570 521
rect 7216 1847 7250 1881
rect 7216 1779 7250 1813
rect 7216 1711 7250 1745
rect 7216 1643 7250 1677
rect 7216 1575 7250 1609
rect 7216 1507 7250 1541
rect 7216 1439 7250 1473
rect 7216 1371 7250 1405
rect 7216 1303 7250 1337
rect 7216 1235 7250 1269
rect 7216 1167 7250 1201
rect 7216 1099 7250 1133
rect 7216 1031 7250 1065
rect 7216 963 7250 997
rect 7216 895 7250 929
rect 7216 827 7250 861
rect 7216 759 7250 793
rect 7216 691 7250 725
rect 7216 623 7250 657
rect 7216 555 7250 589
rect 7379 1847 7413 1881
rect 7379 1779 7413 1813
rect 7379 1711 7413 1745
rect 7379 1643 7413 1677
rect 7379 1575 7413 1609
rect 7379 1507 7413 1541
rect 7379 1439 7413 1473
rect 7379 1371 7413 1405
rect 7379 1303 7413 1337
rect 7379 1235 7413 1269
rect 7379 1167 7413 1201
rect 7379 1099 7413 1133
rect 7379 1031 7413 1065
rect 7379 963 7413 997
rect 7379 895 7413 929
rect 7379 827 7413 861
rect 7379 759 7413 793
rect 7379 691 7413 725
rect 7379 623 7413 657
rect 7379 555 7413 589
rect 7542 1847 7576 1881
rect 7542 1779 7576 1813
rect 7542 1711 7576 1745
rect 7542 1643 7576 1677
rect 7542 1575 7576 1609
rect 7542 1507 7576 1541
rect 7542 1439 7576 1473
rect 7542 1371 7576 1405
rect 7542 1303 7576 1337
rect 7542 1235 7576 1269
rect 7542 1167 7576 1201
rect 7542 1099 7576 1133
rect 7542 1031 7576 1065
rect 7542 963 7576 997
rect 7542 895 7576 929
rect 7542 827 7576 861
rect 7542 759 7576 793
rect 7542 691 7576 725
rect 7542 623 7576 657
rect 7542 555 7576 589
rect 7705 1847 7739 1881
rect 7705 1779 7739 1813
rect 7705 1711 7739 1745
rect 7705 1643 7739 1677
rect 7705 1575 7739 1609
rect 7705 1507 7739 1541
rect 7705 1439 7739 1473
rect 7705 1371 7739 1405
rect 7705 1303 7739 1337
rect 7705 1235 7739 1269
rect 7705 1167 7739 1201
rect 7705 1099 7739 1133
rect 7705 1031 7739 1065
rect 7705 963 7739 997
rect 7705 895 7739 929
rect 7705 827 7739 861
rect 7705 759 7739 793
rect 7705 691 7739 725
rect 7705 623 7739 657
rect 7705 555 7739 589
rect 7868 1847 7902 1881
rect 7868 1779 7902 1813
rect 7868 1711 7902 1745
rect 7868 1643 7902 1677
rect 7868 1575 7902 1609
rect 7868 1507 7902 1541
rect 7868 1439 7902 1473
rect 7868 1371 7902 1405
rect 7868 1303 7902 1337
rect 7868 1235 7902 1269
rect 7868 1167 7902 1201
rect 7868 1099 7902 1133
rect 7868 1031 7902 1065
rect 7868 963 7902 997
rect 7868 895 7902 929
rect 7868 827 7902 861
rect 7868 759 7902 793
rect 7868 691 7902 725
rect 7868 623 7902 657
rect 7868 555 7902 589
rect 8031 1847 8065 1881
rect 8031 1779 8065 1813
rect 8031 1711 8065 1745
rect 8031 1643 8065 1677
rect 8031 1575 8065 1609
rect 8031 1507 8065 1541
rect 8031 1439 8065 1473
rect 8031 1371 8065 1405
rect 8031 1303 8065 1337
rect 8031 1235 8065 1269
rect 8031 1167 8065 1201
rect 8031 1099 8065 1133
rect 8031 1031 8065 1065
rect 8031 963 8065 997
rect 8031 895 8065 929
rect 8031 827 8065 861
rect 8031 759 8065 793
rect 8031 691 8065 725
rect 8031 623 8065 657
rect 8031 555 8065 589
rect 8194 1847 8228 1881
rect 8194 1779 8228 1813
rect 8194 1711 8228 1745
rect 8194 1643 8228 1677
rect 8194 1575 8228 1609
rect 8194 1507 8228 1541
rect 8194 1439 8228 1473
rect 8194 1371 8228 1405
rect 8194 1303 8228 1337
rect 8194 1235 8228 1269
rect 8194 1167 8228 1201
rect 8194 1099 8228 1133
rect 8194 1031 8228 1065
rect 8194 963 8228 997
rect 8194 895 8228 929
rect 8194 827 8228 861
rect 8194 759 8228 793
rect 8194 691 8228 725
rect 8194 623 8228 657
rect 8194 555 8228 589
rect 8357 1847 8391 1881
rect 8357 1779 8391 1813
rect 8357 1711 8391 1745
rect 8357 1643 8391 1677
rect 8357 1575 8391 1609
rect 8357 1507 8391 1541
rect 8357 1439 8391 1473
rect 8357 1371 8391 1405
rect 8357 1303 8391 1337
rect 8357 1235 8391 1269
rect 8357 1167 8391 1201
rect 8357 1099 8391 1133
rect 8357 1031 8391 1065
rect 8357 963 8391 997
rect 8357 895 8391 929
rect 8357 827 8391 861
rect 8357 759 8391 793
rect 8357 691 8391 725
rect 8357 623 8391 657
rect 8357 555 8391 589
rect 8480 1847 8514 1881
rect 8480 1779 8514 1813
rect 8480 1711 8514 1745
rect 8480 1643 8514 1677
rect 8480 1575 8514 1609
rect 8480 1507 8514 1541
rect 8480 1439 8514 1473
rect 8480 1371 8514 1405
rect 8480 1303 8514 1337
rect 8480 1235 8514 1269
rect 8480 1167 8514 1201
rect 8480 1099 8514 1133
rect 8480 1031 8514 1065
rect 8480 963 8514 997
rect 8480 895 8514 929
rect 8480 827 8514 861
rect 8480 759 8514 793
rect 8480 691 8514 725
rect 8480 623 8514 657
rect 8480 555 8514 589
rect 8643 1847 8677 1881
rect 8643 1779 8677 1813
rect 8643 1711 8677 1745
rect 8643 1643 8677 1677
rect 8643 1575 8677 1609
rect 8643 1507 8677 1541
rect 8643 1439 8677 1473
rect 8643 1371 8677 1405
rect 8643 1303 8677 1337
rect 8643 1235 8677 1269
rect 8643 1167 8677 1201
rect 8643 1099 8677 1133
rect 8643 1031 8677 1065
rect 8643 963 8677 997
rect 8643 895 8677 929
rect 8643 827 8677 861
rect 8643 759 8677 793
rect 8643 691 8677 725
rect 8643 623 8677 657
rect 8643 555 8677 589
rect 8806 1847 8840 1881
rect 8806 1779 8840 1813
rect 8806 1711 8840 1745
rect 8806 1643 8840 1677
rect 8806 1575 8840 1609
rect 8806 1507 8840 1541
rect 8806 1439 8840 1473
rect 8806 1371 8840 1405
rect 8806 1303 8840 1337
rect 8806 1235 8840 1269
rect 8806 1167 8840 1201
rect 8806 1099 8840 1133
rect 8806 1031 8840 1065
rect 8806 963 8840 997
rect 8806 895 8840 929
rect 8806 827 8840 861
rect 8806 759 8840 793
rect 8806 691 8840 725
rect 8806 623 8840 657
rect 8806 555 8840 589
rect 8969 1847 9003 1881
rect 8969 1779 9003 1813
rect 8969 1711 9003 1745
rect 8969 1643 9003 1677
rect 8969 1575 9003 1609
rect 8969 1507 9003 1541
rect 8969 1439 9003 1473
rect 8969 1371 9003 1405
rect 8969 1303 9003 1337
rect 8969 1235 9003 1269
rect 8969 1167 9003 1201
rect 8969 1099 9003 1133
rect 8969 1031 9003 1065
rect 8969 963 9003 997
rect 8969 895 9003 929
rect 8969 827 9003 861
rect 8969 759 9003 793
rect 8969 691 9003 725
rect 8969 623 9003 657
rect 8969 555 9003 589
rect 9132 1847 9166 1881
rect 9132 1779 9166 1813
rect 9132 1711 9166 1745
rect 9132 1643 9166 1677
rect 9132 1575 9166 1609
rect 9132 1507 9166 1541
rect 9132 1439 9166 1473
rect 9132 1371 9166 1405
rect 9132 1303 9166 1337
rect 9132 1235 9166 1269
rect 9132 1167 9166 1201
rect 9132 1099 9166 1133
rect 9132 1031 9166 1065
rect 9132 963 9166 997
rect 9132 895 9166 929
rect 9132 827 9166 861
rect 9132 759 9166 793
rect 9132 691 9166 725
rect 9132 623 9166 657
rect 9132 555 9166 589
rect 9295 1847 9329 1881
rect 9295 1779 9329 1813
rect 9295 1711 9329 1745
rect 9295 1643 9329 1677
rect 9295 1575 9329 1609
rect 9295 1507 9329 1541
rect 9295 1439 9329 1473
rect 9295 1371 9329 1405
rect 9295 1303 9329 1337
rect 9295 1235 9329 1269
rect 9295 1167 9329 1201
rect 9295 1099 9329 1133
rect 9295 1031 9329 1065
rect 9295 963 9329 997
rect 9295 895 9329 929
rect 9295 827 9329 861
rect 9295 759 9329 793
rect 9295 691 9329 725
rect 9295 623 9329 657
rect 9295 555 9329 589
rect 9458 1847 9492 1881
rect 9458 1779 9492 1813
rect 9458 1711 9492 1745
rect 9458 1643 9492 1677
rect 9458 1575 9492 1609
rect 9458 1507 9492 1541
rect 9458 1439 9492 1473
rect 9458 1371 9492 1405
rect 9458 1303 9492 1337
rect 9458 1235 9492 1269
rect 9458 1167 9492 1201
rect 9458 1099 9492 1133
rect 9458 1031 9492 1065
rect 9458 963 9492 997
rect 9458 895 9492 929
rect 9458 827 9492 861
rect 9458 759 9492 793
rect 9458 691 9492 725
rect 9458 623 9492 657
rect 9458 555 9492 589
rect 9621 1847 9655 1881
rect 9621 1779 9655 1813
rect 9621 1711 9655 1745
rect 9621 1643 9655 1677
rect 9621 1575 9655 1609
rect 9621 1507 9655 1541
rect 9621 1439 9655 1473
rect 9621 1371 9655 1405
rect 9621 1303 9655 1337
rect 9621 1235 9655 1269
rect 9621 1167 9655 1201
rect 9621 1099 9655 1133
rect 9621 1031 9655 1065
rect 9621 963 9655 997
rect 9621 895 9655 929
rect 9621 827 9655 861
rect 9621 759 9655 793
rect 9621 691 9655 725
rect 9621 623 9655 657
rect 9621 555 9655 589
rect 9784 1847 9818 1881
rect 9784 1779 9818 1813
rect 9784 1711 9818 1745
rect 9784 1643 9818 1677
rect 9784 1575 9818 1609
rect 9784 1507 9818 1541
rect 9784 1439 9818 1473
rect 9784 1371 9818 1405
rect 9784 1303 9818 1337
rect 9784 1235 9818 1269
rect 9784 1167 9818 1201
rect 9784 1099 9818 1133
rect 9784 1031 9818 1065
rect 9784 963 9818 997
rect 9784 895 9818 929
rect 9784 827 9818 861
rect 9784 759 9818 793
rect 9784 691 9818 725
rect 9784 623 9818 657
rect 9784 555 9818 589
<< mvpdiffc >>
rect 362 1779 396 1813
rect 362 1711 396 1745
rect 362 1643 396 1677
rect 362 1575 396 1609
rect 362 1507 396 1541
rect 362 1439 396 1473
rect 362 1371 396 1405
rect 362 1303 396 1337
rect 362 1235 396 1269
rect 362 1167 396 1201
rect 362 1099 396 1133
rect 362 1031 396 1065
rect 362 963 396 997
rect 362 895 396 929
rect 362 827 396 861
rect 362 759 396 793
rect 362 691 396 725
rect 362 623 396 657
rect 362 555 396 589
rect 362 487 396 521
rect 525 1779 559 1813
rect 525 1711 559 1745
rect 525 1643 559 1677
rect 525 1575 559 1609
rect 525 1507 559 1541
rect 525 1439 559 1473
rect 525 1371 559 1405
rect 525 1303 559 1337
rect 525 1235 559 1269
rect 525 1167 559 1201
rect 525 1099 559 1133
rect 525 1031 559 1065
rect 525 963 559 997
rect 525 895 559 929
rect 525 827 559 861
rect 525 759 559 793
rect 525 691 559 725
rect 525 623 559 657
rect 525 555 559 589
rect 525 487 559 521
rect 688 1779 722 1813
rect 688 1711 722 1745
rect 688 1643 722 1677
rect 688 1575 722 1609
rect 688 1507 722 1541
rect 688 1439 722 1473
rect 688 1371 722 1405
rect 688 1303 722 1337
rect 688 1235 722 1269
rect 688 1167 722 1201
rect 688 1099 722 1133
rect 688 1031 722 1065
rect 688 963 722 997
rect 688 895 722 929
rect 688 827 722 861
rect 688 759 722 793
rect 688 691 722 725
rect 688 623 722 657
rect 688 555 722 589
rect 688 487 722 521
rect 851 1779 885 1813
rect 851 1711 885 1745
rect 851 1643 885 1677
rect 851 1575 885 1609
rect 851 1507 885 1541
rect 851 1439 885 1473
rect 851 1371 885 1405
rect 851 1303 885 1337
rect 851 1235 885 1269
rect 851 1167 885 1201
rect 851 1099 885 1133
rect 851 1031 885 1065
rect 851 963 885 997
rect 851 895 885 929
rect 851 827 885 861
rect 851 759 885 793
rect 851 691 885 725
rect 851 623 885 657
rect 851 555 885 589
rect 851 487 885 521
rect 1014 1779 1048 1813
rect 1014 1711 1048 1745
rect 1014 1643 1048 1677
rect 1014 1575 1048 1609
rect 1014 1507 1048 1541
rect 1014 1439 1048 1473
rect 1014 1371 1048 1405
rect 1014 1303 1048 1337
rect 1014 1235 1048 1269
rect 1014 1167 1048 1201
rect 1014 1099 1048 1133
rect 1014 1031 1048 1065
rect 1014 963 1048 997
rect 1014 895 1048 929
rect 1014 827 1048 861
rect 1014 759 1048 793
rect 1014 691 1048 725
rect 1014 623 1048 657
rect 1014 555 1048 589
rect 1014 487 1048 521
rect 1177 1779 1211 1813
rect 1177 1711 1211 1745
rect 1177 1643 1211 1677
rect 1177 1575 1211 1609
rect 1177 1507 1211 1541
rect 1177 1439 1211 1473
rect 1177 1371 1211 1405
rect 1177 1303 1211 1337
rect 1177 1235 1211 1269
rect 1177 1167 1211 1201
rect 1177 1099 1211 1133
rect 1177 1031 1211 1065
rect 1177 963 1211 997
rect 1177 895 1211 929
rect 1177 827 1211 861
rect 1177 759 1211 793
rect 1177 691 1211 725
rect 1177 623 1211 657
rect 1177 555 1211 589
rect 1177 487 1211 521
rect 1340 1779 1374 1813
rect 1340 1711 1374 1745
rect 1340 1643 1374 1677
rect 1340 1575 1374 1609
rect 1340 1507 1374 1541
rect 1340 1439 1374 1473
rect 1340 1371 1374 1405
rect 1340 1303 1374 1337
rect 1340 1235 1374 1269
rect 1340 1167 1374 1201
rect 1340 1099 1374 1133
rect 1340 1031 1374 1065
rect 1340 963 1374 997
rect 1340 895 1374 929
rect 1340 827 1374 861
rect 1340 759 1374 793
rect 1340 691 1374 725
rect 1340 623 1374 657
rect 1340 555 1374 589
rect 1340 487 1374 521
rect 2246 1779 2280 1813
rect 2246 1711 2280 1745
rect 2246 1643 2280 1677
rect 2246 1575 2280 1609
rect 2246 1507 2280 1541
rect 2246 1439 2280 1473
rect 2246 1371 2280 1405
rect 2246 1303 2280 1337
rect 2246 1235 2280 1269
rect 2246 1167 2280 1201
rect 2246 1099 2280 1133
rect 2246 1031 2280 1065
rect 2246 963 2280 997
rect 2246 895 2280 929
rect 2246 827 2280 861
rect 2246 759 2280 793
rect 2246 691 2280 725
rect 2246 623 2280 657
rect 2246 555 2280 589
rect 2246 487 2280 521
rect 2409 1779 2443 1813
rect 2409 1711 2443 1745
rect 2409 1643 2443 1677
rect 2409 1575 2443 1609
rect 2409 1507 2443 1541
rect 2409 1439 2443 1473
rect 2409 1371 2443 1405
rect 2409 1303 2443 1337
rect 2409 1235 2443 1269
rect 2409 1167 2443 1201
rect 2409 1099 2443 1133
rect 2409 1031 2443 1065
rect 2409 963 2443 997
rect 2409 895 2443 929
rect 2409 827 2443 861
rect 2409 759 2443 793
rect 2409 691 2443 725
rect 2409 623 2443 657
rect 2409 555 2443 589
rect 2409 487 2443 521
rect 2572 1779 2606 1813
rect 2572 1711 2606 1745
rect 2572 1643 2606 1677
rect 2572 1575 2606 1609
rect 2572 1507 2606 1541
rect 2572 1439 2606 1473
rect 2572 1371 2606 1405
rect 2572 1303 2606 1337
rect 2572 1235 2606 1269
rect 2572 1167 2606 1201
rect 2572 1099 2606 1133
rect 2572 1031 2606 1065
rect 2572 963 2606 997
rect 2572 895 2606 929
rect 2572 827 2606 861
rect 2572 759 2606 793
rect 2572 691 2606 725
rect 2572 623 2606 657
rect 2572 555 2606 589
rect 2572 487 2606 521
rect 2735 1779 2769 1813
rect 2735 1711 2769 1745
rect 2735 1643 2769 1677
rect 2735 1575 2769 1609
rect 2735 1507 2769 1541
rect 2735 1439 2769 1473
rect 2735 1371 2769 1405
rect 2735 1303 2769 1337
rect 2735 1235 2769 1269
rect 2735 1167 2769 1201
rect 2735 1099 2769 1133
rect 2735 1031 2769 1065
rect 2735 963 2769 997
rect 2735 895 2769 929
rect 2735 827 2769 861
rect 2735 759 2769 793
rect 2735 691 2769 725
rect 2735 623 2769 657
rect 2735 555 2769 589
rect 2735 487 2769 521
rect 2898 1779 2932 1813
rect 2898 1711 2932 1745
rect 2898 1643 2932 1677
rect 2898 1575 2932 1609
rect 2898 1507 2932 1541
rect 2898 1439 2932 1473
rect 2898 1371 2932 1405
rect 2898 1303 2932 1337
rect 2898 1235 2932 1269
rect 2898 1167 2932 1201
rect 2898 1099 2932 1133
rect 2898 1031 2932 1065
rect 2898 963 2932 997
rect 2898 895 2932 929
rect 2898 827 2932 861
rect 2898 759 2932 793
rect 2898 691 2932 725
rect 2898 623 2932 657
rect 2898 555 2932 589
rect 2898 487 2932 521
rect 3061 1779 3095 1813
rect 3061 1711 3095 1745
rect 3061 1643 3095 1677
rect 3061 1575 3095 1609
rect 3061 1507 3095 1541
rect 3061 1439 3095 1473
rect 3061 1371 3095 1405
rect 3061 1303 3095 1337
rect 3061 1235 3095 1269
rect 3061 1167 3095 1201
rect 3061 1099 3095 1133
rect 3061 1031 3095 1065
rect 3061 963 3095 997
rect 3061 895 3095 929
rect 3061 827 3095 861
rect 3061 759 3095 793
rect 3061 691 3095 725
rect 3061 623 3095 657
rect 3061 555 3095 589
rect 3061 487 3095 521
<< psubdiff >>
rect 1647 424 1648 447
rect 1682 424 1720 447
rect 1754 424 1792 447
rect 1826 424 1864 447
rect 1898 424 1899 447
rect 1647 390 1899 424
rect -24 177 78 211
rect 10 143 78 177
rect -24 138 78 143
rect 1647 356 1648 390
rect 1682 356 1720 390
rect 1754 356 1792 390
rect 1826 356 1864 390
rect 1898 356 1899 390
rect 1647 322 1899 356
rect 1647 288 1648 322
rect 1682 288 1720 322
rect 1754 288 1792 322
rect 1826 288 1864 322
rect 1898 288 1899 322
rect 1647 254 1899 288
rect 1647 220 1648 254
rect 1682 220 1720 254
rect 1754 220 1792 254
rect 1826 220 1864 254
rect 1898 220 1899 254
rect 1647 138 1899 220
rect -24 36 44 138
rect 3342 104 3435 138
rect 3342 70 3537 104
rect 3342 36 3376 70
rect 3410 36 3537 70
rect 4005 367 4039 447
rect 6655 435 6689 447
rect 6655 367 6689 401
rect 4005 333 4073 367
rect 4107 333 4141 367
rect 4175 333 4209 367
rect 4243 333 4277 367
rect 4311 333 4345 367
rect 4379 333 4413 367
rect 4447 333 4481 367
rect 4515 333 4549 367
rect 4583 333 4617 367
rect 4651 333 4685 367
rect 4719 333 4753 367
rect 4787 333 4821 367
rect 4855 333 4889 367
rect 4923 333 4957 367
rect 4991 333 5025 367
rect 5059 333 5093 367
rect 5127 333 5161 367
rect 5195 333 5229 367
rect 5263 333 5297 367
rect 5331 333 5365 367
rect 5399 333 5433 367
rect 5467 333 5501 367
rect 5535 333 5569 367
rect 5603 333 5637 367
rect 5671 333 5705 367
rect 5739 333 5773 367
rect 5807 333 5841 367
rect 5875 333 5909 367
rect 5943 333 5977 367
rect 6011 333 6045 367
rect 6079 333 6113 367
rect 6147 333 6181 367
rect 6215 333 6249 367
rect 6283 333 6317 367
rect 6351 333 6385 367
rect 6419 333 6453 367
rect 6487 333 6521 367
rect 6555 333 6689 367
rect 7097 435 7165 447
rect 7199 435 7233 447
rect 7267 435 7301 447
rect 7335 435 7369 447
rect 7403 435 7437 447
rect 7471 435 7505 447
rect 7539 435 7573 447
rect 7607 435 7641 447
rect 7675 435 7709 447
rect 7743 435 7777 447
rect 7811 435 7845 447
rect 7879 435 7913 447
rect 7947 435 7981 447
rect 8015 435 8049 447
rect 8083 435 8117 447
rect 8151 435 8185 447
rect 8219 435 8253 447
rect 8287 435 8321 447
rect 8355 435 8389 447
rect 8423 435 8457 447
rect 8491 435 8525 447
rect 8559 435 8593 447
rect 8627 435 8661 447
rect 8695 435 8729 447
rect 8763 435 8797 447
rect 8831 435 8865 447
rect 8899 435 8933 447
rect 8967 435 9001 447
rect 9035 435 9069 447
rect 9103 435 9137 447
rect 9171 435 9205 447
rect 9239 435 9273 447
rect 9307 435 9341 447
rect 9375 435 9409 447
rect 9443 435 9477 447
rect 9511 435 9545 447
rect 9579 435 9613 447
rect 9647 435 9681 447
rect 9715 435 9749 447
rect 9783 435 9817 447
rect 9851 435 9885 447
rect 9919 435 9997 447
<< nsubdiff >>
rect 237 395 271 447
rect 1459 395 1493 429
rect 237 361 305 395
rect 339 361 373 395
rect 407 361 441 395
rect 475 361 509 395
rect 543 361 577 395
rect 611 361 645 395
rect 679 361 713 395
rect 747 361 781 395
rect 815 361 849 395
rect 883 361 917 395
rect 951 361 985 395
rect 1019 361 1053 395
rect 1087 361 1121 395
rect 1155 361 1189 395
rect 1223 361 1257 395
rect 1291 361 1325 395
rect 1359 361 1493 395
rect 3180 434 3282 447
rect 3180 400 3248 434
rect 3180 393 3282 400
rect 2154 359 2228 393
rect 2052 325 2228 359
rect 2052 291 2160 325
rect 2194 291 2228 325
rect 3214 291 3282 393
rect 3750 418 3852 447
rect 10160 438 10228 447
rect 10160 322 10262 336
rect 10160 288 10228 322
rect 10160 254 10262 288
rect 10160 248 10228 254
rect 7010 182 7032 248
rect 6842 180 7032 182
rect 6842 146 6910 180
rect 6944 146 7032 180
rect 10194 220 10228 248
rect 10194 146 10262 220
rect 3852 112 3918 146
rect 3750 78 3918 112
rect 3750 44 3850 78
rect 3884 44 3918 78
rect 6876 44 6944 146
<< mvpsubdiff >>
rect -24 2260 69 2362
rect 3503 2260 3537 2362
rect -24 2226 78 2260
rect 1647 2226 1899 2260
rect 1647 2192 1648 2226
rect 1682 2192 1720 2226
rect 1754 2192 1792 2226
rect 1826 2192 1864 2226
rect 1898 2192 1899 2226
rect 1647 2158 1899 2192
rect 1647 2124 1648 2158
rect 1682 2124 1720 2158
rect 1754 2124 1792 2158
rect 1826 2124 1864 2158
rect 1898 2124 1899 2158
rect -24 1265 78 1376
rect 1647 2090 1899 2124
rect 3435 2178 3537 2260
rect 1647 2056 1648 2090
rect 1682 2056 1720 2090
rect 1754 2056 1792 2090
rect 1826 2056 1864 2090
rect 1898 2056 1899 2090
rect 1647 2022 1899 2056
rect 1647 1988 1648 2022
rect 1682 1988 1720 2022
rect 1754 1988 1792 2022
rect 1826 1988 1864 2022
rect 1898 1988 1899 2022
rect 1647 1954 1899 1988
rect 1647 1920 1648 1954
rect 1682 1920 1720 1954
rect 1754 1920 1792 1954
rect 1826 1920 1864 1954
rect 1898 1920 1899 1954
rect 1647 1886 1899 1920
rect 1647 1852 1648 1886
rect 1682 1852 1720 1886
rect 1754 1852 1792 1886
rect 1826 1852 1864 1886
rect 1898 1852 1899 1886
rect 1647 1818 1899 1852
rect 1647 1784 1648 1818
rect 1682 1784 1720 1818
rect 1754 1784 1792 1818
rect 1826 1784 1864 1818
rect 1898 1784 1899 1818
rect 1647 1750 1899 1784
rect 1647 1716 1648 1750
rect 1682 1716 1720 1750
rect 1754 1716 1792 1750
rect 1826 1716 1864 1750
rect 1898 1716 1899 1750
rect 1647 1682 1899 1716
rect 1647 1648 1648 1682
rect 1682 1648 1720 1682
rect 1754 1648 1792 1682
rect 1826 1648 1864 1682
rect 1898 1648 1899 1682
rect 1647 1614 1899 1648
rect 1647 1580 1648 1614
rect 1682 1580 1720 1614
rect 1754 1580 1792 1614
rect 1826 1580 1864 1614
rect 1898 1580 1899 1614
rect 1647 1546 1899 1580
rect 1647 1512 1648 1546
rect 1682 1512 1720 1546
rect 1754 1512 1792 1546
rect 1826 1512 1864 1546
rect 1898 1512 1899 1546
rect 1647 1478 1899 1512
rect 1647 1444 1648 1478
rect 1682 1444 1720 1478
rect 1754 1444 1792 1478
rect 1826 1444 1864 1478
rect 1898 1444 1899 1478
rect 1647 1410 1899 1444
rect 1647 1376 1648 1410
rect 1682 1376 1720 1410
rect 1754 1376 1792 1410
rect 1826 1376 1864 1410
rect 1898 1376 1899 1410
rect 1647 1342 1899 1376
rect 1647 1308 1648 1342
rect 1682 1308 1720 1342
rect 1754 1308 1792 1342
rect 1826 1308 1864 1342
rect 1898 1308 1899 1342
rect 1647 1274 1899 1308
rect 1647 1240 1648 1274
rect 1682 1240 1720 1274
rect 1754 1240 1792 1274
rect 1826 1240 1864 1274
rect 1898 1240 1899 1274
rect 1647 1206 1899 1240
rect 1647 1172 1648 1206
rect 1682 1172 1720 1206
rect 1754 1172 1792 1206
rect 1826 1172 1864 1206
rect 1898 1172 1899 1206
rect 1647 1138 1899 1172
rect 1647 1104 1648 1138
rect 1682 1104 1720 1138
rect 1754 1104 1792 1138
rect 1826 1104 1864 1138
rect 1898 1104 1899 1138
rect 1647 1070 1899 1104
rect 1647 1036 1648 1070
rect 1682 1036 1720 1070
rect 1754 1036 1792 1070
rect 1826 1036 1864 1070
rect 1898 1036 1899 1070
rect 1647 1002 1899 1036
rect 1647 968 1648 1002
rect 1682 968 1720 1002
rect 1754 968 1792 1002
rect 1826 968 1864 1002
rect 1898 968 1899 1002
rect 1647 934 1899 968
rect 1647 900 1648 934
rect 1682 900 1720 934
rect 1754 900 1792 934
rect 1826 900 1864 934
rect 1898 900 1899 934
rect 1647 866 1899 900
rect 1647 832 1648 866
rect 1682 832 1720 866
rect 1754 832 1792 866
rect 1826 832 1864 866
rect 1898 832 1899 866
rect 1647 798 1899 832
rect 1647 764 1648 798
rect 1682 764 1720 798
rect 1754 764 1792 798
rect 1826 764 1864 798
rect 1898 764 1899 798
rect 1647 730 1899 764
rect 1647 696 1648 730
rect 1682 696 1720 730
rect 1754 696 1792 730
rect 1826 696 1864 730
rect 1898 696 1899 730
rect 1647 662 1899 696
rect 1647 628 1648 662
rect 1682 628 1720 662
rect 1754 628 1792 662
rect 1826 628 1864 662
rect 1898 628 1899 662
rect 1647 594 1899 628
rect 1647 560 1648 594
rect 1682 560 1720 594
rect 1754 560 1792 594
rect 1826 560 1864 594
rect 1898 560 1899 594
rect 1647 526 1899 560
rect 1647 492 1648 526
rect 1682 492 1720 526
rect 1754 492 1792 526
rect 1826 492 1864 526
rect 1898 492 1899 526
rect 1647 458 1899 492
rect 1647 447 1648 458
rect 1682 447 1720 458
rect 1754 447 1792 458
rect 1826 447 1864 458
rect 1898 447 1899 458
rect 4005 2039 4139 2073
rect 4173 2039 4207 2073
rect 4241 2039 4275 2073
rect 4309 2039 4343 2073
rect 4377 2039 4411 2073
rect 4445 2039 4479 2073
rect 4513 2039 4547 2073
rect 4581 2039 4615 2073
rect 4649 2039 4683 2073
rect 4717 2039 4751 2073
rect 4785 2039 4819 2073
rect 4853 2039 4887 2073
rect 4921 2039 4955 2073
rect 4989 2039 5023 2073
rect 5057 2039 5091 2073
rect 5125 2039 5159 2073
rect 5193 2039 5227 2073
rect 5261 2039 5295 2073
rect 5329 2039 5363 2073
rect 5397 2039 5431 2073
rect 5465 2039 5499 2073
rect 5533 2039 5567 2073
rect 5601 2039 5635 2073
rect 5669 2039 5703 2073
rect 5737 2039 5771 2073
rect 5805 2039 5839 2073
rect 5873 2039 5907 2073
rect 5941 2039 5975 2073
rect 6009 2039 6043 2073
rect 6077 2039 6111 2073
rect 6145 2039 6179 2073
rect 6213 2039 6247 2073
rect 6281 2039 6315 2073
rect 6349 2039 6383 2073
rect 6417 2039 6451 2073
rect 6485 2039 6519 2073
rect 6553 2039 6587 2073
rect 6621 2039 6689 2073
rect 4005 2005 4039 2039
rect 6655 1999 6689 2039
rect 4005 1937 4039 1971
rect 4005 1869 4039 1903
rect 6655 1931 6689 1965
rect 4005 1801 4039 1835
rect 4005 1733 4039 1767
rect 4005 1665 4039 1699
rect 4005 1597 4039 1631
rect 4005 1529 4039 1563
rect 4005 1461 4039 1495
rect 4005 1393 4039 1427
rect 4005 1325 4039 1359
rect 4005 1257 4039 1291
rect 4005 1189 4039 1223
rect 4005 1121 4039 1155
rect 4005 1053 4039 1087
rect 4005 985 4039 1019
rect 4005 917 4039 951
rect 4005 849 4039 883
rect 4005 781 4039 815
rect 4005 713 4039 747
rect 4005 645 4039 679
rect 4005 486 4039 611
rect 6655 1863 6689 1897
rect 6655 1795 6689 1829
rect 6655 1727 6689 1761
rect 6655 1659 6689 1693
rect 6655 1591 6689 1625
rect 6655 1523 6689 1557
rect 6655 1455 6689 1489
rect 6655 1387 6689 1421
rect 6655 1319 6689 1353
rect 6655 1251 6689 1285
rect 6655 1183 6689 1217
rect 6655 1115 6689 1149
rect 6655 1047 6689 1081
rect 6655 979 6689 1013
rect 6655 911 6689 945
rect 6655 843 6689 877
rect 6655 775 6689 809
rect 6655 707 6689 741
rect 6655 639 6689 673
rect 6655 571 6689 605
rect 6655 503 6689 537
rect 4005 447 4039 452
rect 6655 447 6689 469
rect 7097 2073 7175 2107
rect 7209 2073 7243 2107
rect 7277 2073 7311 2107
rect 7345 2073 7379 2107
rect 7413 2073 7447 2107
rect 7481 2073 7515 2107
rect 7549 2073 7583 2107
rect 7617 2073 7651 2107
rect 7685 2073 7719 2107
rect 7753 2073 7787 2107
rect 7821 2073 7855 2107
rect 7889 2073 7923 2107
rect 7957 2073 7991 2107
rect 8025 2073 8059 2107
rect 8093 2073 8127 2107
rect 8161 2073 8195 2107
rect 8229 2073 8263 2107
rect 8297 2073 8331 2107
rect 8365 2073 8399 2107
rect 8433 2073 8467 2107
rect 8501 2073 8535 2107
rect 8569 2073 8603 2107
rect 8637 2073 8671 2107
rect 8705 2073 8739 2107
rect 8773 2073 8807 2107
rect 8841 2073 8875 2107
rect 8909 2073 8943 2107
rect 8977 2073 9011 2107
rect 9045 2073 9079 2107
rect 9113 2073 9147 2107
rect 9181 2073 9215 2107
rect 9249 2073 9283 2107
rect 9317 2073 9351 2107
rect 9385 2073 9419 2107
rect 9453 2073 9487 2107
rect 9521 2073 9555 2107
rect 9589 2073 9623 2107
rect 9657 2073 9691 2107
rect 9725 2073 9759 2107
rect 9793 2073 9827 2107
rect 9861 2073 9895 2107
rect 9929 2073 9997 2107
rect 7097 2039 7131 2073
rect 7097 1971 7131 2005
rect 9963 2033 9997 2073
rect 9963 1965 9997 1999
rect 7097 1903 7131 1937
rect 7097 1835 7131 1869
rect 7097 1767 7131 1801
rect 7097 1699 7131 1733
rect 7097 1631 7131 1665
rect 7097 1563 7131 1597
rect 7097 1495 7131 1529
rect 7097 1427 7131 1461
rect 7097 1359 7131 1393
rect 7097 1291 7131 1325
rect 7097 1223 7131 1257
rect 7097 1155 7131 1189
rect 7097 1087 7131 1121
rect 7097 1019 7131 1053
rect 7097 951 7131 985
rect 7097 883 7131 917
rect 7097 815 7131 849
rect 7097 747 7131 781
rect 7097 679 7131 713
rect 7097 554 7131 645
rect 9963 1897 9997 1931
rect 9963 1829 9997 1863
rect 9963 1761 9997 1795
rect 9963 1693 9997 1727
rect 9963 1625 9997 1659
rect 9963 1557 9997 1591
rect 9963 1489 9997 1523
rect 9963 1421 9997 1455
rect 9963 1353 9997 1387
rect 9963 1285 9997 1319
rect 9963 1217 9997 1251
rect 9963 1149 9997 1183
rect 9963 1081 9997 1115
rect 9963 1013 9997 1047
rect 9963 945 9997 979
rect 9963 877 9997 911
rect 9963 809 9997 843
rect 9963 741 9997 775
rect 9963 673 9997 707
rect 9963 605 9997 639
rect 7097 469 7131 520
rect 9963 537 9997 571
rect 9963 469 9997 503
rect 7097 447 7165 469
rect 7199 447 7233 469
rect 7267 447 7301 469
rect 7335 447 7369 469
rect 7403 447 7437 469
rect 7471 447 7505 469
rect 7539 447 7573 469
rect 7607 447 7641 469
rect 7675 447 7709 469
rect 7743 447 7777 469
rect 7811 447 7845 469
rect 7879 447 7913 469
rect 7947 447 7981 469
rect 8015 447 8049 469
rect 8083 447 8117 469
rect 8151 447 8185 469
rect 8219 447 8253 469
rect 8287 447 8321 469
rect 8355 447 8389 469
rect 8423 447 8457 469
rect 8491 447 8525 469
rect 8559 447 8593 469
rect 8627 447 8661 469
rect 8695 447 8729 469
rect 8763 447 8797 469
rect 8831 447 8865 469
rect 8899 447 8933 469
rect 8967 447 9001 469
rect 9035 447 9069 469
rect 9103 447 9137 469
rect 9171 447 9205 469
rect 9239 447 9273 469
rect 9307 447 9341 469
rect 9375 447 9409 469
rect 9443 447 9477 469
rect 9511 447 9545 469
rect 9579 447 9613 469
rect 9647 447 9681 469
rect 9715 447 9749 469
rect 9783 447 9817 469
rect 9851 447 9885 469
rect 9919 447 9997 469
<< mvnsubdiff >>
rect 237 2057 371 2091
rect 405 2057 439 2091
rect 473 2057 507 2091
rect 541 2057 575 2091
rect 609 2057 643 2091
rect 677 2057 711 2091
rect 745 2057 779 2091
rect 813 2057 847 2091
rect 881 2057 915 2091
rect 949 2057 983 2091
rect 1017 2057 1051 2091
rect 1085 2057 1119 2091
rect 1153 2057 1187 2091
rect 1221 2057 1255 2091
rect 1289 2057 1323 2091
rect 1357 2057 1391 2091
rect 1425 2057 1493 2091
rect 237 2023 271 2057
rect 237 1955 271 1989
rect 237 1887 271 1921
rect 1459 1959 1493 2057
rect 1459 1891 1493 1925
rect 237 1819 271 1853
rect 237 1751 271 1785
rect 237 1683 271 1717
rect 237 1615 271 1649
rect 237 1547 271 1581
rect 237 1479 271 1513
rect 237 1411 271 1445
rect 237 1343 271 1377
rect 237 1275 271 1309
rect 237 1123 271 1241
rect 237 1055 271 1089
rect 237 987 271 1021
rect 237 919 271 953
rect 237 851 271 885
rect 237 783 271 817
rect 237 715 271 749
rect 237 647 271 681
rect 237 579 271 613
rect 237 511 271 545
rect 237 447 271 477
rect 1459 1823 1493 1857
rect 1459 1755 1493 1789
rect 1459 1687 1493 1721
rect 1459 1619 1493 1653
rect 1459 1551 1493 1585
rect 1459 1483 1493 1517
rect 1459 1415 1493 1449
rect 1459 1347 1493 1381
rect 1459 1279 1493 1313
rect 1459 1211 1493 1245
rect 1459 1143 1493 1177
rect 1459 1075 1493 1109
rect 1459 1007 1493 1041
rect 1459 939 1493 973
rect 1459 871 1493 905
rect 1459 803 1493 837
rect 1459 735 1493 769
rect 1459 667 1493 701
rect 1459 599 1493 633
rect 1459 531 1493 565
rect 1459 463 1493 497
rect 2052 2025 2120 2107
rect 2086 2005 2120 2025
rect 3106 2073 3140 2107
rect 3174 2073 3282 2107
rect 3106 2039 3282 2073
rect 3106 2005 3180 2039
rect 2086 1991 2154 2005
rect 2052 1957 2154 1991
rect 3180 910 3282 985
rect 3180 447 3282 468
rect 3750 2260 3818 2362
rect 10108 2294 10262 2362
rect 10108 2274 10228 2294
rect 10108 2260 10160 2274
rect 3750 2254 3852 2260
rect 3784 2220 3852 2254
rect 3750 2186 3852 2220
rect 3750 447 3852 452
rect 6842 661 6944 696
rect 6876 627 6910 661
rect 6842 592 6944 627
rect 6876 558 6910 592
rect 6842 523 6944 558
rect 6876 489 6910 523
rect 6842 454 6944 489
rect 6876 420 6910 454
rect 10160 458 10262 472
rect 10160 447 10228 458
rect 6842 385 6944 420
rect 6876 351 6910 385
rect 6842 316 6944 351
rect 6876 282 6910 316
rect 6842 248 6944 282
rect 6876 214 6964 248
rect 6998 214 7010 248
rect 6842 182 7010 214
<< psubdiffcont >>
rect -24 211 78 447
rect 1648 424 1682 447
rect 1720 424 1754 447
rect 1792 424 1826 447
rect 1864 424 1898 447
rect -24 143 10 177
rect 1648 356 1682 390
rect 1720 356 1754 390
rect 1792 356 1826 390
rect 1864 356 1898 390
rect 1648 288 1682 322
rect 1720 288 1754 322
rect 1792 288 1826 322
rect 1864 288 1898 322
rect 1648 220 1682 254
rect 1720 220 1754 254
rect 1792 220 1826 254
rect 1864 220 1898 254
rect 44 36 3342 138
rect 3435 104 3537 447
rect 3376 36 3410 70
rect 6655 401 6689 435
rect 4073 333 4107 367
rect 4141 333 4175 367
rect 4209 333 4243 367
rect 4277 333 4311 367
rect 4345 333 4379 367
rect 4413 333 4447 367
rect 4481 333 4515 367
rect 4549 333 4583 367
rect 4617 333 4651 367
rect 4685 333 4719 367
rect 4753 333 4787 367
rect 4821 333 4855 367
rect 4889 333 4923 367
rect 4957 333 4991 367
rect 5025 333 5059 367
rect 5093 333 5127 367
rect 5161 333 5195 367
rect 5229 333 5263 367
rect 5297 333 5331 367
rect 5365 333 5399 367
rect 5433 333 5467 367
rect 5501 333 5535 367
rect 5569 333 5603 367
rect 5637 333 5671 367
rect 5705 333 5739 367
rect 5773 333 5807 367
rect 5841 333 5875 367
rect 5909 333 5943 367
rect 5977 333 6011 367
rect 6045 333 6079 367
rect 6113 333 6147 367
rect 6181 333 6215 367
rect 6249 333 6283 367
rect 6317 333 6351 367
rect 6385 333 6419 367
rect 6453 333 6487 367
rect 6521 333 6555 367
rect 7165 435 7199 447
rect 7233 435 7267 447
rect 7301 435 7335 447
rect 7369 435 7403 447
rect 7437 435 7471 447
rect 7505 435 7539 447
rect 7573 435 7607 447
rect 7641 435 7675 447
rect 7709 435 7743 447
rect 7777 435 7811 447
rect 7845 435 7879 447
rect 7913 435 7947 447
rect 7981 435 8015 447
rect 8049 435 8083 447
rect 8117 435 8151 447
rect 8185 435 8219 447
rect 8253 435 8287 447
rect 8321 435 8355 447
rect 8389 435 8423 447
rect 8457 435 8491 447
rect 8525 435 8559 447
rect 8593 435 8627 447
rect 8661 435 8695 447
rect 8729 435 8763 447
rect 8797 435 8831 447
rect 8865 435 8899 447
rect 8933 435 8967 447
rect 9001 435 9035 447
rect 9069 435 9103 447
rect 9137 435 9171 447
rect 9205 435 9239 447
rect 9273 435 9307 447
rect 9341 435 9375 447
rect 9409 435 9443 447
rect 9477 435 9511 447
rect 9545 435 9579 447
rect 9613 435 9647 447
rect 9681 435 9715 447
rect 9749 435 9783 447
rect 9817 435 9851 447
rect 9885 435 9919 447
<< nsubdiffcont >>
rect 1459 429 1493 447
rect 305 361 339 395
rect 373 361 407 395
rect 441 361 475 395
rect 509 361 543 395
rect 577 361 611 395
rect 645 361 679 395
rect 713 361 747 395
rect 781 361 815 395
rect 849 361 883 395
rect 917 361 951 395
rect 985 361 1019 395
rect 1053 361 1087 395
rect 1121 361 1155 395
rect 1189 361 1223 395
rect 1257 361 1291 395
rect 1325 361 1359 395
rect 2052 359 2154 447
rect 3248 400 3282 434
rect 2160 291 2194 325
rect 2228 291 3214 393
rect 3750 112 3852 418
rect 10228 438 10262 447
rect 10160 336 10262 438
rect 10228 288 10262 322
rect 6910 146 6944 180
rect 7032 146 10194 248
rect 10228 220 10262 254
rect 3850 44 3884 78
rect 3918 44 6876 146
<< mvpsubdiffcont >>
rect 69 2260 3503 2362
rect -24 1376 78 2226
rect 1648 2192 1682 2226
rect 1720 2192 1754 2226
rect 1792 2192 1826 2226
rect 1864 2192 1898 2226
rect 1648 2124 1682 2158
rect 1720 2124 1754 2158
rect 1792 2124 1826 2158
rect 1864 2124 1898 2158
rect -24 447 78 1265
rect 1648 2056 1682 2090
rect 1720 2056 1754 2090
rect 1792 2056 1826 2090
rect 1864 2056 1898 2090
rect 1648 1988 1682 2022
rect 1720 1988 1754 2022
rect 1792 1988 1826 2022
rect 1864 1988 1898 2022
rect 1648 1920 1682 1954
rect 1720 1920 1754 1954
rect 1792 1920 1826 1954
rect 1864 1920 1898 1954
rect 1648 1852 1682 1886
rect 1720 1852 1754 1886
rect 1792 1852 1826 1886
rect 1864 1852 1898 1886
rect 1648 1784 1682 1818
rect 1720 1784 1754 1818
rect 1792 1784 1826 1818
rect 1864 1784 1898 1818
rect 1648 1716 1682 1750
rect 1720 1716 1754 1750
rect 1792 1716 1826 1750
rect 1864 1716 1898 1750
rect 1648 1648 1682 1682
rect 1720 1648 1754 1682
rect 1792 1648 1826 1682
rect 1864 1648 1898 1682
rect 1648 1580 1682 1614
rect 1720 1580 1754 1614
rect 1792 1580 1826 1614
rect 1864 1580 1898 1614
rect 1648 1512 1682 1546
rect 1720 1512 1754 1546
rect 1792 1512 1826 1546
rect 1864 1512 1898 1546
rect 1648 1444 1682 1478
rect 1720 1444 1754 1478
rect 1792 1444 1826 1478
rect 1864 1444 1898 1478
rect 1648 1376 1682 1410
rect 1720 1376 1754 1410
rect 1792 1376 1826 1410
rect 1864 1376 1898 1410
rect 1648 1308 1682 1342
rect 1720 1308 1754 1342
rect 1792 1308 1826 1342
rect 1864 1308 1898 1342
rect 1648 1240 1682 1274
rect 1720 1240 1754 1274
rect 1792 1240 1826 1274
rect 1864 1240 1898 1274
rect 1648 1172 1682 1206
rect 1720 1172 1754 1206
rect 1792 1172 1826 1206
rect 1864 1172 1898 1206
rect 1648 1104 1682 1138
rect 1720 1104 1754 1138
rect 1792 1104 1826 1138
rect 1864 1104 1898 1138
rect 1648 1036 1682 1070
rect 1720 1036 1754 1070
rect 1792 1036 1826 1070
rect 1864 1036 1898 1070
rect 1648 968 1682 1002
rect 1720 968 1754 1002
rect 1792 968 1826 1002
rect 1864 968 1898 1002
rect 1648 900 1682 934
rect 1720 900 1754 934
rect 1792 900 1826 934
rect 1864 900 1898 934
rect 1648 832 1682 866
rect 1720 832 1754 866
rect 1792 832 1826 866
rect 1864 832 1898 866
rect 1648 764 1682 798
rect 1720 764 1754 798
rect 1792 764 1826 798
rect 1864 764 1898 798
rect 1648 696 1682 730
rect 1720 696 1754 730
rect 1792 696 1826 730
rect 1864 696 1898 730
rect 1648 628 1682 662
rect 1720 628 1754 662
rect 1792 628 1826 662
rect 1864 628 1898 662
rect 1648 560 1682 594
rect 1720 560 1754 594
rect 1792 560 1826 594
rect 1864 560 1898 594
rect 1648 492 1682 526
rect 1720 492 1754 526
rect 1792 492 1826 526
rect 1864 492 1898 526
rect 1648 447 1682 458
rect 1720 447 1754 458
rect 1792 447 1826 458
rect 1864 447 1898 458
rect 3435 447 3537 2178
rect 4139 2039 4173 2073
rect 4207 2039 4241 2073
rect 4275 2039 4309 2073
rect 4343 2039 4377 2073
rect 4411 2039 4445 2073
rect 4479 2039 4513 2073
rect 4547 2039 4581 2073
rect 4615 2039 4649 2073
rect 4683 2039 4717 2073
rect 4751 2039 4785 2073
rect 4819 2039 4853 2073
rect 4887 2039 4921 2073
rect 4955 2039 4989 2073
rect 5023 2039 5057 2073
rect 5091 2039 5125 2073
rect 5159 2039 5193 2073
rect 5227 2039 5261 2073
rect 5295 2039 5329 2073
rect 5363 2039 5397 2073
rect 5431 2039 5465 2073
rect 5499 2039 5533 2073
rect 5567 2039 5601 2073
rect 5635 2039 5669 2073
rect 5703 2039 5737 2073
rect 5771 2039 5805 2073
rect 5839 2039 5873 2073
rect 5907 2039 5941 2073
rect 5975 2039 6009 2073
rect 6043 2039 6077 2073
rect 6111 2039 6145 2073
rect 6179 2039 6213 2073
rect 6247 2039 6281 2073
rect 6315 2039 6349 2073
rect 6383 2039 6417 2073
rect 6451 2039 6485 2073
rect 6519 2039 6553 2073
rect 6587 2039 6621 2073
rect 4005 1971 4039 2005
rect 4005 1903 4039 1937
rect 6655 1965 6689 1999
rect 6655 1897 6689 1931
rect 4005 1835 4039 1869
rect 4005 1767 4039 1801
rect 4005 1699 4039 1733
rect 4005 1631 4039 1665
rect 4005 1563 4039 1597
rect 4005 1495 4039 1529
rect 4005 1427 4039 1461
rect 4005 1359 4039 1393
rect 4005 1291 4039 1325
rect 4005 1223 4039 1257
rect 4005 1155 4039 1189
rect 4005 1087 4039 1121
rect 4005 1019 4039 1053
rect 4005 951 4039 985
rect 4005 883 4039 917
rect 4005 815 4039 849
rect 4005 747 4039 781
rect 4005 679 4039 713
rect 4005 611 4039 645
rect 4005 452 4039 486
rect 6655 1829 6689 1863
rect 6655 1761 6689 1795
rect 6655 1693 6689 1727
rect 6655 1625 6689 1659
rect 6655 1557 6689 1591
rect 6655 1489 6689 1523
rect 6655 1421 6689 1455
rect 6655 1353 6689 1387
rect 6655 1285 6689 1319
rect 6655 1217 6689 1251
rect 6655 1149 6689 1183
rect 6655 1081 6689 1115
rect 6655 1013 6689 1047
rect 6655 945 6689 979
rect 6655 877 6689 911
rect 6655 809 6689 843
rect 6655 741 6689 775
rect 6655 673 6689 707
rect 6655 605 6689 639
rect 6655 537 6689 571
rect 6655 469 6689 503
rect 7175 2073 7209 2107
rect 7243 2073 7277 2107
rect 7311 2073 7345 2107
rect 7379 2073 7413 2107
rect 7447 2073 7481 2107
rect 7515 2073 7549 2107
rect 7583 2073 7617 2107
rect 7651 2073 7685 2107
rect 7719 2073 7753 2107
rect 7787 2073 7821 2107
rect 7855 2073 7889 2107
rect 7923 2073 7957 2107
rect 7991 2073 8025 2107
rect 8059 2073 8093 2107
rect 8127 2073 8161 2107
rect 8195 2073 8229 2107
rect 8263 2073 8297 2107
rect 8331 2073 8365 2107
rect 8399 2073 8433 2107
rect 8467 2073 8501 2107
rect 8535 2073 8569 2107
rect 8603 2073 8637 2107
rect 8671 2073 8705 2107
rect 8739 2073 8773 2107
rect 8807 2073 8841 2107
rect 8875 2073 8909 2107
rect 8943 2073 8977 2107
rect 9011 2073 9045 2107
rect 9079 2073 9113 2107
rect 9147 2073 9181 2107
rect 9215 2073 9249 2107
rect 9283 2073 9317 2107
rect 9351 2073 9385 2107
rect 9419 2073 9453 2107
rect 9487 2073 9521 2107
rect 9555 2073 9589 2107
rect 9623 2073 9657 2107
rect 9691 2073 9725 2107
rect 9759 2073 9793 2107
rect 9827 2073 9861 2107
rect 9895 2073 9929 2107
rect 7097 2005 7131 2039
rect 7097 1937 7131 1971
rect 9963 1999 9997 2033
rect 7097 1869 7131 1903
rect 7097 1801 7131 1835
rect 7097 1733 7131 1767
rect 7097 1665 7131 1699
rect 7097 1597 7131 1631
rect 7097 1529 7131 1563
rect 7097 1461 7131 1495
rect 7097 1393 7131 1427
rect 7097 1325 7131 1359
rect 7097 1257 7131 1291
rect 7097 1189 7131 1223
rect 7097 1121 7131 1155
rect 7097 1053 7131 1087
rect 7097 985 7131 1019
rect 7097 917 7131 951
rect 7097 849 7131 883
rect 7097 781 7131 815
rect 7097 713 7131 747
rect 7097 645 7131 679
rect 7097 520 7131 554
rect 9963 1931 9997 1965
rect 9963 1863 9997 1897
rect 9963 1795 9997 1829
rect 9963 1727 9997 1761
rect 9963 1659 9997 1693
rect 9963 1591 9997 1625
rect 9963 1523 9997 1557
rect 9963 1455 9997 1489
rect 9963 1387 9997 1421
rect 9963 1319 9997 1353
rect 9963 1251 9997 1285
rect 9963 1183 9997 1217
rect 9963 1115 9997 1149
rect 9963 1047 9997 1081
rect 9963 979 9997 1013
rect 9963 911 9997 945
rect 9963 843 9997 877
rect 9963 775 9997 809
rect 9963 707 9997 741
rect 9963 639 9997 673
rect 9963 571 9997 605
rect 9963 503 9997 537
rect 7165 447 7199 469
rect 7233 447 7267 469
rect 7301 447 7335 469
rect 7369 447 7403 469
rect 7437 447 7471 469
rect 7505 447 7539 469
rect 7573 447 7607 469
rect 7641 447 7675 469
rect 7709 447 7743 469
rect 7777 447 7811 469
rect 7845 447 7879 469
rect 7913 447 7947 469
rect 7981 447 8015 469
rect 8049 447 8083 469
rect 8117 447 8151 469
rect 8185 447 8219 469
rect 8253 447 8287 469
rect 8321 447 8355 469
rect 8389 447 8423 469
rect 8457 447 8491 469
rect 8525 447 8559 469
rect 8593 447 8627 469
rect 8661 447 8695 469
rect 8729 447 8763 469
rect 8797 447 8831 469
rect 8865 447 8899 469
rect 8933 447 8967 469
rect 9001 447 9035 469
rect 9069 447 9103 469
rect 9137 447 9171 469
rect 9205 447 9239 469
rect 9273 447 9307 469
rect 9341 447 9375 469
rect 9409 447 9443 469
rect 9477 447 9511 469
rect 9545 447 9579 469
rect 9613 447 9647 469
rect 9681 447 9715 469
rect 9749 447 9783 469
rect 9817 447 9851 469
rect 9885 447 9919 469
<< mvnsubdiffcont >>
rect 371 2057 405 2091
rect 439 2057 473 2091
rect 507 2057 541 2091
rect 575 2057 609 2091
rect 643 2057 677 2091
rect 711 2057 745 2091
rect 779 2057 813 2091
rect 847 2057 881 2091
rect 915 2057 949 2091
rect 983 2057 1017 2091
rect 1051 2057 1085 2091
rect 1119 2057 1153 2091
rect 1187 2057 1221 2091
rect 1255 2057 1289 2091
rect 1323 2057 1357 2091
rect 1391 2057 1425 2091
rect 237 1989 271 2023
rect 237 1921 271 1955
rect 237 1853 271 1887
rect 1459 1925 1493 1959
rect 237 1785 271 1819
rect 237 1717 271 1751
rect 237 1649 271 1683
rect 237 1581 271 1615
rect 237 1513 271 1547
rect 237 1445 271 1479
rect 237 1377 271 1411
rect 237 1309 271 1343
rect 237 1241 271 1275
rect 237 1089 271 1123
rect 237 1021 271 1055
rect 237 953 271 987
rect 237 885 271 919
rect 237 817 271 851
rect 237 749 271 783
rect 237 681 271 715
rect 237 613 271 647
rect 237 545 271 579
rect 237 477 271 511
rect 1459 1857 1493 1891
rect 1459 1789 1493 1823
rect 1459 1721 1493 1755
rect 1459 1653 1493 1687
rect 1459 1585 1493 1619
rect 1459 1517 1493 1551
rect 1459 1449 1493 1483
rect 1459 1381 1493 1415
rect 1459 1313 1493 1347
rect 1459 1245 1493 1279
rect 1459 1177 1493 1211
rect 1459 1109 1493 1143
rect 1459 1041 1493 1075
rect 1459 973 1493 1007
rect 1459 905 1493 939
rect 1459 837 1493 871
rect 1459 769 1493 803
rect 1459 701 1493 735
rect 1459 633 1493 667
rect 1459 565 1493 599
rect 1459 497 1493 531
rect 1459 447 1493 463
rect 2052 1991 2086 2025
rect 2120 2005 3106 2107
rect 3140 2073 3174 2107
rect 2052 447 2154 1957
rect 3180 985 3282 2039
rect 3180 468 3282 910
rect 3818 2260 10108 2362
rect 10228 2274 10262 2294
rect 3750 2220 3784 2254
rect 3750 452 3852 2186
rect 6842 696 6944 2260
rect 6842 627 6876 661
rect 6910 627 6944 661
rect 6842 558 6876 592
rect 6910 558 6944 592
rect 6842 489 6876 523
rect 6910 489 6944 523
rect 6842 420 6876 454
rect 6910 420 6944 454
rect 10160 472 10262 2274
rect 10228 447 10262 458
rect 6842 351 6876 385
rect 6910 351 6944 385
rect 6842 282 6876 316
rect 6910 282 6944 316
rect 6842 214 6876 248
rect 6964 214 6998 248
<< poly >>
rect 414 1957 1322 1973
rect 414 1923 430 1957
rect 464 1923 501 1957
rect 535 1923 572 1957
rect 606 1923 642 1957
rect 676 1923 712 1957
rect 746 1923 782 1957
rect 816 1923 852 1957
rect 886 1923 922 1957
rect 956 1923 992 1957
rect 1026 1923 1062 1957
rect 1096 1923 1132 1957
rect 1166 1923 1202 1957
rect 1236 1923 1272 1957
rect 1306 1923 1322 1957
rect 414 1907 1322 1923
rect 414 1875 514 1907
rect 570 1875 670 1907
rect 740 1875 840 1907
rect 896 1875 996 1907
rect 1066 1875 1166 1907
rect 1222 1875 1322 1907
rect 414 443 514 475
rect 570 443 670 475
rect 740 443 840 475
rect 896 443 996 475
rect 1066 443 1166 475
rect 1222 443 1322 475
rect 2291 1957 3043 1973
rect 2291 1923 2307 1957
rect 2341 1923 2376 1957
rect 2410 1923 2445 1957
rect 2479 1923 2514 1957
rect 2548 1923 2583 1957
rect 2617 1923 2652 1957
rect 2686 1923 2721 1957
rect 2755 1923 2789 1957
rect 2823 1923 2857 1957
rect 2891 1923 2925 1957
rect 2959 1923 2993 1957
rect 3027 1923 3043 1957
rect 2291 1907 3043 1923
rect 2291 1875 2391 1907
rect 2461 1875 2561 1907
rect 2617 1875 2717 1907
rect 2787 1875 2887 1907
rect 2943 1875 3043 1907
rect 2291 443 2391 475
rect 2461 443 2561 475
rect 2617 443 2717 475
rect 2787 443 2887 475
rect 2943 443 3043 475
rect 4176 1957 5254 1973
rect 4176 1923 4192 1957
rect 4226 1923 4264 1957
rect 4298 1923 4336 1957
rect 4370 1923 4408 1957
rect 4442 1923 4480 1957
rect 4514 1923 4552 1957
rect 4586 1923 4624 1957
rect 4658 1923 4696 1957
rect 4730 1923 4768 1957
rect 4802 1923 4840 1957
rect 4874 1923 4912 1957
rect 4946 1923 4985 1957
rect 5019 1923 5058 1957
rect 5092 1923 5131 1957
rect 5165 1923 5204 1957
rect 5238 1923 5254 1957
rect 4176 1907 5254 1923
rect 4176 1875 4276 1907
rect 4346 1875 4446 1907
rect 4502 1875 4602 1907
rect 4672 1875 4772 1907
rect 4828 1875 4928 1907
rect 4998 1875 5098 1907
rect 5154 1875 5254 1907
rect 5447 1957 6525 1973
rect 5447 1923 5463 1957
rect 5497 1923 5536 1957
rect 5570 1923 5609 1957
rect 5643 1923 5682 1957
rect 5716 1923 5755 1957
rect 5789 1923 5827 1957
rect 5861 1923 5899 1957
rect 5933 1923 5971 1957
rect 6005 1923 6043 1957
rect 6077 1923 6115 1957
rect 6149 1923 6187 1957
rect 6221 1923 6259 1957
rect 6293 1923 6331 1957
rect 6365 1923 6403 1957
rect 6437 1923 6475 1957
rect 6509 1923 6525 1957
rect 5447 1907 6525 1923
rect 5447 1875 5547 1907
rect 5603 1875 5703 1907
rect 5773 1875 5873 1907
rect 5929 1875 6029 1907
rect 6099 1875 6199 1907
rect 6255 1875 6355 1907
rect 6425 1875 6525 1907
rect 4176 443 4276 475
rect 4346 443 4446 475
rect 4502 443 4602 475
rect 4672 443 4772 475
rect 4828 443 4928 475
rect 4998 443 5098 475
rect 5154 443 5254 475
rect 5447 443 5547 475
rect 5603 443 5703 475
rect 5773 443 5873 475
rect 5929 443 6029 475
rect 6099 443 6199 475
rect 6255 443 6355 475
rect 6425 443 6525 475
rect 7261 2025 8339 2041
rect 7261 1991 7277 2025
rect 7311 1991 7350 2025
rect 7384 1991 7423 2025
rect 7457 1991 7496 2025
rect 7530 1991 7569 2025
rect 7603 1991 7641 2025
rect 7675 1991 7713 2025
rect 7747 1991 7785 2025
rect 7819 1991 7857 2025
rect 7891 1991 7929 2025
rect 7963 1991 8001 2025
rect 8035 1991 8073 2025
rect 8107 1991 8145 2025
rect 8179 1991 8217 2025
rect 8251 1991 8289 2025
rect 8323 1991 8339 2025
rect 7261 1975 8339 1991
rect 7261 1943 7361 1975
rect 7431 1943 7531 1975
rect 7587 1943 7687 1975
rect 7757 1943 7857 1975
rect 7913 1943 8013 1975
rect 8083 1943 8183 1975
rect 8239 1943 8339 1975
rect 8532 2025 9766 2041
rect 8532 1991 8548 2025
rect 8582 1991 8617 2025
rect 8651 1991 8686 2025
rect 8720 1991 8755 2025
rect 8789 1991 8824 2025
rect 8858 1991 8893 2025
rect 8927 1991 8962 2025
rect 8996 1991 9031 2025
rect 9065 1991 9100 2025
rect 9134 1991 9169 2025
rect 9203 1991 9238 2025
rect 9272 1991 9307 2025
rect 9341 1991 9376 2025
rect 9410 1991 9444 2025
rect 9478 1991 9512 2025
rect 9546 1991 9580 2025
rect 9614 1991 9648 2025
rect 9682 1991 9716 2025
rect 9750 1991 9766 2025
rect 8532 1975 9766 1991
rect 8532 1943 8632 1975
rect 8688 1943 8788 1975
rect 8858 1943 8958 1975
rect 9014 1943 9114 1975
rect 9184 1943 9284 1975
rect 9340 1943 9440 1975
rect 9510 1943 9610 1975
rect 9666 1943 9766 1975
rect 7261 511 7361 543
rect 7431 511 7531 543
rect 7587 511 7687 543
rect 7757 511 7857 543
rect 7913 511 8013 543
rect 8083 511 8183 543
rect 8239 511 8339 543
rect 8532 511 8632 543
rect 8688 511 8788 543
rect 8858 511 8958 543
rect 9014 511 9114 543
rect 9184 511 9284 543
rect 9340 511 9440 543
rect 9510 511 9610 543
rect 9666 511 9766 543
<< polycont >>
rect 430 1923 464 1957
rect 501 1923 535 1957
rect 572 1923 606 1957
rect 642 1923 676 1957
rect 712 1923 746 1957
rect 782 1923 816 1957
rect 852 1923 886 1957
rect 922 1923 956 1957
rect 992 1923 1026 1957
rect 1062 1923 1096 1957
rect 1132 1923 1166 1957
rect 1202 1923 1236 1957
rect 1272 1923 1306 1957
rect 2307 1923 2341 1957
rect 2376 1923 2410 1957
rect 2445 1923 2479 1957
rect 2514 1923 2548 1957
rect 2583 1923 2617 1957
rect 2652 1923 2686 1957
rect 2721 1923 2755 1957
rect 2789 1923 2823 1957
rect 2857 1923 2891 1957
rect 2925 1923 2959 1957
rect 2993 1923 3027 1957
rect 4192 1923 4226 1957
rect 4264 1923 4298 1957
rect 4336 1923 4370 1957
rect 4408 1923 4442 1957
rect 4480 1923 4514 1957
rect 4552 1923 4586 1957
rect 4624 1923 4658 1957
rect 4696 1923 4730 1957
rect 4768 1923 4802 1957
rect 4840 1923 4874 1957
rect 4912 1923 4946 1957
rect 4985 1923 5019 1957
rect 5058 1923 5092 1957
rect 5131 1923 5165 1957
rect 5204 1923 5238 1957
rect 5463 1923 5497 1957
rect 5536 1923 5570 1957
rect 5609 1923 5643 1957
rect 5682 1923 5716 1957
rect 5755 1923 5789 1957
rect 5827 1923 5861 1957
rect 5899 1923 5933 1957
rect 5971 1923 6005 1957
rect 6043 1923 6077 1957
rect 6115 1923 6149 1957
rect 6187 1923 6221 1957
rect 6259 1923 6293 1957
rect 6331 1923 6365 1957
rect 6403 1923 6437 1957
rect 6475 1923 6509 1957
rect 7277 1991 7311 2025
rect 7350 1991 7384 2025
rect 7423 1991 7457 2025
rect 7496 1991 7530 2025
rect 7569 1991 7603 2025
rect 7641 1991 7675 2025
rect 7713 1991 7747 2025
rect 7785 1991 7819 2025
rect 7857 1991 7891 2025
rect 7929 1991 7963 2025
rect 8001 1991 8035 2025
rect 8073 1991 8107 2025
rect 8145 1991 8179 2025
rect 8217 1991 8251 2025
rect 8289 1991 8323 2025
rect 8548 1991 8582 2025
rect 8617 1991 8651 2025
rect 8686 1991 8720 2025
rect 8755 1991 8789 2025
rect 8824 1991 8858 2025
rect 8893 1991 8927 2025
rect 8962 1991 8996 2025
rect 9031 1991 9065 2025
rect 9100 1991 9134 2025
rect 9169 1991 9203 2025
rect 9238 1991 9272 2025
rect 9307 1991 9341 2025
rect 9376 1991 9410 2025
rect 9444 1991 9478 2025
rect 9512 1991 9546 2025
rect 9580 1991 9614 2025
rect 9648 1991 9682 2025
rect 9716 1991 9750 2025
<< locali >>
rect -24 2328 69 2362
rect -24 2294 54 2328
rect -24 2260 69 2294
rect -24 2226 78 2260
rect 1641 2228 1905 2260
rect -24 1372 10 1376
rect 44 1372 78 1376
rect -24 1332 78 1372
rect -24 1298 10 1332
rect 44 1298 78 1332
rect -24 1265 78 1298
rect 181 2091 1549 2101
rect 181 2073 371 2091
rect 405 2073 439 2091
rect 181 2039 329 2073
rect 363 2057 371 2073
rect 437 2057 439 2073
rect 473 2073 507 2091
rect 541 2073 575 2091
rect 609 2073 643 2091
rect 677 2073 711 2091
rect 745 2073 779 2091
rect 473 2057 477 2073
rect 541 2057 551 2073
rect 609 2057 625 2073
rect 677 2057 699 2073
rect 745 2057 773 2073
rect 813 2057 847 2091
rect 881 2057 915 2091
rect 949 2073 983 2091
rect 1017 2073 1051 2091
rect 1085 2073 1119 2091
rect 1153 2073 1187 2091
rect 1221 2073 1255 2091
rect 955 2057 983 2073
rect 1029 2057 1051 2073
rect 1103 2057 1119 2073
rect 1177 2057 1187 2073
rect 1252 2057 1255 2073
rect 1289 2073 1323 2091
rect 1357 2073 1391 2091
rect 1425 2073 1549 2091
rect 1289 2057 1293 2073
rect 1357 2057 1368 2073
rect 1425 2057 1443 2073
rect 363 2039 403 2057
rect 437 2039 477 2057
rect 511 2039 551 2057
rect 585 2039 625 2057
rect 659 2039 699 2057
rect 733 2039 773 2057
rect 807 2039 847 2057
rect 881 2039 921 2057
rect 955 2039 995 2057
rect 1029 2039 1069 2057
rect 1103 2039 1143 2057
rect 1177 2039 1218 2057
rect 1252 2039 1293 2057
rect 1327 2039 1368 2057
rect 1402 2039 1443 2057
rect 1477 2039 1549 2073
rect 181 2029 1549 2039
rect 181 1995 209 2029
rect 243 2023 1549 2029
rect 271 2011 1549 2023
rect 181 1989 237 1995
rect 181 1955 271 1989
rect 1459 1959 1549 2011
rect 181 1921 209 1955
rect 414 1923 427 1957
rect 464 1923 501 1957
rect 540 1923 572 1957
rect 619 1923 642 1957
rect 698 1923 712 1957
rect 776 1923 782 1957
rect 816 1923 820 1957
rect 886 1923 898 1957
rect 956 1923 976 1957
rect 1026 1923 1054 1957
rect 1096 1923 1132 1957
rect 1166 1923 1202 1957
rect 1244 1923 1272 1957
rect 1493 1955 1549 1959
rect 181 1887 271 1921
rect 181 1881 237 1887
rect 181 1847 209 1881
rect 1459 1921 1487 1925
rect 1521 1921 1549 1955
rect 1459 1891 1549 1921
rect 1493 1882 1549 1891
rect 243 1847 271 1853
rect 181 1819 271 1847
rect 181 1807 237 1819
rect 181 1773 209 1807
rect 243 1773 271 1785
rect 181 1751 271 1773
rect 181 1733 237 1751
rect 181 1699 209 1733
rect 243 1699 271 1717
rect 181 1683 271 1699
rect 181 1659 237 1683
rect 181 1625 209 1659
rect 243 1625 271 1649
rect 181 1615 271 1625
rect 181 1585 237 1615
rect 181 1551 209 1585
rect 243 1551 271 1581
rect 181 1547 271 1551
rect 181 1513 237 1547
rect 181 1511 271 1513
rect 181 1477 209 1511
rect 243 1479 271 1511
rect 181 1445 237 1477
rect 181 1437 271 1445
rect 181 1403 209 1437
rect 243 1411 271 1437
rect 181 1377 237 1403
rect 181 1363 271 1377
rect 181 1329 209 1363
rect 243 1343 271 1363
rect 181 1309 237 1329
rect 181 1289 271 1309
rect 181 1255 209 1289
rect 243 1275 271 1289
rect 181 1241 237 1255
rect 181 1215 271 1241
rect 181 1181 209 1215
rect 243 1181 271 1215
rect 181 1142 271 1181
rect 181 1108 209 1142
rect 243 1123 271 1142
rect 181 1089 237 1108
rect 181 1069 271 1089
rect 181 1035 209 1069
rect 243 1055 271 1069
rect 181 1021 237 1035
rect 181 996 271 1021
rect 181 962 209 996
rect 243 987 271 996
rect 181 953 237 962
rect 181 923 271 953
rect 181 889 209 923
rect 243 919 271 923
rect 181 885 237 889
rect 181 851 271 885
rect 181 850 237 851
rect 181 816 209 850
rect 243 816 271 817
rect 181 783 271 816
rect 181 777 237 783
rect 181 743 209 777
rect 243 743 271 749
rect 181 715 271 743
rect 181 704 237 715
rect 181 670 209 704
rect 243 670 271 681
rect 181 647 271 670
rect 181 631 237 647
rect 181 597 209 631
rect 243 597 271 613
rect 181 579 271 597
rect 181 558 237 579
rect 181 524 209 558
rect 243 524 271 545
rect 181 511 271 524
rect 181 485 237 511
rect 181 451 209 485
rect 243 451 271 477
rect 362 1813 396 1839
rect 362 1745 396 1767
rect 362 1677 396 1695
rect 362 1609 396 1623
rect 362 1541 396 1551
rect 362 1473 396 1479
rect 362 1405 396 1407
rect 362 1369 396 1371
rect 362 1297 396 1303
rect 362 1225 396 1235
rect 362 1153 396 1167
rect 362 1081 396 1099
rect 362 1009 396 1031
rect 362 937 396 963
rect 362 865 396 895
rect 362 793 396 827
rect 362 725 396 759
rect 362 657 396 687
rect 362 589 396 615
rect 362 521 396 543
rect 525 1813 559 1839
rect 525 1745 559 1767
rect 525 1677 559 1695
rect 525 1609 559 1623
rect 525 1541 559 1551
rect 525 1473 559 1479
rect 525 1405 559 1407
rect 525 1369 559 1371
rect 525 1297 559 1303
rect 525 1225 559 1235
rect 525 1153 559 1167
rect 525 1081 559 1099
rect 525 1009 559 1031
rect 525 937 559 963
rect 525 865 559 895
rect 525 793 559 827
rect 525 725 559 759
rect 525 657 559 687
rect 525 589 559 615
rect 525 521 559 543
rect 688 1813 722 1839
rect 688 1745 722 1767
rect 688 1677 722 1695
rect 688 1609 722 1623
rect 688 1541 722 1551
rect 688 1473 722 1479
rect 688 1405 722 1407
rect 688 1369 722 1371
rect 688 1297 722 1303
rect 688 1225 722 1235
rect 688 1153 722 1167
rect 688 1081 722 1099
rect 688 1009 722 1031
rect 688 937 722 963
rect 688 865 722 895
rect 688 793 722 827
rect 688 725 722 759
rect 688 657 722 687
rect 688 589 722 615
rect 688 521 722 543
rect 851 1813 885 1839
rect 851 1745 885 1767
rect 851 1677 885 1695
rect 851 1609 885 1623
rect 851 1541 885 1551
rect 851 1473 885 1479
rect 851 1405 885 1407
rect 851 1369 885 1371
rect 851 1297 885 1303
rect 851 1225 885 1235
rect 851 1153 885 1167
rect 851 1081 885 1099
rect 851 1009 885 1031
rect 851 937 885 963
rect 851 865 885 895
rect 851 793 885 827
rect 851 725 885 759
rect 851 657 885 687
rect 851 589 885 615
rect 851 521 885 543
rect 1014 1813 1048 1839
rect 1014 1745 1048 1767
rect 1014 1677 1048 1695
rect 1014 1609 1048 1623
rect 1014 1541 1048 1551
rect 1014 1473 1048 1479
rect 1014 1405 1048 1407
rect 1014 1369 1048 1371
rect 1014 1297 1048 1303
rect 1014 1225 1048 1235
rect 1014 1153 1048 1167
rect 1014 1081 1048 1099
rect 1014 1009 1048 1031
rect 1014 937 1048 963
rect 1014 865 1048 895
rect 1014 793 1048 827
rect 1014 725 1048 759
rect 1014 657 1048 687
rect 1014 589 1048 615
rect 1014 521 1048 543
rect 1177 1813 1211 1839
rect 1177 1745 1211 1767
rect 1177 1677 1211 1695
rect 1177 1609 1211 1623
rect 1177 1541 1211 1551
rect 1177 1473 1211 1479
rect 1177 1405 1211 1407
rect 1177 1369 1211 1371
rect 1177 1297 1211 1303
rect 1177 1225 1211 1235
rect 1177 1153 1211 1167
rect 1177 1081 1211 1099
rect 1177 1009 1211 1031
rect 1177 937 1211 963
rect 1177 865 1211 895
rect 1177 793 1211 827
rect 1177 725 1211 759
rect 1177 657 1211 687
rect 1177 589 1211 615
rect 1177 521 1211 543
rect 1340 1813 1374 1839
rect 1340 1745 1374 1767
rect 1340 1677 1374 1695
rect 1340 1609 1374 1623
rect 1340 1541 1374 1551
rect 1340 1473 1374 1479
rect 1340 1405 1374 1407
rect 1340 1369 1374 1371
rect 1340 1297 1374 1303
rect 1340 1225 1374 1235
rect 1340 1153 1374 1167
rect 1340 1081 1374 1099
rect 1340 1009 1374 1031
rect 1340 937 1374 963
rect 1340 865 1374 895
rect 1340 793 1374 827
rect 1340 725 1374 759
rect 1340 657 1374 687
rect 1340 589 1374 615
rect 1340 521 1374 543
rect 1459 1848 1487 1857
rect 1521 1848 1549 1882
rect 1459 1823 1549 1848
rect 1493 1809 1549 1823
rect 1459 1775 1487 1789
rect 1521 1775 1549 1809
rect 1459 1755 1549 1775
rect 1493 1736 1549 1755
rect 1459 1702 1487 1721
rect 1521 1702 1549 1736
rect 1459 1687 1549 1702
rect 1493 1663 1549 1687
rect 1459 1629 1487 1653
rect 1521 1629 1549 1663
rect 1459 1619 1549 1629
rect 1493 1590 1549 1619
rect 1459 1556 1487 1585
rect 1521 1556 1549 1590
rect 1459 1551 1549 1556
rect 1493 1517 1549 1551
rect 1459 1483 1487 1517
rect 1521 1483 1549 1517
rect 1493 1449 1549 1483
rect 1459 1444 1549 1449
rect 1459 1415 1487 1444
rect 1521 1410 1549 1444
rect 1493 1381 1549 1410
rect 1459 1371 1549 1381
rect 1459 1347 1487 1371
rect 1521 1337 1549 1371
rect 1493 1313 1549 1337
rect 1459 1298 1549 1313
rect 1459 1279 1487 1298
rect 1521 1264 1549 1298
rect 1493 1245 1549 1264
rect 1459 1225 1549 1245
rect 1459 1211 1487 1225
rect 1521 1191 1549 1225
rect 1493 1177 1549 1191
rect 1459 1151 1549 1177
rect 1459 1143 1487 1151
rect 1521 1117 1549 1151
rect 1493 1109 1549 1117
rect 1459 1077 1549 1109
rect 1459 1075 1487 1077
rect 1521 1043 1549 1077
rect 1493 1041 1549 1043
rect 1459 1007 1549 1041
rect 1493 1003 1549 1007
rect 1459 969 1487 973
rect 1521 969 1549 1003
rect 1459 939 1549 969
rect 1493 929 1549 939
rect 1459 895 1487 905
rect 1521 895 1549 929
rect 1459 871 1549 895
rect 1493 855 1549 871
rect 1459 821 1487 837
rect 1521 821 1549 855
rect 1459 803 1549 821
rect 1493 781 1549 803
rect 1459 747 1487 769
rect 1521 747 1549 781
rect 1459 735 1549 747
rect 1493 707 1549 735
rect 1459 673 1487 701
rect 1521 673 1549 707
rect 1459 667 1549 673
rect 1493 633 1549 667
rect 1459 599 1487 633
rect 1521 599 1549 633
rect 1493 565 1549 599
rect 1459 559 1549 565
rect 1459 531 1487 559
rect 1521 525 1549 559
rect 1493 497 1549 525
rect 1459 485 1549 497
rect 181 395 271 451
rect 1459 463 1487 485
rect 1521 451 1549 485
rect 1493 429 1549 451
rect 1459 411 1549 429
rect 1459 395 1487 411
rect 181 367 305 395
rect 181 333 253 367
rect 287 361 305 367
rect 339 367 373 395
rect 407 367 441 395
rect 339 361 347 367
rect 407 361 440 367
rect 475 361 509 395
rect 543 367 577 395
rect 611 367 645 395
rect 567 361 577 367
rect 643 361 645 367
rect 679 367 713 395
rect 747 367 781 395
rect 815 367 849 395
rect 883 367 917 395
rect 679 361 685 367
rect 747 361 761 367
rect 815 361 837 367
rect 883 361 913 367
rect 951 361 985 395
rect 1019 367 1053 395
rect 1087 367 1121 395
rect 1155 367 1189 395
rect 1223 367 1257 395
rect 1291 367 1325 395
rect 1023 361 1053 367
rect 1099 361 1121 367
rect 1174 361 1189 367
rect 1249 361 1257 367
rect 1324 361 1325 367
rect 1359 377 1487 395
rect 1521 377 1549 411
rect 1359 367 1549 377
rect 1359 361 1365 367
rect 287 333 347 361
rect 381 333 440 361
rect 474 333 533 361
rect 567 333 609 361
rect 643 333 685 361
rect 719 333 761 361
rect 795 333 837 361
rect 871 333 913 361
rect 947 333 989 361
rect 1023 333 1065 361
rect 1099 333 1140 361
rect 1174 333 1215 361
rect 1249 333 1290 361
rect 1324 333 1365 361
rect 1399 333 1549 367
rect 181 305 1549 333
rect 1641 754 1648 2228
rect 1898 754 1905 2228
rect 3435 2250 3469 2260
rect 3503 2250 3537 2362
rect 3435 2210 3537 2250
rect 3435 2178 3469 2210
rect 3503 2178 3537 2210
rect 1641 730 1905 754
rect 1641 681 1648 730
rect 1682 681 1720 730
rect 1754 681 1792 730
rect 1826 681 1864 730
rect 1898 681 1905 730
rect 1641 662 1905 681
rect 1641 608 1648 662
rect 1682 608 1720 662
rect 1754 608 1792 662
rect 1826 608 1864 662
rect 1898 608 1905 662
rect 1641 594 1905 608
rect 1641 535 1648 594
rect 1682 535 1720 594
rect 1754 535 1792 594
rect 1826 535 1864 594
rect 1898 535 1905 594
rect 1641 526 1905 535
rect 1641 462 1648 526
rect 1682 462 1720 526
rect 1754 462 1792 526
rect 1826 462 1864 526
rect 1898 462 1905 526
rect 1641 458 1905 462
rect 1641 424 1648 458
rect 1682 424 1720 458
rect 1754 424 1792 458
rect 1826 424 1864 458
rect 1898 424 1905 458
rect 1641 423 1905 424
rect 1641 356 1648 423
rect 1682 356 1720 423
rect 1754 356 1792 423
rect 1826 356 1864 423
rect 1898 356 1905 423
rect 1641 350 1905 356
rect -24 188 10 211
rect 44 188 78 211
rect -24 177 78 188
rect 10 148 78 177
rect -24 114 10 143
rect 44 138 78 148
rect 1641 288 1648 350
rect 1682 288 1720 350
rect 1754 288 1792 350
rect 1826 288 1864 350
rect 1898 288 1905 350
rect 2052 2029 2120 2107
rect 3106 2073 3140 2107
rect 3174 2073 3282 2107
rect 3135 2039 3176 2073
rect 3210 2039 3282 2073
rect 2052 2025 2092 2029
rect 2086 1995 2092 2025
rect 3106 2005 3180 2039
rect 2126 1995 2154 2005
rect 2086 1991 2154 1995
rect 2052 1957 2154 1991
rect 2291 1923 2303 1957
rect 2341 1923 2376 1957
rect 2416 1923 2445 1957
rect 2495 1923 2514 1957
rect 2574 1923 2583 1957
rect 2617 1923 2619 1957
rect 2686 1923 2697 1957
rect 2755 1923 2775 1957
rect 2823 1923 2853 1957
rect 2891 1923 2925 1957
rect 2965 1923 2993 1957
rect 2246 1813 2280 1839
rect 2246 1745 2280 1767
rect 2246 1677 2280 1695
rect 2246 1609 2280 1623
rect 2246 1541 2280 1551
rect 2246 1473 2280 1479
rect 2246 1405 2280 1407
rect 2246 1369 2280 1371
rect 2246 1297 2280 1303
rect 2246 1225 2280 1235
rect 2246 1153 2280 1167
rect 2246 1081 2280 1099
rect 2246 1009 2280 1031
rect 2246 937 2280 963
rect 2246 865 2280 895
rect 2246 793 2280 827
rect 2246 725 2280 759
rect 2246 657 2280 687
rect 2246 589 2280 615
rect 2246 521 2280 543
rect 2409 1813 2443 1839
rect 2409 1745 2443 1767
rect 2409 1677 2443 1695
rect 2409 1609 2443 1623
rect 2409 1541 2443 1551
rect 2409 1473 2443 1479
rect 2409 1405 2443 1407
rect 2409 1369 2443 1371
rect 2409 1297 2443 1303
rect 2409 1225 2443 1235
rect 2409 1153 2443 1167
rect 2409 1081 2443 1099
rect 2409 1009 2443 1031
rect 2409 937 2443 963
rect 2409 865 2443 895
rect 2409 793 2443 827
rect 2409 725 2443 759
rect 2409 657 2443 687
rect 2409 589 2443 615
rect 2409 521 2443 543
rect 2572 1813 2606 1839
rect 2572 1745 2606 1767
rect 2572 1677 2606 1695
rect 2572 1609 2606 1623
rect 2572 1541 2606 1551
rect 2572 1473 2606 1479
rect 2572 1405 2606 1407
rect 2572 1369 2606 1371
rect 2572 1297 2606 1303
rect 2572 1225 2606 1235
rect 2572 1153 2606 1167
rect 2572 1081 2606 1099
rect 2572 1009 2606 1031
rect 2572 937 2606 963
rect 2572 865 2606 895
rect 2572 793 2606 827
rect 2572 725 2606 759
rect 2572 657 2606 687
rect 2572 589 2606 615
rect 2572 521 2606 543
rect 2735 1813 2769 1839
rect 2735 1745 2769 1767
rect 2735 1677 2769 1695
rect 2735 1609 2769 1623
rect 2735 1541 2769 1551
rect 2735 1473 2769 1479
rect 2735 1405 2769 1407
rect 2735 1369 2769 1371
rect 2735 1297 2769 1303
rect 2735 1225 2769 1235
rect 2735 1153 2769 1167
rect 2735 1081 2769 1099
rect 2735 1009 2769 1031
rect 2735 937 2769 963
rect 2735 865 2769 895
rect 2735 793 2769 827
rect 2735 725 2769 759
rect 2735 657 2769 687
rect 2735 589 2769 615
rect 2735 521 2769 543
rect 2898 1813 2932 1839
rect 2898 1745 2932 1767
rect 2898 1677 2932 1695
rect 2898 1609 2932 1623
rect 2898 1541 2932 1551
rect 2898 1473 2932 1479
rect 2898 1405 2932 1407
rect 2898 1369 2932 1371
rect 2898 1297 2932 1303
rect 2898 1225 2932 1235
rect 2898 1153 2932 1167
rect 2898 1081 2932 1099
rect 2898 1009 2932 1031
rect 2898 937 2932 963
rect 2898 865 2932 895
rect 2898 793 2932 827
rect 2898 725 2932 759
rect 2898 657 2932 687
rect 2898 589 2932 615
rect 2898 521 2932 543
rect 3061 1813 3095 1839
rect 3061 1745 3095 1767
rect 3061 1677 3095 1695
rect 3061 1609 3095 1623
rect 3061 1541 3095 1551
rect 3061 1473 3095 1479
rect 3061 1405 3095 1407
rect 3061 1369 3095 1371
rect 3061 1297 3095 1303
rect 3061 1225 3095 1235
rect 3061 1153 3095 1167
rect 3061 1081 3095 1099
rect 3061 1009 3095 1031
rect 3061 937 3095 963
rect 3061 865 3095 895
rect 3061 793 3095 827
rect 3061 725 3095 759
rect 3061 657 3095 687
rect 3061 589 3095 615
rect 3061 521 3095 543
rect 3180 969 3220 985
rect 3254 969 3282 985
rect 3180 929 3282 969
rect 3180 910 3220 929
rect 3254 910 3282 929
rect 3180 451 3220 468
rect 3254 451 3282 468
rect 3180 434 3282 451
rect 3180 411 3248 434
rect 3180 395 3220 411
rect 2154 393 2450 395
rect 2492 393 3220 395
rect 2154 367 2228 393
rect 3214 377 3220 393
rect 3254 377 3282 400
rect 2052 333 2136 359
rect 2170 333 2228 367
rect 2052 325 2228 333
rect 2052 291 2160 325
rect 2194 291 2228 325
rect 3214 291 3282 377
rect 1641 277 1905 288
rect 1641 220 1648 277
rect 1682 220 1720 277
rect 1754 220 1792 277
rect 1826 220 1864 277
rect 1898 220 1905 277
rect 1641 204 1905 220
rect 1641 170 1648 204
rect 1682 170 1720 204
rect 1754 170 1792 204
rect 1826 170 1864 204
rect 1898 170 1905 204
rect 1641 138 1905 170
rect -24 36 44 114
rect 3342 104 3435 138
rect 3342 70 3351 104
rect 3385 70 3425 104
rect 3459 70 3537 104
rect 3342 36 3376 70
rect 3410 36 3537 70
rect 3750 2260 3818 2362
rect 10108 2328 10262 2362
rect 10108 2294 10145 2328
rect 10179 2294 10262 2328
rect 3750 2254 3852 2260
rect 3784 2220 3852 2254
rect 3750 2210 3852 2220
rect 3750 2186 3784 2210
rect 3818 2186 3852 2210
rect 10108 2274 10228 2294
rect 10108 2260 10160 2274
rect 3750 418 3784 452
rect 3818 418 3852 452
rect 4005 2039 4099 2073
rect 4133 2039 4139 2073
rect 4173 2039 4179 2073
rect 4241 2039 4252 2073
rect 4309 2039 4325 2073
rect 4377 2039 4398 2073
rect 4445 2039 4471 2073
rect 4513 2039 4544 2073
rect 4581 2039 4615 2073
rect 4651 2039 4683 2073
rect 4724 2039 4751 2073
rect 4797 2039 4819 2073
rect 4870 2039 4887 2073
rect 4943 2039 4955 2073
rect 5016 2039 5023 2073
rect 5089 2039 5091 2073
rect 5125 2039 5128 2073
rect 5193 2039 5201 2073
rect 5261 2039 5274 2073
rect 5329 2039 5347 2073
rect 5397 2039 5420 2073
rect 5465 2039 5493 2073
rect 5533 2039 5566 2073
rect 5601 2039 5635 2073
rect 5673 2039 5703 2073
rect 5746 2039 5771 2073
rect 5819 2039 5839 2073
rect 5892 2039 5907 2073
rect 5965 2039 5975 2073
rect 6038 2039 6043 2073
rect 6145 2039 6150 2073
rect 6213 2039 6223 2073
rect 6281 2039 6295 2073
rect 6349 2039 6367 2073
rect 6417 2039 6439 2073
rect 6485 2039 6511 2073
rect 6553 2039 6583 2073
rect 6621 2039 6689 2073
rect 4005 2005 4039 2039
rect 4005 1937 4039 1965
rect 6655 2001 6689 2039
rect 4226 1923 4250 1957
rect 4298 1923 4323 1957
rect 4370 1923 4396 1957
rect 4442 1923 4469 1957
rect 4514 1923 4542 1957
rect 4586 1923 4615 1957
rect 4658 1923 4688 1957
rect 4730 1923 4768 1957
rect 4802 1923 4840 1957
rect 4874 1923 4912 1957
rect 4946 1923 4985 1957
rect 5019 1923 5058 1957
rect 5092 1923 5131 1957
rect 5165 1923 5204 1957
rect 5238 1923 5254 1957
rect 5447 1923 5459 1957
rect 5497 1923 5535 1957
rect 5570 1923 5609 1957
rect 5645 1923 5682 1957
rect 5721 1923 5755 1957
rect 5797 1923 5827 1957
rect 5872 1923 5899 1957
rect 5947 1923 5971 1957
rect 6022 1923 6043 1957
rect 6077 1923 6115 1957
rect 6149 1923 6187 1957
rect 6221 1923 6259 1957
rect 6293 1923 6331 1957
rect 6365 1923 6403 1957
rect 6437 1923 6475 1957
rect 6509 1923 6525 1957
rect 6655 1931 6689 1965
rect 4005 1869 4039 1891
rect 4005 1801 4039 1817
rect 4005 1733 4039 1743
rect 4005 1665 4039 1669
rect 4005 1629 4039 1631
rect 4005 1555 4039 1563
rect 4005 1481 4039 1495
rect 4005 1407 4039 1427
rect 4005 1333 4039 1359
rect 4005 1259 4039 1291
rect 4005 1189 4039 1223
rect 4005 1121 4039 1151
rect 4005 1053 4039 1077
rect 4005 985 4039 1003
rect 4005 917 4039 929
rect 4005 849 4039 855
rect 4005 814 4039 815
rect 4005 739 4039 747
rect 4005 664 4039 679
rect 4005 589 4039 611
rect 4005 514 4039 555
rect 4131 1813 4165 1839
rect 4131 1745 4165 1767
rect 4131 1677 4165 1695
rect 4131 1609 4165 1623
rect 4131 1541 4165 1551
rect 4131 1473 4165 1479
rect 4131 1405 4165 1407
rect 4131 1369 4165 1371
rect 4131 1297 4165 1303
rect 4131 1225 4165 1235
rect 4131 1153 4165 1167
rect 4131 1081 4165 1099
rect 4131 1009 4165 1031
rect 4131 937 4165 963
rect 4131 865 4165 895
rect 4131 793 4165 827
rect 4131 725 4165 759
rect 4131 657 4165 687
rect 4131 589 4165 615
rect 4131 521 4165 543
rect 4294 1813 4328 1839
rect 4294 1745 4328 1767
rect 4294 1677 4328 1695
rect 4294 1609 4328 1623
rect 4294 1541 4328 1551
rect 4294 1473 4328 1479
rect 4294 1405 4328 1407
rect 4294 1369 4328 1371
rect 4294 1297 4328 1303
rect 4294 1225 4328 1235
rect 4294 1153 4328 1167
rect 4294 1081 4328 1099
rect 4294 1009 4328 1031
rect 4294 937 4328 963
rect 4294 865 4328 895
rect 4294 793 4328 827
rect 4294 725 4328 759
rect 4294 657 4328 687
rect 4294 589 4328 615
rect 4294 521 4328 543
rect 4457 1813 4491 1839
rect 4457 1745 4491 1767
rect 4457 1677 4491 1695
rect 4457 1609 4491 1623
rect 4457 1541 4491 1551
rect 4457 1473 4491 1479
rect 4457 1405 4491 1407
rect 4457 1369 4491 1371
rect 4457 1297 4491 1303
rect 4457 1225 4491 1235
rect 4457 1153 4491 1167
rect 4457 1081 4491 1099
rect 4457 1009 4491 1031
rect 4457 937 4491 963
rect 4457 865 4491 895
rect 4457 793 4491 827
rect 4457 725 4491 759
rect 4457 657 4491 687
rect 4457 589 4491 615
rect 4457 521 4491 543
rect 4620 1813 4654 1839
rect 4620 1745 4654 1767
rect 4620 1677 4654 1695
rect 4620 1609 4654 1623
rect 4620 1541 4654 1551
rect 4620 1473 4654 1479
rect 4620 1405 4654 1407
rect 4620 1369 4654 1371
rect 4620 1297 4654 1303
rect 4620 1225 4654 1235
rect 4620 1153 4654 1167
rect 4620 1081 4654 1099
rect 4620 1009 4654 1031
rect 4620 937 4654 963
rect 4620 865 4654 895
rect 4620 793 4654 827
rect 4620 725 4654 759
rect 4620 657 4654 687
rect 4620 589 4654 615
rect 4620 521 4654 543
rect 4783 1813 4817 1839
rect 4783 1745 4817 1767
rect 4783 1677 4817 1695
rect 4783 1609 4817 1623
rect 4783 1541 4817 1551
rect 4783 1473 4817 1479
rect 4783 1405 4817 1407
rect 4783 1369 4817 1371
rect 4783 1297 4817 1303
rect 4783 1225 4817 1235
rect 4783 1153 4817 1167
rect 4783 1081 4817 1099
rect 4783 1009 4817 1031
rect 4783 937 4817 963
rect 4783 865 4817 895
rect 4783 793 4817 827
rect 4783 725 4817 759
rect 4783 657 4817 687
rect 4783 589 4817 615
rect 4783 521 4817 543
rect 4946 1813 4980 1839
rect 4946 1745 4980 1767
rect 4946 1677 4980 1695
rect 4946 1609 4980 1623
rect 4946 1541 4980 1551
rect 4946 1473 4980 1479
rect 4946 1405 4980 1407
rect 4946 1369 4980 1371
rect 4946 1297 4980 1303
rect 4946 1225 4980 1235
rect 4946 1153 4980 1167
rect 4946 1081 4980 1099
rect 4946 1009 4980 1031
rect 4946 937 4980 963
rect 4946 865 4980 895
rect 4946 793 4980 827
rect 4946 725 4980 759
rect 4946 657 4980 687
rect 4946 589 4980 615
rect 4946 521 4980 543
rect 5109 1813 5143 1839
rect 5109 1745 5143 1767
rect 5109 1677 5143 1695
rect 5109 1609 5143 1623
rect 5109 1541 5143 1551
rect 5109 1473 5143 1479
rect 5109 1405 5143 1407
rect 5109 1369 5143 1371
rect 5109 1297 5143 1303
rect 5109 1225 5143 1235
rect 5109 1153 5143 1167
rect 5109 1081 5143 1099
rect 5109 1009 5143 1031
rect 5109 937 5143 963
rect 5109 865 5143 895
rect 5109 793 5143 827
rect 5109 725 5143 759
rect 5109 657 5143 687
rect 5109 589 5143 615
rect 5109 521 5143 543
rect 5272 1813 5306 1839
rect 5272 1745 5306 1767
rect 5272 1677 5306 1695
rect 5272 1609 5306 1623
rect 5272 1541 5306 1551
rect 5272 1473 5306 1479
rect 5272 1405 5306 1407
rect 5272 1369 5306 1371
rect 5272 1297 5306 1303
rect 5272 1225 5306 1235
rect 5272 1153 5306 1167
rect 5272 1081 5306 1099
rect 5272 1009 5306 1031
rect 5272 937 5306 963
rect 5272 865 5306 895
rect 5272 793 5306 827
rect 5272 725 5306 759
rect 5272 657 5306 687
rect 5272 589 5306 615
rect 5272 521 5306 543
rect 5395 1813 5429 1839
rect 5395 1745 5429 1767
rect 5395 1677 5429 1695
rect 5395 1609 5429 1623
rect 5395 1541 5429 1551
rect 5395 1473 5429 1479
rect 5395 1405 5429 1407
rect 5395 1369 5429 1371
rect 5395 1297 5429 1303
rect 5395 1225 5429 1235
rect 5395 1153 5429 1167
rect 5395 1081 5429 1099
rect 5395 1009 5429 1031
rect 5395 937 5429 963
rect 5395 865 5429 895
rect 5395 793 5429 827
rect 5395 725 5429 759
rect 5395 657 5429 687
rect 5395 589 5429 615
rect 5395 521 5429 543
rect 5558 1813 5592 1839
rect 5558 1745 5592 1767
rect 5558 1677 5592 1695
rect 5558 1609 5592 1623
rect 5558 1541 5592 1551
rect 5558 1473 5592 1479
rect 5558 1405 5592 1407
rect 5558 1369 5592 1371
rect 5558 1297 5592 1303
rect 5558 1225 5592 1235
rect 5558 1153 5592 1167
rect 5558 1081 5592 1099
rect 5558 1009 5592 1031
rect 5558 937 5592 963
rect 5558 865 5592 895
rect 5558 793 5592 827
rect 5558 725 5592 759
rect 5558 657 5592 687
rect 5558 589 5592 615
rect 5558 521 5592 543
rect 5721 1813 5755 1839
rect 5721 1745 5755 1767
rect 5721 1677 5755 1695
rect 5721 1609 5755 1623
rect 5721 1541 5755 1551
rect 5721 1473 5755 1479
rect 5721 1405 5755 1407
rect 5721 1369 5755 1371
rect 5721 1297 5755 1303
rect 5721 1225 5755 1235
rect 5721 1153 5755 1167
rect 5721 1081 5755 1099
rect 5721 1009 5755 1031
rect 5721 937 5755 963
rect 5721 865 5755 895
rect 5721 793 5755 827
rect 5721 725 5755 759
rect 5721 657 5755 687
rect 5721 589 5755 615
rect 5721 521 5755 543
rect 5884 1813 5918 1839
rect 5884 1745 5918 1767
rect 5884 1677 5918 1695
rect 5884 1609 5918 1623
rect 5884 1541 5918 1551
rect 5884 1473 5918 1479
rect 5884 1405 5918 1407
rect 5884 1369 5918 1371
rect 5884 1297 5918 1303
rect 5884 1225 5918 1235
rect 5884 1153 5918 1167
rect 5884 1081 5918 1099
rect 5884 1009 5918 1031
rect 5884 937 5918 963
rect 5884 865 5918 895
rect 5884 793 5918 827
rect 5884 725 5918 759
rect 5884 657 5918 687
rect 5884 589 5918 615
rect 5884 521 5918 543
rect 6047 1813 6081 1839
rect 6047 1745 6081 1767
rect 6047 1677 6081 1695
rect 6047 1609 6081 1623
rect 6047 1541 6081 1551
rect 6047 1473 6081 1479
rect 6047 1405 6081 1407
rect 6047 1369 6081 1371
rect 6047 1297 6081 1303
rect 6047 1225 6081 1235
rect 6047 1153 6081 1167
rect 6047 1081 6081 1099
rect 6047 1009 6081 1031
rect 6047 937 6081 963
rect 6047 865 6081 895
rect 6047 793 6081 827
rect 6047 725 6081 759
rect 6047 657 6081 687
rect 6047 589 6081 615
rect 6047 521 6081 543
rect 6210 1813 6244 1839
rect 6210 1745 6244 1767
rect 6210 1677 6244 1695
rect 6210 1609 6244 1623
rect 6210 1541 6244 1551
rect 6210 1473 6244 1479
rect 6210 1405 6244 1407
rect 6210 1369 6244 1371
rect 6210 1297 6244 1303
rect 6210 1225 6244 1235
rect 6210 1153 6244 1167
rect 6210 1081 6244 1099
rect 6210 1009 6244 1031
rect 6210 937 6244 963
rect 6210 865 6244 895
rect 6210 793 6244 827
rect 6210 725 6244 759
rect 6210 657 6244 687
rect 6210 589 6244 615
rect 6210 521 6244 543
rect 6373 1813 6407 1839
rect 6373 1745 6407 1767
rect 6373 1677 6407 1695
rect 6373 1609 6407 1623
rect 6373 1541 6407 1551
rect 6373 1473 6407 1479
rect 6373 1405 6407 1407
rect 6373 1369 6407 1371
rect 6373 1297 6407 1303
rect 6373 1225 6407 1235
rect 6373 1153 6407 1167
rect 6373 1081 6407 1099
rect 6373 1009 6407 1031
rect 6373 937 6407 963
rect 6373 865 6407 895
rect 6373 793 6407 827
rect 6373 725 6407 759
rect 6373 657 6407 687
rect 6373 589 6407 615
rect 6373 521 6407 543
rect 6536 1813 6570 1839
rect 6536 1745 6570 1767
rect 6536 1677 6570 1695
rect 6536 1609 6570 1623
rect 6536 1541 6570 1551
rect 6536 1473 6570 1479
rect 6536 1405 6570 1407
rect 6536 1369 6570 1371
rect 6536 1297 6570 1303
rect 6536 1225 6570 1235
rect 6536 1153 6570 1167
rect 6536 1081 6570 1099
rect 6536 1009 6570 1031
rect 6536 937 6570 963
rect 6536 865 6570 895
rect 6536 793 6570 827
rect 6536 725 6570 759
rect 6536 657 6570 687
rect 6536 589 6570 615
rect 6536 521 6570 543
rect 6655 1863 6689 1892
rect 6655 1795 6689 1817
rect 6655 1727 6689 1742
rect 6655 1659 6689 1667
rect 6655 1591 6689 1592
rect 6655 1551 6689 1557
rect 6655 1477 6689 1489
rect 6655 1403 6689 1421
rect 6655 1329 6689 1353
rect 6655 1255 6689 1285
rect 6655 1183 6689 1217
rect 6655 1115 6689 1147
rect 6655 1047 6689 1073
rect 6655 979 6689 999
rect 6655 911 6689 925
rect 6655 843 6689 851
rect 6655 775 6689 777
rect 6655 737 6689 741
rect 6655 663 6689 673
rect 6655 589 6689 605
rect 6655 515 6689 537
rect 4005 439 4039 452
rect 4005 367 4039 405
rect 6655 441 6689 469
rect 6655 367 6689 401
rect 4005 333 4073 367
rect 4112 333 4141 367
rect 4185 333 4209 367
rect 4258 333 4277 367
rect 4331 333 4345 367
rect 4404 333 4413 367
rect 4477 333 4481 367
rect 4515 333 4516 367
rect 4583 333 4589 367
rect 4651 333 4662 367
rect 4719 333 4735 367
rect 4787 333 4808 367
rect 4855 333 4881 367
rect 4923 333 4955 367
rect 4991 333 5025 367
rect 5063 333 5093 367
rect 5137 333 5161 367
rect 5211 333 5229 367
rect 5285 333 5297 367
rect 5359 333 5365 367
rect 5467 333 5473 367
rect 5535 333 5547 367
rect 5603 333 5621 367
rect 5671 333 5695 367
rect 5739 333 5769 367
rect 5807 333 5841 367
rect 5877 333 5909 367
rect 5951 333 5977 367
rect 6025 333 6045 367
rect 6099 333 6113 367
rect 6173 333 6181 367
rect 6247 333 6249 367
rect 6283 333 6287 367
rect 6351 333 6361 367
rect 6419 333 6435 367
rect 6487 333 6509 367
rect 6555 333 6583 367
rect 6617 333 6689 367
rect 6842 668 6944 696
rect 6842 661 6876 668
rect 6910 661 6944 668
rect 6876 627 6910 634
rect 6842 595 6944 627
rect 6842 592 6876 595
rect 6910 592 6944 595
rect 6876 558 6910 561
rect 6842 523 6944 558
rect 6876 522 6910 523
rect 6842 488 6876 489
rect 6910 488 6944 489
rect 6842 454 6944 488
rect 6876 449 6910 454
rect 6842 415 6876 420
rect 7091 2107 10003 2113
rect 7091 2073 7170 2107
rect 7209 2073 7243 2107
rect 7277 2073 7311 2107
rect 7350 2073 7379 2107
rect 7423 2073 7447 2107
rect 7497 2073 7515 2107
rect 7571 2073 7583 2107
rect 7645 2073 7651 2107
rect 7753 2073 7759 2107
rect 7821 2073 7833 2107
rect 7889 2073 7907 2107
rect 7957 2073 7981 2107
rect 8025 2073 8055 2107
rect 8093 2073 8127 2107
rect 8163 2073 8195 2107
rect 8237 2073 8263 2107
rect 8311 2073 8331 2107
rect 8385 2073 8399 2107
rect 8459 2073 8467 2107
rect 8533 2073 8535 2107
rect 8569 2073 8573 2107
rect 8637 2073 8647 2107
rect 8705 2073 8721 2107
rect 8773 2073 8795 2107
rect 8841 2073 8869 2107
rect 8909 2073 8943 2107
rect 8977 2073 9011 2107
rect 9051 2073 9079 2107
rect 9125 2073 9147 2107
rect 9199 2073 9215 2107
rect 9273 2073 9283 2107
rect 9347 2073 9351 2107
rect 9385 2073 9387 2107
rect 9453 2073 9461 2107
rect 9521 2073 9535 2107
rect 9589 2073 9623 2107
rect 9679 2073 9691 2107
rect 9725 2073 9727 2107
rect 9793 2073 9809 2107
rect 9861 2073 9891 2107
rect 9929 2073 10003 2107
rect 7091 2067 10003 2073
rect 7091 2039 7137 2067
rect 7091 2001 7097 2039
rect 7131 2001 7137 2039
rect 9957 2033 10003 2067
rect 7091 1971 7137 2001
rect 7261 1991 7273 2025
rect 7311 1991 7346 2025
rect 7384 1991 7419 2025
rect 7457 1991 7492 2025
rect 7530 1991 7565 2025
rect 7603 1991 7638 2025
rect 7675 1991 7711 2025
rect 7747 1991 7784 2025
rect 7819 1991 7857 2025
rect 7891 1991 7929 2025
rect 7964 1991 8001 2025
rect 8037 1991 8073 2025
rect 8109 1991 8145 2025
rect 8181 1991 8217 2025
rect 8251 1991 8289 2025
rect 8323 1991 8339 2025
rect 8532 1991 8544 2025
rect 8582 1991 8617 2025
rect 8653 1991 8686 2025
rect 8728 1991 8755 2025
rect 8803 1991 8824 2025
rect 8878 1991 8893 2025
rect 8952 1991 8962 2025
rect 9026 1991 9031 2025
rect 9065 1991 9066 2025
rect 9134 1991 9140 2025
rect 9203 1991 9214 2025
rect 9272 1991 9288 2025
rect 9341 1991 9362 2025
rect 9410 1991 9436 2025
rect 9478 1991 9510 2025
rect 9546 1991 9580 2025
rect 9618 1991 9648 2025
rect 9692 1991 9716 2025
rect 9957 1999 9963 2033
rect 9997 1999 10003 2033
rect 7091 1926 7097 1971
rect 7131 1926 7137 1971
rect 9957 1965 10003 1999
rect 7091 1903 7137 1926
rect 7091 1851 7097 1903
rect 7131 1851 7137 1903
rect 7091 1835 7137 1851
rect 7091 1776 7097 1835
rect 7131 1776 7137 1835
rect 7091 1767 7137 1776
rect 7091 1701 7097 1767
rect 7131 1701 7137 1767
rect 7091 1699 7137 1701
rect 7091 1665 7097 1699
rect 7131 1665 7137 1699
rect 7091 1660 7137 1665
rect 7091 1597 7097 1660
rect 7131 1597 7137 1660
rect 7091 1585 7137 1597
rect 7091 1529 7097 1585
rect 7131 1529 7137 1585
rect 7091 1510 7137 1529
rect 7091 1461 7097 1510
rect 7131 1461 7137 1510
rect 7091 1435 7137 1461
rect 7091 1393 7097 1435
rect 7131 1393 7137 1435
rect 7091 1360 7137 1393
rect 7091 1325 7097 1360
rect 7131 1325 7137 1360
rect 7091 1291 7137 1325
rect 7091 1251 7097 1291
rect 7131 1251 7137 1291
rect 7091 1223 7137 1251
rect 7091 1176 7097 1223
rect 7131 1176 7137 1223
rect 7091 1155 7137 1176
rect 7091 1101 7097 1155
rect 7131 1101 7137 1155
rect 7091 1087 7137 1101
rect 7091 1027 7097 1087
rect 7131 1027 7137 1087
rect 7091 1019 7137 1027
rect 7091 953 7097 1019
rect 7131 953 7137 1019
rect 7091 951 7137 953
rect 7091 917 7097 951
rect 7131 917 7137 951
rect 7091 913 7137 917
rect 7091 849 7097 913
rect 7131 849 7137 913
rect 7091 839 7137 849
rect 7091 781 7097 839
rect 7131 781 7137 839
rect 7091 765 7137 781
rect 7091 713 7097 765
rect 7131 713 7137 765
rect 7091 691 7137 713
rect 7091 645 7097 691
rect 7131 645 7137 691
rect 7091 617 7137 645
rect 7091 583 7097 617
rect 7131 583 7137 617
rect 7091 554 7137 583
rect 7091 509 7097 554
rect 7131 509 7137 554
rect 7216 1881 7250 1907
rect 7216 1813 7250 1835
rect 7216 1745 7250 1763
rect 7216 1677 7250 1691
rect 7216 1609 7250 1619
rect 7216 1541 7250 1547
rect 7216 1473 7250 1475
rect 7216 1437 7250 1439
rect 7216 1365 7250 1371
rect 7216 1293 7250 1303
rect 7216 1221 7250 1235
rect 7216 1149 7250 1167
rect 7216 1077 7250 1099
rect 7216 1005 7250 1031
rect 7216 933 7250 963
rect 7216 861 7250 895
rect 7216 793 7250 827
rect 7216 725 7250 755
rect 7216 657 7250 683
rect 7216 589 7250 611
rect 7379 1881 7413 1907
rect 7379 1813 7413 1835
rect 7379 1745 7413 1763
rect 7379 1677 7413 1691
rect 7379 1609 7413 1619
rect 7379 1541 7413 1547
rect 7379 1473 7413 1475
rect 7379 1437 7413 1439
rect 7379 1365 7413 1371
rect 7379 1293 7413 1303
rect 7379 1221 7413 1235
rect 7379 1149 7413 1167
rect 7379 1077 7413 1099
rect 7379 1005 7413 1031
rect 7379 933 7413 963
rect 7379 861 7413 895
rect 7379 793 7413 827
rect 7379 725 7413 755
rect 7379 657 7413 683
rect 7379 589 7413 611
rect 7542 1881 7576 1907
rect 7542 1813 7576 1835
rect 7542 1745 7576 1763
rect 7542 1677 7576 1691
rect 7542 1609 7576 1619
rect 7542 1541 7576 1547
rect 7542 1473 7576 1475
rect 7542 1437 7576 1439
rect 7542 1365 7576 1371
rect 7542 1293 7576 1303
rect 7542 1221 7576 1235
rect 7542 1149 7576 1167
rect 7542 1077 7576 1099
rect 7542 1005 7576 1031
rect 7542 933 7576 963
rect 7542 861 7576 895
rect 7542 793 7576 827
rect 7542 725 7576 755
rect 7542 657 7576 683
rect 7542 589 7576 611
rect 7705 1881 7739 1907
rect 7705 1813 7739 1835
rect 7705 1745 7739 1763
rect 7705 1677 7739 1691
rect 7705 1609 7739 1619
rect 7705 1541 7739 1547
rect 7705 1473 7739 1475
rect 7705 1437 7739 1439
rect 7705 1365 7739 1371
rect 7705 1293 7739 1303
rect 7705 1221 7739 1235
rect 7705 1149 7739 1167
rect 7705 1077 7739 1099
rect 7705 1005 7739 1031
rect 7705 933 7739 963
rect 7705 861 7739 895
rect 7705 793 7739 827
rect 7705 725 7739 755
rect 7705 657 7739 683
rect 7705 589 7739 611
rect 7868 1881 7902 1907
rect 7868 1813 7902 1835
rect 7868 1745 7902 1763
rect 7868 1677 7902 1691
rect 7868 1609 7902 1619
rect 7868 1541 7902 1547
rect 7868 1473 7902 1475
rect 7868 1437 7902 1439
rect 7868 1365 7902 1371
rect 7868 1293 7902 1303
rect 7868 1221 7902 1235
rect 7868 1149 7902 1167
rect 7868 1077 7902 1099
rect 7868 1005 7902 1031
rect 7868 933 7902 963
rect 7868 861 7902 895
rect 7868 793 7902 827
rect 7868 725 7902 755
rect 7868 657 7902 683
rect 7868 589 7902 611
rect 8031 1881 8065 1907
rect 8031 1813 8065 1835
rect 8031 1745 8065 1763
rect 8031 1677 8065 1691
rect 8031 1609 8065 1619
rect 8031 1541 8065 1547
rect 8031 1473 8065 1475
rect 8031 1437 8065 1439
rect 8031 1365 8065 1371
rect 8031 1293 8065 1303
rect 8031 1221 8065 1235
rect 8031 1149 8065 1167
rect 8031 1077 8065 1099
rect 8031 1005 8065 1031
rect 8031 933 8065 963
rect 8031 861 8065 895
rect 8031 793 8065 827
rect 8031 725 8065 755
rect 8031 657 8065 683
rect 8031 589 8065 611
rect 8194 1881 8228 1907
rect 8194 1813 8228 1835
rect 8194 1745 8228 1763
rect 8194 1677 8228 1691
rect 8194 1609 8228 1619
rect 8194 1541 8228 1547
rect 8194 1473 8228 1475
rect 8194 1437 8228 1439
rect 8194 1365 8228 1371
rect 8194 1293 8228 1303
rect 8194 1221 8228 1235
rect 8194 1149 8228 1167
rect 8194 1077 8228 1099
rect 8194 1005 8228 1031
rect 8194 933 8228 963
rect 8194 861 8228 895
rect 8194 793 8228 827
rect 8194 725 8228 755
rect 8194 657 8228 683
rect 8194 589 8228 611
rect 8357 1881 8391 1907
rect 9957 1925 9963 1965
rect 9997 1925 10003 1965
rect 8357 1813 8391 1835
rect 8357 1745 8391 1763
rect 8357 1677 8391 1691
rect 8357 1609 8391 1619
rect 8357 1541 8391 1547
rect 8357 1473 8391 1475
rect 8357 1437 8391 1439
rect 8357 1365 8391 1371
rect 8357 1293 8391 1303
rect 8357 1221 8391 1235
rect 8357 1149 8391 1167
rect 8357 1077 8391 1099
rect 8357 1005 8391 1031
rect 8357 933 8391 963
rect 8357 861 8391 895
rect 8357 793 8391 827
rect 8357 725 8391 755
rect 8357 657 8391 683
rect 8357 589 8391 611
rect 9957 1897 10003 1925
rect 8480 1824 8514 1847
rect 8480 1749 8514 1779
rect 8480 1677 8514 1711
rect 8480 1609 8514 1640
rect 8480 1541 8514 1565
rect 8480 1473 8514 1490
rect 8480 1405 8514 1415
rect 8480 1337 8514 1340
rect 8480 1299 8514 1303
rect 8480 1224 8514 1235
rect 8480 1149 8514 1167
rect 8480 1073 8514 1099
rect 8480 997 8514 1031
rect 8480 929 8514 963
rect 8480 861 8514 887
rect 8480 793 8514 811
rect 8480 725 8514 735
rect 8480 657 8514 659
rect 8480 617 8514 623
rect 8480 541 8514 555
rect 7091 475 7137 509
rect 8643 1824 8677 1847
rect 8643 1751 8677 1779
rect 8643 1678 8677 1711
rect 8643 1609 8677 1643
rect 8643 1541 8677 1571
rect 8643 1473 8677 1497
rect 8643 1405 8677 1423
rect 8643 1337 8677 1349
rect 8643 1269 8677 1303
rect 8643 1201 8677 1235
rect 8643 1133 8677 1167
rect 8643 1065 8677 1099
rect 8643 997 8677 1031
rect 8643 929 8677 963
rect 8643 861 8677 895
rect 8643 793 8677 827
rect 8643 725 8677 759
rect 8643 657 8677 691
rect 8643 589 8677 623
rect 8643 539 8677 555
rect 8806 1881 8840 1897
rect 8806 1813 8840 1847
rect 8806 1745 8840 1779
rect 8806 1677 8840 1711
rect 8806 1609 8840 1643
rect 8806 1541 8840 1575
rect 8806 1473 8840 1507
rect 8806 1405 8840 1439
rect 8806 1337 8840 1371
rect 8806 1269 8840 1303
rect 8806 1201 8840 1235
rect 8806 1133 8840 1167
rect 8806 1087 8840 1099
rect 8806 1009 8840 1031
rect 8806 931 8840 963
rect 8806 861 8840 895
rect 8806 793 8840 819
rect 8806 725 8840 741
rect 8806 657 8840 663
rect 8806 619 8840 623
rect 8806 541 8840 555
rect 8480 475 8514 507
rect 8969 1824 9003 1847
rect 8969 1751 9003 1779
rect 8969 1678 9003 1711
rect 8969 1609 9003 1643
rect 8969 1541 9003 1571
rect 8969 1473 9003 1497
rect 8969 1405 9003 1423
rect 8969 1337 9003 1349
rect 8969 1269 9003 1303
rect 8969 1201 9003 1235
rect 8969 1133 9003 1167
rect 8969 1065 9003 1099
rect 8969 997 9003 1031
rect 8969 929 9003 963
rect 8969 861 9003 895
rect 8969 793 9003 827
rect 8969 725 9003 759
rect 8969 657 9003 691
rect 8969 589 9003 623
rect 8969 539 9003 555
rect 9132 1881 9166 1897
rect 9132 1813 9166 1847
rect 9132 1745 9166 1779
rect 9132 1677 9166 1711
rect 9132 1609 9166 1643
rect 9132 1541 9166 1575
rect 9132 1473 9166 1507
rect 9132 1405 9166 1439
rect 9132 1337 9166 1371
rect 9132 1269 9166 1303
rect 9132 1201 9166 1235
rect 9132 1133 9166 1167
rect 9132 1087 9166 1099
rect 9132 1009 9166 1031
rect 9132 931 9166 963
rect 9132 861 9166 895
rect 9132 793 9166 819
rect 9132 725 9166 741
rect 9132 657 9166 663
rect 9132 619 9166 623
rect 9132 541 9166 555
rect 8806 475 8840 507
rect 9295 1824 9329 1847
rect 9295 1751 9329 1779
rect 9295 1678 9329 1711
rect 9295 1609 9329 1643
rect 9295 1541 9329 1571
rect 9295 1473 9329 1497
rect 9295 1405 9329 1423
rect 9295 1337 9329 1349
rect 9295 1269 9329 1303
rect 9295 1201 9329 1235
rect 9295 1133 9329 1167
rect 9295 1065 9329 1099
rect 9295 997 9329 1031
rect 9295 929 9329 963
rect 9295 861 9329 895
rect 9295 793 9329 827
rect 9295 725 9329 759
rect 9295 657 9329 691
rect 9295 589 9329 623
rect 9295 539 9329 555
rect 9458 1881 9492 1897
rect 9458 1813 9492 1847
rect 9458 1745 9492 1779
rect 9458 1677 9492 1711
rect 9458 1609 9492 1643
rect 9458 1541 9492 1575
rect 9458 1473 9492 1507
rect 9458 1405 9492 1439
rect 9458 1337 9492 1371
rect 9458 1269 9492 1303
rect 9458 1201 9492 1235
rect 9458 1133 9492 1167
rect 9458 1087 9492 1099
rect 9458 1009 9492 1031
rect 9458 931 9492 963
rect 9458 861 9492 895
rect 9458 793 9492 819
rect 9458 725 9492 741
rect 9458 657 9492 663
rect 9458 619 9492 623
rect 9458 541 9492 555
rect 9132 475 9166 507
rect 9621 1824 9655 1847
rect 9621 1751 9655 1779
rect 9621 1678 9655 1711
rect 9621 1609 9655 1643
rect 9621 1541 9655 1571
rect 9621 1473 9655 1497
rect 9621 1405 9655 1423
rect 9621 1337 9655 1349
rect 9621 1269 9655 1303
rect 9621 1201 9655 1235
rect 9621 1133 9655 1167
rect 9621 1065 9655 1099
rect 9621 997 9655 1031
rect 9621 929 9655 963
rect 9621 861 9655 895
rect 9621 793 9655 827
rect 9621 725 9655 759
rect 9621 657 9655 691
rect 9621 589 9655 623
rect 9621 539 9655 555
rect 9784 1881 9818 1897
rect 9784 1813 9818 1847
rect 9784 1745 9818 1779
rect 9784 1677 9818 1711
rect 9784 1609 9818 1643
rect 9784 1541 9818 1575
rect 9784 1473 9818 1507
rect 9784 1405 9818 1439
rect 9784 1337 9818 1371
rect 9784 1269 9818 1303
rect 9784 1201 9818 1235
rect 9784 1133 9818 1167
rect 9784 1087 9818 1099
rect 9784 1009 9818 1031
rect 9784 931 9818 963
rect 9784 861 9818 895
rect 9784 793 9818 819
rect 9784 725 9818 741
rect 9784 657 9818 663
rect 9784 619 9818 623
rect 9784 541 9818 555
rect 9458 475 9492 507
rect 9784 475 9818 507
rect 9957 1851 9963 1897
rect 9997 1851 10003 1897
rect 9957 1829 10003 1851
rect 9957 1777 9963 1829
rect 9997 1777 10003 1829
rect 9957 1761 10003 1777
rect 9957 1703 9963 1761
rect 9997 1703 10003 1761
rect 9957 1693 10003 1703
rect 9957 1629 9963 1693
rect 9997 1629 10003 1693
rect 9957 1625 10003 1629
rect 9957 1591 9963 1625
rect 9997 1591 10003 1625
rect 9957 1589 10003 1591
rect 9957 1523 9963 1589
rect 9997 1523 10003 1589
rect 9957 1515 10003 1523
rect 9957 1455 9963 1515
rect 9997 1455 10003 1515
rect 9957 1441 10003 1455
rect 9957 1387 9963 1441
rect 9997 1387 10003 1441
rect 9957 1366 10003 1387
rect 9957 1319 9963 1366
rect 9997 1319 10003 1366
rect 9957 1291 10003 1319
rect 9957 1251 9963 1291
rect 9997 1251 10003 1291
rect 9957 1217 10003 1251
rect 9957 1182 9963 1217
rect 9997 1182 10003 1217
rect 9957 1149 10003 1182
rect 9957 1107 9963 1149
rect 9997 1107 10003 1149
rect 9957 1081 10003 1107
rect 9957 1032 9963 1081
rect 9997 1032 10003 1081
rect 9957 1013 10003 1032
rect 9957 957 9963 1013
rect 9997 957 10003 1013
rect 9957 945 10003 957
rect 9957 882 9963 945
rect 9997 882 10003 945
rect 9957 877 10003 882
rect 9957 843 9963 877
rect 9997 843 10003 877
rect 9957 841 10003 843
rect 9957 775 9963 841
rect 9997 775 10003 841
rect 9957 766 10003 775
rect 9957 707 9963 766
rect 9997 707 10003 766
rect 9957 691 10003 707
rect 9957 639 9963 691
rect 9997 639 10003 691
rect 9957 616 10003 639
rect 9957 571 9963 616
rect 9997 571 10003 616
rect 9957 541 10003 571
rect 9957 503 9963 541
rect 9997 503 10003 541
rect 9957 475 10003 503
rect 7091 469 10003 475
rect 7091 435 7165 469
rect 7203 435 7233 469
rect 7277 435 7301 469
rect 7351 435 7369 469
rect 7425 435 7437 469
rect 7499 435 7505 469
rect 7607 435 7613 469
rect 7675 435 7687 469
rect 7743 435 7761 469
rect 7811 435 7835 469
rect 7879 435 7909 469
rect 7947 435 7981 469
rect 8017 435 8049 469
rect 8091 435 8117 469
rect 8165 435 8185 469
rect 8239 435 8253 469
rect 8313 435 8321 469
rect 8387 435 8389 469
rect 8423 435 8427 469
rect 8491 435 8501 469
rect 8559 435 8575 469
rect 8627 435 8649 469
rect 8695 435 8722 469
rect 8763 435 8795 469
rect 8831 435 8865 469
rect 8902 435 8933 469
rect 8975 435 9001 469
rect 9048 435 9069 469
rect 9121 435 9137 469
rect 9194 435 9205 469
rect 9267 435 9273 469
rect 9340 435 9341 469
rect 9375 435 9379 469
rect 9443 435 9452 469
rect 9511 435 9525 469
rect 9579 435 9598 469
rect 9647 435 9671 469
rect 9715 435 9744 469
rect 9783 435 9817 469
rect 9851 435 9885 469
rect 9924 435 10003 469
rect 7091 429 10003 435
rect 10160 443 10189 472
rect 10223 458 10262 472
rect 10223 443 10228 458
rect 10160 438 10228 443
rect 6910 415 6944 420
rect 6842 385 6944 415
rect 6876 376 6910 385
rect 6842 342 6876 351
rect 6910 342 6944 351
rect 6842 316 6944 342
rect 6876 303 6910 316
rect 6842 269 6876 282
rect 6910 269 6944 282
rect 6842 248 6944 269
rect 10160 331 10262 336
rect 10160 297 10189 331
rect 10223 322 10262 331
rect 10223 297 10228 322
rect 10160 288 10228 297
rect 10160 258 10262 288
rect 10160 248 10189 258
rect 10223 254 10262 258
rect 6876 230 6964 248
rect 6842 196 6876 214
rect 6910 214 6964 230
rect 6998 214 7032 248
rect 10223 224 10228 254
rect 10194 220 10228 224
rect 6910 196 6956 214
rect 6842 180 6956 196
rect 6990 180 7029 214
rect 6842 146 6910 180
rect 6944 146 7032 180
rect 10194 146 10262 220
rect 3852 112 3918 146
rect 3750 78 3902 112
rect 3750 44 3850 78
rect 3884 44 3918 78
rect 6876 44 6944 146
<< viali >>
rect 54 2294 69 2328
rect 69 2294 88 2328
rect 148 2294 182 2328
rect 241 2294 275 2328
rect 334 2294 368 2328
rect 410 2294 444 2328
rect 484 2294 518 2328
rect 558 2294 592 2328
rect 632 2294 666 2328
rect 706 2294 740 2328
rect 780 2294 814 2328
rect 854 2294 888 2328
rect 928 2294 962 2328
rect 1002 2294 1036 2328
rect 1076 2294 1110 2328
rect 1150 2294 1184 2328
rect 1224 2294 1258 2328
rect 1298 2294 1332 2328
rect 1372 2294 1406 2328
rect 1446 2294 1480 2328
rect 1520 2294 1554 2328
rect 1594 2294 1628 2328
rect 1668 2294 1702 2328
rect 1742 2294 1776 2328
rect 1816 2294 1850 2328
rect 1890 2294 1924 2328
rect 1964 2294 1998 2328
rect 2037 2294 2071 2328
rect 2110 2294 2144 2328
rect 2183 2294 2217 2328
rect 2256 2294 2290 2328
rect 2329 2294 2363 2328
rect 2402 2294 2436 2328
rect 2475 2294 2509 2328
rect 2548 2294 2582 2328
rect 2621 2294 2655 2328
rect 2694 2294 2728 2328
rect 2767 2294 2801 2328
rect 2840 2294 2874 2328
rect 2913 2294 2947 2328
rect 2986 2294 3020 2328
rect 3059 2294 3093 2328
rect 3132 2294 3166 2328
rect 3205 2294 3239 2328
rect 3278 2294 3312 2328
rect 3351 2294 3385 2328
rect 3469 2260 3503 2284
rect 10 2176 44 2210
rect 10 2103 44 2137
rect 10 2030 44 2064
rect 10 1957 44 1991
rect 10 1884 44 1918
rect 10 1811 44 1845
rect 10 1738 44 1772
rect 10 1665 44 1699
rect 10 1592 44 1626
rect 10 1519 44 1553
rect 10 1446 44 1480
rect 10 1376 44 1406
rect 10 1372 44 1376
rect 10 1298 44 1332
rect 10 1224 44 1258
rect 10 1150 44 1184
rect 10 1076 44 1110
rect 10 1002 44 1036
rect 10 928 44 962
rect 10 854 44 888
rect 10 780 44 814
rect 10 706 44 740
rect 10 632 44 666
rect 10 558 44 592
rect 10 484 44 518
rect 10 410 44 444
rect 10 336 44 370
rect 329 2039 363 2073
rect 403 2057 405 2073
rect 405 2057 437 2073
rect 477 2057 507 2073
rect 507 2057 511 2073
rect 551 2057 575 2073
rect 575 2057 585 2073
rect 625 2057 643 2073
rect 643 2057 659 2073
rect 699 2057 711 2073
rect 711 2057 733 2073
rect 773 2057 779 2073
rect 779 2057 807 2073
rect 847 2057 881 2073
rect 921 2057 949 2073
rect 949 2057 955 2073
rect 995 2057 1017 2073
rect 1017 2057 1029 2073
rect 1069 2057 1085 2073
rect 1085 2057 1103 2073
rect 1143 2057 1153 2073
rect 1153 2057 1177 2073
rect 1218 2057 1221 2073
rect 1221 2057 1252 2073
rect 1293 2057 1323 2073
rect 1323 2057 1327 2073
rect 1368 2057 1391 2073
rect 1391 2057 1402 2073
rect 403 2039 437 2057
rect 477 2039 511 2057
rect 551 2039 585 2057
rect 625 2039 659 2057
rect 699 2039 733 2057
rect 773 2039 807 2057
rect 847 2039 881 2057
rect 921 2039 955 2057
rect 995 2039 1029 2057
rect 1069 2039 1103 2057
rect 1143 2039 1177 2057
rect 1218 2039 1252 2057
rect 1293 2039 1327 2057
rect 1368 2039 1402 2057
rect 1443 2039 1477 2073
rect 209 2023 243 2029
rect 209 1995 237 2023
rect 237 1995 243 2023
rect 209 1921 237 1955
rect 237 1921 243 1955
rect 427 1923 430 1957
rect 430 1923 461 1957
rect 506 1923 535 1957
rect 535 1923 540 1957
rect 585 1923 606 1957
rect 606 1923 619 1957
rect 664 1923 676 1957
rect 676 1923 698 1957
rect 742 1923 746 1957
rect 746 1923 776 1957
rect 820 1923 852 1957
rect 852 1923 854 1957
rect 898 1923 922 1957
rect 922 1923 932 1957
rect 976 1923 992 1957
rect 992 1923 1010 1957
rect 1054 1923 1062 1957
rect 1062 1923 1088 1957
rect 1132 1923 1166 1957
rect 1210 1923 1236 1957
rect 1236 1923 1244 1957
rect 1288 1923 1306 1957
rect 1306 1923 1322 1957
rect 1487 1925 1493 1955
rect 1493 1925 1521 1955
rect 209 1853 237 1881
rect 237 1853 243 1881
rect 1487 1921 1521 1925
rect 209 1847 243 1853
rect 209 1785 237 1807
rect 237 1785 243 1807
rect 209 1773 243 1785
rect 209 1717 237 1733
rect 237 1717 243 1733
rect 209 1699 243 1717
rect 209 1649 237 1659
rect 237 1649 243 1659
rect 209 1625 243 1649
rect 209 1581 237 1585
rect 237 1581 243 1585
rect 209 1551 243 1581
rect 209 1479 243 1511
rect 209 1477 237 1479
rect 237 1477 243 1479
rect 209 1411 243 1437
rect 209 1403 237 1411
rect 237 1403 243 1411
rect 209 1343 243 1363
rect 209 1329 237 1343
rect 237 1329 243 1343
rect 209 1275 243 1289
rect 209 1255 237 1275
rect 237 1255 243 1275
rect 209 1181 243 1215
rect 209 1123 243 1142
rect 209 1108 237 1123
rect 237 1108 243 1123
rect 209 1055 243 1069
rect 209 1035 237 1055
rect 237 1035 243 1055
rect 209 987 243 996
rect 209 962 237 987
rect 237 962 243 987
rect 209 919 243 923
rect 209 889 237 919
rect 237 889 243 919
rect 209 817 237 850
rect 237 817 243 850
rect 209 816 243 817
rect 209 749 237 777
rect 237 749 243 777
rect 209 743 243 749
rect 209 681 237 704
rect 237 681 243 704
rect 209 670 243 681
rect 209 613 237 631
rect 237 613 243 631
rect 209 597 243 613
rect 209 545 237 558
rect 237 545 243 558
rect 209 524 243 545
rect 209 477 237 485
rect 237 477 243 485
rect 209 451 243 477
rect 362 1839 396 1873
rect 362 1779 396 1801
rect 362 1767 396 1779
rect 362 1711 396 1729
rect 362 1695 396 1711
rect 362 1643 396 1657
rect 362 1623 396 1643
rect 362 1575 396 1585
rect 362 1551 396 1575
rect 362 1507 396 1513
rect 362 1479 396 1507
rect 362 1439 396 1441
rect 362 1407 396 1439
rect 362 1337 396 1369
rect 362 1335 396 1337
rect 362 1269 396 1297
rect 362 1263 396 1269
rect 362 1201 396 1225
rect 362 1191 396 1201
rect 362 1133 396 1153
rect 362 1119 396 1133
rect 362 1065 396 1081
rect 362 1047 396 1065
rect 362 997 396 1009
rect 362 975 396 997
rect 362 929 396 937
rect 362 903 396 929
rect 362 861 396 865
rect 362 831 396 861
rect 362 759 396 793
rect 362 691 396 721
rect 362 687 396 691
rect 362 623 396 649
rect 362 615 396 623
rect 362 555 396 577
rect 362 543 396 555
rect 362 487 396 505
rect 362 471 396 487
rect 525 1839 559 1873
rect 525 1779 559 1801
rect 525 1767 559 1779
rect 525 1711 559 1729
rect 525 1695 559 1711
rect 525 1643 559 1657
rect 525 1623 559 1643
rect 525 1575 559 1585
rect 525 1551 559 1575
rect 525 1507 559 1513
rect 525 1479 559 1507
rect 525 1439 559 1441
rect 525 1407 559 1439
rect 525 1337 559 1369
rect 525 1335 559 1337
rect 525 1269 559 1297
rect 525 1263 559 1269
rect 525 1201 559 1225
rect 525 1191 559 1201
rect 525 1133 559 1153
rect 525 1119 559 1133
rect 525 1065 559 1081
rect 525 1047 559 1065
rect 525 997 559 1009
rect 525 975 559 997
rect 525 929 559 937
rect 525 903 559 929
rect 525 861 559 865
rect 525 831 559 861
rect 525 759 559 793
rect 525 691 559 721
rect 525 687 559 691
rect 525 623 559 649
rect 525 615 559 623
rect 525 555 559 577
rect 525 543 559 555
rect 525 487 559 505
rect 525 471 559 487
rect 688 1839 722 1873
rect 688 1779 722 1801
rect 688 1767 722 1779
rect 688 1711 722 1729
rect 688 1695 722 1711
rect 688 1643 722 1657
rect 688 1623 722 1643
rect 688 1575 722 1585
rect 688 1551 722 1575
rect 688 1507 722 1513
rect 688 1479 722 1507
rect 688 1439 722 1441
rect 688 1407 722 1439
rect 688 1337 722 1369
rect 688 1335 722 1337
rect 688 1269 722 1297
rect 688 1263 722 1269
rect 688 1201 722 1225
rect 688 1191 722 1201
rect 688 1133 722 1153
rect 688 1119 722 1133
rect 688 1065 722 1081
rect 688 1047 722 1065
rect 688 997 722 1009
rect 688 975 722 997
rect 688 929 722 937
rect 688 903 722 929
rect 688 861 722 865
rect 688 831 722 861
rect 688 759 722 793
rect 688 691 722 721
rect 688 687 722 691
rect 688 623 722 649
rect 688 615 722 623
rect 688 555 722 577
rect 688 543 722 555
rect 688 487 722 505
rect 688 471 722 487
rect 851 1839 885 1873
rect 851 1779 885 1801
rect 851 1767 885 1779
rect 851 1711 885 1729
rect 851 1695 885 1711
rect 851 1643 885 1657
rect 851 1623 885 1643
rect 851 1575 885 1585
rect 851 1551 885 1575
rect 851 1507 885 1513
rect 851 1479 885 1507
rect 851 1439 885 1441
rect 851 1407 885 1439
rect 851 1337 885 1369
rect 851 1335 885 1337
rect 851 1269 885 1297
rect 851 1263 885 1269
rect 851 1201 885 1225
rect 851 1191 885 1201
rect 851 1133 885 1153
rect 851 1119 885 1133
rect 851 1065 885 1081
rect 851 1047 885 1065
rect 851 997 885 1009
rect 851 975 885 997
rect 851 929 885 937
rect 851 903 885 929
rect 851 861 885 865
rect 851 831 885 861
rect 851 759 885 793
rect 851 691 885 721
rect 851 687 885 691
rect 851 623 885 649
rect 851 615 885 623
rect 851 555 885 577
rect 851 543 885 555
rect 851 487 885 505
rect 851 471 885 487
rect 1014 1839 1048 1873
rect 1014 1779 1048 1801
rect 1014 1767 1048 1779
rect 1014 1711 1048 1729
rect 1014 1695 1048 1711
rect 1014 1643 1048 1657
rect 1014 1623 1048 1643
rect 1014 1575 1048 1585
rect 1014 1551 1048 1575
rect 1014 1507 1048 1513
rect 1014 1479 1048 1507
rect 1014 1439 1048 1441
rect 1014 1407 1048 1439
rect 1014 1337 1048 1369
rect 1014 1335 1048 1337
rect 1014 1269 1048 1297
rect 1014 1263 1048 1269
rect 1014 1201 1048 1225
rect 1014 1191 1048 1201
rect 1014 1133 1048 1153
rect 1014 1119 1048 1133
rect 1014 1065 1048 1081
rect 1014 1047 1048 1065
rect 1014 997 1048 1009
rect 1014 975 1048 997
rect 1014 929 1048 937
rect 1014 903 1048 929
rect 1014 861 1048 865
rect 1014 831 1048 861
rect 1014 759 1048 793
rect 1014 691 1048 721
rect 1014 687 1048 691
rect 1014 623 1048 649
rect 1014 615 1048 623
rect 1014 555 1048 577
rect 1014 543 1048 555
rect 1014 487 1048 505
rect 1014 471 1048 487
rect 1177 1839 1211 1873
rect 1177 1779 1211 1801
rect 1177 1767 1211 1779
rect 1177 1711 1211 1729
rect 1177 1695 1211 1711
rect 1177 1643 1211 1657
rect 1177 1623 1211 1643
rect 1177 1575 1211 1585
rect 1177 1551 1211 1575
rect 1177 1507 1211 1513
rect 1177 1479 1211 1507
rect 1177 1439 1211 1441
rect 1177 1407 1211 1439
rect 1177 1337 1211 1369
rect 1177 1335 1211 1337
rect 1177 1269 1211 1297
rect 1177 1263 1211 1269
rect 1177 1201 1211 1225
rect 1177 1191 1211 1201
rect 1177 1133 1211 1153
rect 1177 1119 1211 1133
rect 1177 1065 1211 1081
rect 1177 1047 1211 1065
rect 1177 997 1211 1009
rect 1177 975 1211 997
rect 1177 929 1211 937
rect 1177 903 1211 929
rect 1177 861 1211 865
rect 1177 831 1211 861
rect 1177 759 1211 793
rect 1177 691 1211 721
rect 1177 687 1211 691
rect 1177 623 1211 649
rect 1177 615 1211 623
rect 1177 555 1211 577
rect 1177 543 1211 555
rect 1177 487 1211 505
rect 1177 471 1211 487
rect 1340 1839 1374 1873
rect 1340 1779 1374 1801
rect 1340 1767 1374 1779
rect 1340 1711 1374 1729
rect 1340 1695 1374 1711
rect 1340 1643 1374 1657
rect 1340 1623 1374 1643
rect 1340 1575 1374 1585
rect 1340 1551 1374 1575
rect 1340 1507 1374 1513
rect 1340 1479 1374 1507
rect 1340 1439 1374 1441
rect 1340 1407 1374 1439
rect 1340 1337 1374 1369
rect 1340 1335 1374 1337
rect 1340 1269 1374 1297
rect 1340 1263 1374 1269
rect 1340 1201 1374 1225
rect 1340 1191 1374 1201
rect 1340 1133 1374 1153
rect 1340 1119 1374 1133
rect 1340 1065 1374 1081
rect 1340 1047 1374 1065
rect 1340 997 1374 1009
rect 1340 975 1374 997
rect 1340 929 1374 937
rect 1340 903 1374 929
rect 1340 861 1374 865
rect 1340 831 1374 861
rect 1340 759 1374 793
rect 1340 691 1374 721
rect 1340 687 1374 691
rect 1340 623 1374 649
rect 1340 615 1374 623
rect 1340 555 1374 577
rect 1340 543 1374 555
rect 1340 487 1374 505
rect 1340 471 1374 487
rect 1487 1857 1493 1882
rect 1493 1857 1521 1882
rect 1487 1848 1521 1857
rect 1487 1789 1493 1809
rect 1493 1789 1521 1809
rect 1487 1775 1521 1789
rect 1487 1721 1493 1736
rect 1493 1721 1521 1736
rect 1487 1702 1521 1721
rect 1487 1653 1493 1663
rect 1493 1653 1521 1663
rect 1487 1629 1521 1653
rect 1487 1585 1493 1590
rect 1493 1585 1521 1590
rect 1487 1556 1521 1585
rect 1487 1483 1521 1517
rect 1487 1415 1521 1444
rect 1487 1410 1493 1415
rect 1493 1410 1521 1415
rect 1487 1347 1521 1371
rect 1487 1337 1493 1347
rect 1493 1337 1521 1347
rect 1487 1279 1521 1298
rect 1487 1264 1493 1279
rect 1493 1264 1521 1279
rect 1487 1211 1521 1225
rect 1487 1191 1493 1211
rect 1493 1191 1521 1211
rect 1487 1143 1521 1151
rect 1487 1117 1493 1143
rect 1493 1117 1521 1143
rect 1487 1075 1521 1077
rect 1487 1043 1493 1075
rect 1493 1043 1521 1075
rect 1487 973 1493 1003
rect 1493 973 1521 1003
rect 1487 969 1521 973
rect 1487 905 1493 929
rect 1493 905 1521 929
rect 1487 895 1521 905
rect 1487 837 1493 855
rect 1493 837 1521 855
rect 1487 821 1521 837
rect 1487 769 1493 781
rect 1493 769 1521 781
rect 1487 747 1521 769
rect 1487 701 1493 707
rect 1493 701 1521 707
rect 1487 673 1521 701
rect 1487 599 1521 633
rect 1487 531 1521 559
rect 1487 525 1493 531
rect 1493 525 1521 531
rect 1487 463 1521 485
rect 1487 451 1493 463
rect 1493 451 1521 463
rect 253 333 287 367
rect 347 361 373 367
rect 373 361 381 367
rect 440 361 441 367
rect 441 361 474 367
rect 533 361 543 367
rect 543 361 567 367
rect 609 361 611 367
rect 611 361 643 367
rect 685 361 713 367
rect 713 361 719 367
rect 761 361 781 367
rect 781 361 795 367
rect 837 361 849 367
rect 849 361 871 367
rect 913 361 917 367
rect 917 361 947 367
rect 989 361 1019 367
rect 1019 361 1023 367
rect 1065 361 1087 367
rect 1087 361 1099 367
rect 1140 361 1155 367
rect 1155 361 1174 367
rect 1215 361 1223 367
rect 1223 361 1249 367
rect 1290 361 1291 367
rect 1291 361 1324 367
rect 1487 377 1521 411
rect 347 333 381 361
rect 440 333 474 361
rect 533 333 567 361
rect 609 333 643 361
rect 685 333 719 361
rect 761 333 795 361
rect 837 333 871 361
rect 913 333 947 361
rect 989 333 1023 361
rect 1065 333 1099 361
rect 1140 333 1174 361
rect 1215 333 1249 361
rect 1290 333 1324 361
rect 1365 333 1399 367
rect 1648 2226 1898 2228
rect 1648 2192 1682 2226
rect 1682 2192 1720 2226
rect 1720 2192 1754 2226
rect 1754 2192 1792 2226
rect 1792 2192 1826 2226
rect 1826 2192 1864 2226
rect 1864 2192 1898 2226
rect 1648 2158 1898 2192
rect 1648 2124 1682 2158
rect 1682 2124 1720 2158
rect 1720 2124 1754 2158
rect 1754 2124 1792 2158
rect 1792 2124 1826 2158
rect 1826 2124 1864 2158
rect 1864 2124 1898 2158
rect 1648 2090 1898 2124
rect 1648 2056 1682 2090
rect 1682 2056 1720 2090
rect 1720 2056 1754 2090
rect 1754 2056 1792 2090
rect 1792 2056 1826 2090
rect 1826 2056 1864 2090
rect 1864 2056 1898 2090
rect 1648 2022 1898 2056
rect 1648 1988 1682 2022
rect 1682 1988 1720 2022
rect 1720 1988 1754 2022
rect 1754 1988 1792 2022
rect 1792 1988 1826 2022
rect 1826 1988 1864 2022
rect 1864 1988 1898 2022
rect 1648 1954 1898 1988
rect 1648 1920 1682 1954
rect 1682 1920 1720 1954
rect 1720 1920 1754 1954
rect 1754 1920 1792 1954
rect 1792 1920 1826 1954
rect 1826 1920 1864 1954
rect 1864 1920 1898 1954
rect 1648 1886 1898 1920
rect 1648 1852 1682 1886
rect 1682 1852 1720 1886
rect 1720 1852 1754 1886
rect 1754 1852 1792 1886
rect 1792 1852 1826 1886
rect 1826 1852 1864 1886
rect 1864 1852 1898 1886
rect 1648 1818 1898 1852
rect 1648 1784 1682 1818
rect 1682 1784 1720 1818
rect 1720 1784 1754 1818
rect 1754 1784 1792 1818
rect 1792 1784 1826 1818
rect 1826 1784 1864 1818
rect 1864 1784 1898 1818
rect 1648 1750 1898 1784
rect 1648 1716 1682 1750
rect 1682 1716 1720 1750
rect 1720 1716 1754 1750
rect 1754 1716 1792 1750
rect 1792 1716 1826 1750
rect 1826 1716 1864 1750
rect 1864 1716 1898 1750
rect 1648 1682 1898 1716
rect 1648 1648 1682 1682
rect 1682 1648 1720 1682
rect 1720 1648 1754 1682
rect 1754 1648 1792 1682
rect 1792 1648 1826 1682
rect 1826 1648 1864 1682
rect 1864 1648 1898 1682
rect 1648 1614 1898 1648
rect 1648 1580 1682 1614
rect 1682 1580 1720 1614
rect 1720 1580 1754 1614
rect 1754 1580 1792 1614
rect 1792 1580 1826 1614
rect 1826 1580 1864 1614
rect 1864 1580 1898 1614
rect 1648 1546 1898 1580
rect 1648 1512 1682 1546
rect 1682 1512 1720 1546
rect 1720 1512 1754 1546
rect 1754 1512 1792 1546
rect 1792 1512 1826 1546
rect 1826 1512 1864 1546
rect 1864 1512 1898 1546
rect 1648 1478 1898 1512
rect 1648 1444 1682 1478
rect 1682 1444 1720 1478
rect 1720 1444 1754 1478
rect 1754 1444 1792 1478
rect 1792 1444 1826 1478
rect 1826 1444 1864 1478
rect 1864 1444 1898 1478
rect 1648 1410 1898 1444
rect 1648 1376 1682 1410
rect 1682 1376 1720 1410
rect 1720 1376 1754 1410
rect 1754 1376 1792 1410
rect 1792 1376 1826 1410
rect 1826 1376 1864 1410
rect 1864 1376 1898 1410
rect 1648 1342 1898 1376
rect 1648 1308 1682 1342
rect 1682 1308 1720 1342
rect 1720 1308 1754 1342
rect 1754 1308 1792 1342
rect 1792 1308 1826 1342
rect 1826 1308 1864 1342
rect 1864 1308 1898 1342
rect 1648 1274 1898 1308
rect 1648 1240 1682 1274
rect 1682 1240 1720 1274
rect 1720 1240 1754 1274
rect 1754 1240 1792 1274
rect 1792 1240 1826 1274
rect 1826 1240 1864 1274
rect 1864 1240 1898 1274
rect 1648 1206 1898 1240
rect 1648 1172 1682 1206
rect 1682 1172 1720 1206
rect 1720 1172 1754 1206
rect 1754 1172 1792 1206
rect 1792 1172 1826 1206
rect 1826 1172 1864 1206
rect 1864 1172 1898 1206
rect 1648 1138 1898 1172
rect 1648 1104 1682 1138
rect 1682 1104 1720 1138
rect 1720 1104 1754 1138
rect 1754 1104 1792 1138
rect 1792 1104 1826 1138
rect 1826 1104 1864 1138
rect 1864 1104 1898 1138
rect 1648 1070 1898 1104
rect 1648 1036 1682 1070
rect 1682 1036 1720 1070
rect 1720 1036 1754 1070
rect 1754 1036 1792 1070
rect 1792 1036 1826 1070
rect 1826 1036 1864 1070
rect 1864 1036 1898 1070
rect 1648 1002 1898 1036
rect 1648 968 1682 1002
rect 1682 968 1720 1002
rect 1720 968 1754 1002
rect 1754 968 1792 1002
rect 1792 968 1826 1002
rect 1826 968 1864 1002
rect 1864 968 1898 1002
rect 1648 934 1898 968
rect 1648 900 1682 934
rect 1682 900 1720 934
rect 1720 900 1754 934
rect 1754 900 1792 934
rect 1792 900 1826 934
rect 1826 900 1864 934
rect 1864 900 1898 934
rect 1648 866 1898 900
rect 1648 832 1682 866
rect 1682 832 1720 866
rect 1720 832 1754 866
rect 1754 832 1792 866
rect 1792 832 1826 866
rect 1826 832 1864 866
rect 1864 832 1898 866
rect 1648 798 1898 832
rect 1648 764 1682 798
rect 1682 764 1720 798
rect 1720 764 1754 798
rect 1754 764 1792 798
rect 1792 764 1826 798
rect 1826 764 1864 798
rect 1864 764 1898 798
rect 1648 754 1898 764
rect 3469 2250 3503 2260
rect 3469 2178 3503 2210
rect 3469 2176 3503 2178
rect 1648 696 1682 715
rect 1648 681 1682 696
rect 1720 696 1754 715
rect 1720 681 1754 696
rect 1792 696 1826 715
rect 1792 681 1826 696
rect 1864 696 1898 715
rect 1864 681 1898 696
rect 1648 628 1682 642
rect 1648 608 1682 628
rect 1720 628 1754 642
rect 1720 608 1754 628
rect 1792 628 1826 642
rect 1792 608 1826 628
rect 1864 628 1898 642
rect 1864 608 1898 628
rect 1648 560 1682 569
rect 1648 535 1682 560
rect 1720 560 1754 569
rect 1720 535 1754 560
rect 1792 560 1826 569
rect 1792 535 1826 560
rect 1864 560 1898 569
rect 1864 535 1898 560
rect 1648 492 1682 496
rect 1648 462 1682 492
rect 1720 492 1754 496
rect 1720 462 1754 492
rect 1792 492 1826 496
rect 1792 462 1826 492
rect 1864 492 1898 496
rect 1864 462 1898 492
rect 1648 390 1682 423
rect 1648 389 1682 390
rect 1720 390 1754 423
rect 1720 389 1754 390
rect 1792 390 1826 423
rect 1792 389 1826 390
rect 1864 390 1898 423
rect 1864 389 1898 390
rect 10 262 44 296
rect 10 211 44 222
rect 10 188 44 211
rect 10 114 44 148
rect 1648 322 1682 350
rect 1648 316 1682 322
rect 1720 322 1754 350
rect 1720 316 1754 322
rect 1792 322 1826 350
rect 1792 316 1826 322
rect 1864 322 1898 350
rect 1864 316 1898 322
rect 2212 2039 2246 2073
rect 2286 2039 2320 2073
rect 2360 2039 2394 2073
rect 2434 2039 2468 2073
rect 2508 2039 2542 2073
rect 2582 2039 2616 2073
rect 2656 2039 2690 2073
rect 2730 2039 2764 2073
rect 2804 2039 2838 2073
rect 2878 2039 2912 2073
rect 2952 2039 2986 2073
rect 3026 2039 3060 2073
rect 3101 2039 3106 2073
rect 3106 2039 3135 2073
rect 3176 2039 3210 2073
rect 2092 2005 2120 2029
rect 2120 2005 2126 2029
rect 2092 1995 2126 2005
rect 2092 1921 2126 1955
rect 2303 1923 2307 1957
rect 2307 1923 2337 1957
rect 2382 1923 2410 1957
rect 2410 1923 2416 1957
rect 2461 1923 2479 1957
rect 2479 1923 2495 1957
rect 2540 1923 2548 1957
rect 2548 1923 2574 1957
rect 2619 1923 2652 1957
rect 2652 1923 2653 1957
rect 2697 1923 2721 1957
rect 2721 1923 2731 1957
rect 2775 1923 2789 1957
rect 2789 1923 2809 1957
rect 2853 1923 2857 1957
rect 2857 1923 2887 1957
rect 2931 1923 2959 1957
rect 2959 1923 2965 1957
rect 3009 1923 3027 1957
rect 3027 1923 3043 1957
rect 2092 1847 2126 1881
rect 3220 1921 3254 1955
rect 2092 1773 2126 1807
rect 2092 1699 2126 1733
rect 2092 1625 2126 1659
rect 2092 1551 2126 1585
rect 2092 1477 2126 1511
rect 2092 1403 2126 1437
rect 2092 1329 2126 1363
rect 2092 1255 2126 1289
rect 2092 1181 2126 1215
rect 2092 1108 2126 1142
rect 2092 1035 2126 1069
rect 2092 962 2126 996
rect 2092 889 2126 923
rect 2092 816 2126 850
rect 2092 743 2126 777
rect 2092 670 2126 704
rect 2092 597 2126 631
rect 2092 524 2126 558
rect 2092 451 2126 485
rect 2246 1839 2280 1873
rect 2246 1779 2280 1801
rect 2246 1767 2280 1779
rect 2246 1711 2280 1729
rect 2246 1695 2280 1711
rect 2246 1643 2280 1657
rect 2246 1623 2280 1643
rect 2246 1575 2280 1585
rect 2246 1551 2280 1575
rect 2246 1507 2280 1513
rect 2246 1479 2280 1507
rect 2246 1439 2280 1441
rect 2246 1407 2280 1439
rect 2246 1337 2280 1369
rect 2246 1335 2280 1337
rect 2246 1269 2280 1297
rect 2246 1263 2280 1269
rect 2246 1201 2280 1225
rect 2246 1191 2280 1201
rect 2246 1133 2280 1153
rect 2246 1119 2280 1133
rect 2246 1065 2280 1081
rect 2246 1047 2280 1065
rect 2246 997 2280 1009
rect 2246 975 2280 997
rect 2246 929 2280 937
rect 2246 903 2280 929
rect 2246 861 2280 865
rect 2246 831 2280 861
rect 2246 759 2280 793
rect 2246 691 2280 721
rect 2246 687 2280 691
rect 2246 623 2280 649
rect 2246 615 2280 623
rect 2246 555 2280 577
rect 2246 543 2280 555
rect 2246 487 2280 505
rect 2246 471 2280 487
rect 2409 1839 2443 1873
rect 2409 1779 2443 1801
rect 2409 1767 2443 1779
rect 2409 1711 2443 1729
rect 2409 1695 2443 1711
rect 2409 1643 2443 1657
rect 2409 1623 2443 1643
rect 2409 1575 2443 1585
rect 2409 1551 2443 1575
rect 2409 1507 2443 1513
rect 2409 1479 2443 1507
rect 2409 1439 2443 1441
rect 2409 1407 2443 1439
rect 2409 1337 2443 1369
rect 2409 1335 2443 1337
rect 2409 1269 2443 1297
rect 2409 1263 2443 1269
rect 2409 1201 2443 1225
rect 2409 1191 2443 1201
rect 2409 1133 2443 1153
rect 2409 1119 2443 1133
rect 2409 1065 2443 1081
rect 2409 1047 2443 1065
rect 2409 997 2443 1009
rect 2409 975 2443 997
rect 2409 929 2443 937
rect 2409 903 2443 929
rect 2409 861 2443 865
rect 2409 831 2443 861
rect 2409 759 2443 793
rect 2409 691 2443 721
rect 2409 687 2443 691
rect 2409 623 2443 649
rect 2409 615 2443 623
rect 2409 555 2443 577
rect 2409 543 2443 555
rect 2409 487 2443 505
rect 2409 471 2443 487
rect 2572 1839 2606 1873
rect 2572 1779 2606 1801
rect 2572 1767 2606 1779
rect 2572 1711 2606 1729
rect 2572 1695 2606 1711
rect 2572 1643 2606 1657
rect 2572 1623 2606 1643
rect 2572 1575 2606 1585
rect 2572 1551 2606 1575
rect 2572 1507 2606 1513
rect 2572 1479 2606 1507
rect 2572 1439 2606 1441
rect 2572 1407 2606 1439
rect 2572 1337 2606 1369
rect 2572 1335 2606 1337
rect 2572 1269 2606 1297
rect 2572 1263 2606 1269
rect 2572 1201 2606 1225
rect 2572 1191 2606 1201
rect 2572 1133 2606 1153
rect 2572 1119 2606 1133
rect 2572 1065 2606 1081
rect 2572 1047 2606 1065
rect 2572 997 2606 1009
rect 2572 975 2606 997
rect 2572 929 2606 937
rect 2572 903 2606 929
rect 2572 861 2606 865
rect 2572 831 2606 861
rect 2572 759 2606 793
rect 2572 691 2606 721
rect 2572 687 2606 691
rect 2572 623 2606 649
rect 2572 615 2606 623
rect 2572 555 2606 577
rect 2572 543 2606 555
rect 2572 487 2606 505
rect 2572 471 2606 487
rect 2735 1839 2769 1873
rect 2735 1779 2769 1801
rect 2735 1767 2769 1779
rect 2735 1711 2769 1729
rect 2735 1695 2769 1711
rect 2735 1643 2769 1657
rect 2735 1623 2769 1643
rect 2735 1575 2769 1585
rect 2735 1551 2769 1575
rect 2735 1507 2769 1513
rect 2735 1479 2769 1507
rect 2735 1439 2769 1441
rect 2735 1407 2769 1439
rect 2735 1337 2769 1369
rect 2735 1335 2769 1337
rect 2735 1269 2769 1297
rect 2735 1263 2769 1269
rect 2735 1201 2769 1225
rect 2735 1191 2769 1201
rect 2735 1133 2769 1153
rect 2735 1119 2769 1133
rect 2735 1065 2769 1081
rect 2735 1047 2769 1065
rect 2735 997 2769 1009
rect 2735 975 2769 997
rect 2735 929 2769 937
rect 2735 903 2769 929
rect 2735 861 2769 865
rect 2735 831 2769 861
rect 2735 759 2769 793
rect 2735 691 2769 721
rect 2735 687 2769 691
rect 2735 623 2769 649
rect 2735 615 2769 623
rect 2735 555 2769 577
rect 2735 543 2769 555
rect 2735 487 2769 505
rect 2735 471 2769 487
rect 2898 1839 2932 1873
rect 2898 1779 2932 1801
rect 2898 1767 2932 1779
rect 2898 1711 2932 1729
rect 2898 1695 2932 1711
rect 2898 1643 2932 1657
rect 2898 1623 2932 1643
rect 2898 1575 2932 1585
rect 2898 1551 2932 1575
rect 2898 1507 2932 1513
rect 2898 1479 2932 1507
rect 2898 1439 2932 1441
rect 2898 1407 2932 1439
rect 2898 1337 2932 1369
rect 2898 1335 2932 1337
rect 2898 1269 2932 1297
rect 2898 1263 2932 1269
rect 2898 1201 2932 1225
rect 2898 1191 2932 1201
rect 2898 1133 2932 1153
rect 2898 1119 2932 1133
rect 2898 1065 2932 1081
rect 2898 1047 2932 1065
rect 2898 997 2932 1009
rect 2898 975 2932 997
rect 2898 929 2932 937
rect 2898 903 2932 929
rect 2898 861 2932 865
rect 2898 831 2932 861
rect 2898 759 2932 793
rect 2898 691 2932 721
rect 2898 687 2932 691
rect 2898 623 2932 649
rect 2898 615 2932 623
rect 2898 555 2932 577
rect 2898 543 2932 555
rect 2898 487 2932 505
rect 2898 471 2932 487
rect 3061 1839 3095 1873
rect 3061 1779 3095 1801
rect 3061 1767 3095 1779
rect 3061 1711 3095 1729
rect 3061 1695 3095 1711
rect 3061 1643 3095 1657
rect 3061 1623 3095 1643
rect 3061 1575 3095 1585
rect 3061 1551 3095 1575
rect 3061 1507 3095 1513
rect 3061 1479 3095 1507
rect 3061 1439 3095 1441
rect 3061 1407 3095 1439
rect 3061 1337 3095 1369
rect 3061 1335 3095 1337
rect 3061 1269 3095 1297
rect 3061 1263 3095 1269
rect 3061 1201 3095 1225
rect 3061 1191 3095 1201
rect 3061 1133 3095 1153
rect 3061 1119 3095 1133
rect 3061 1065 3095 1081
rect 3061 1047 3095 1065
rect 3061 997 3095 1009
rect 3061 975 3095 997
rect 3061 929 3095 937
rect 3061 903 3095 929
rect 3061 861 3095 865
rect 3061 831 3095 861
rect 3061 759 3095 793
rect 3061 691 3095 721
rect 3061 687 3095 691
rect 3061 623 3095 649
rect 3061 615 3095 623
rect 3061 555 3095 577
rect 3061 543 3095 555
rect 3061 487 3095 505
rect 3061 471 3095 487
rect 3220 1848 3254 1882
rect 3220 1775 3254 1809
rect 3220 1702 3254 1736
rect 3220 1629 3254 1663
rect 3220 1556 3254 1590
rect 3220 1483 3254 1517
rect 3220 1410 3254 1444
rect 3220 1337 3254 1371
rect 3220 1264 3254 1298
rect 3220 1191 3254 1225
rect 3220 1117 3254 1151
rect 3220 1043 3254 1077
rect 3220 985 3254 1003
rect 3220 969 3254 985
rect 3220 910 3254 929
rect 3220 895 3254 910
rect 3220 821 3254 855
rect 3220 747 3254 781
rect 3220 673 3254 707
rect 3220 599 3254 633
rect 3220 525 3254 559
rect 3220 468 3254 485
rect 3220 451 3254 468
rect 3220 400 3248 411
rect 3248 400 3254 411
rect 3220 377 3254 400
rect 2136 359 2154 367
rect 2154 359 2170 367
rect 2136 333 2170 359
rect 2230 333 2264 367
rect 2323 333 2357 367
rect 2416 333 2450 367
rect 2492 333 2526 367
rect 2568 333 2602 367
rect 2644 333 2678 367
rect 2720 333 2754 367
rect 2796 333 2830 367
rect 2872 333 2906 367
rect 2948 333 2982 367
rect 3023 333 3057 367
rect 3098 333 3132 367
rect 3469 2102 3503 2136
rect 3469 2028 3503 2062
rect 3469 1954 3503 1988
rect 3469 1880 3503 1914
rect 3469 1806 3503 1840
rect 3469 1732 3503 1766
rect 3469 1658 3503 1692
rect 3469 1584 3503 1618
rect 3469 1510 3503 1544
rect 3469 1436 3503 1470
rect 3469 1362 3503 1396
rect 3469 1288 3503 1322
rect 3469 1214 3503 1248
rect 3469 1140 3503 1174
rect 3469 1066 3503 1100
rect 3469 992 3503 1026
rect 3469 918 3503 952
rect 3469 845 3503 879
rect 3469 772 3503 806
rect 3469 699 3503 733
rect 3469 626 3503 660
rect 3469 553 3503 587
rect 3469 480 3503 514
rect 3469 407 3503 441
rect 3469 334 3503 368
rect 1648 254 1682 277
rect 1648 243 1682 254
rect 1720 254 1754 277
rect 1720 243 1754 254
rect 1792 254 1826 277
rect 1792 243 1826 254
rect 1864 254 1898 277
rect 1864 243 1898 254
rect 1648 170 1682 204
rect 1720 170 1754 204
rect 1792 170 1826 204
rect 1864 170 1898 204
rect 3469 261 3503 295
rect 3469 188 3503 222
rect 128 70 162 104
rect 201 70 235 104
rect 274 70 308 104
rect 347 70 381 104
rect 420 70 454 104
rect 493 70 527 104
rect 566 70 600 104
rect 639 70 673 104
rect 712 70 746 104
rect 785 70 819 104
rect 858 70 892 104
rect 931 70 965 104
rect 1004 70 1038 104
rect 1077 70 1111 104
rect 1150 70 1184 104
rect 1223 70 1257 104
rect 1296 70 1330 104
rect 1369 70 1403 104
rect 1442 70 1476 104
rect 1515 70 1549 104
rect 1588 70 1622 104
rect 1661 70 1695 104
rect 1734 70 1768 104
rect 1807 70 1841 104
rect 1880 70 1914 104
rect 1953 70 1987 104
rect 2026 70 2060 104
rect 2099 70 2133 104
rect 2172 70 2206 104
rect 2245 70 2279 104
rect 2318 70 2352 104
rect 2391 70 2425 104
rect 2464 70 2498 104
rect 2537 70 2571 104
rect 2611 70 2645 104
rect 2685 70 2719 104
rect 2759 70 2793 104
rect 2833 70 2867 104
rect 2907 70 2941 104
rect 2981 70 3015 104
rect 3055 70 3089 104
rect 3129 70 3163 104
rect 3203 70 3237 104
rect 3277 70 3311 104
rect 3351 70 3385 104
rect 3425 70 3459 104
rect 3828 2294 3862 2328
rect 3922 2294 3956 2328
rect 4015 2294 4049 2328
rect 4108 2294 4142 2328
rect 4184 2294 4218 2328
rect 4258 2294 4292 2328
rect 4332 2294 4366 2328
rect 4406 2294 4440 2328
rect 4480 2294 4514 2328
rect 4554 2294 4588 2328
rect 4628 2294 4662 2328
rect 4702 2294 4736 2328
rect 4776 2294 4810 2328
rect 4850 2294 4884 2328
rect 4924 2294 4958 2328
rect 4998 2294 5032 2328
rect 5072 2294 5106 2328
rect 5146 2294 5180 2328
rect 5220 2294 5254 2328
rect 5294 2294 5328 2328
rect 5368 2294 5402 2328
rect 5442 2294 5476 2328
rect 5516 2294 5550 2328
rect 5590 2294 5624 2328
rect 5663 2294 5697 2328
rect 5736 2294 5770 2328
rect 5809 2294 5843 2328
rect 5882 2294 5916 2328
rect 5955 2294 5989 2328
rect 6028 2294 6062 2328
rect 6101 2294 6135 2328
rect 6174 2294 6208 2328
rect 6247 2294 6281 2328
rect 6320 2294 6354 2328
rect 6393 2294 6427 2328
rect 6466 2294 6500 2328
rect 6539 2294 6573 2328
rect 6612 2294 6646 2328
rect 6685 2294 6719 2328
rect 6758 2294 6792 2328
rect 6956 2294 6990 2328
rect 7028 2294 7062 2328
rect 7100 2294 7134 2328
rect 7172 2294 7206 2328
rect 7244 2294 7278 2328
rect 7316 2294 7350 2328
rect 7388 2294 7422 2328
rect 7460 2294 7494 2328
rect 7532 2294 7566 2328
rect 7604 2294 7638 2328
rect 7676 2294 7710 2328
rect 7748 2294 7782 2328
rect 7820 2294 7854 2328
rect 7892 2294 7926 2328
rect 7964 2294 7998 2328
rect 8036 2294 8070 2328
rect 8108 2294 8142 2328
rect 8181 2294 8215 2328
rect 8254 2294 8288 2328
rect 8327 2294 8361 2328
rect 8400 2294 8434 2328
rect 8473 2294 8507 2328
rect 8546 2294 8580 2328
rect 8619 2294 8653 2328
rect 8692 2294 8726 2328
rect 8765 2294 8799 2328
rect 8838 2294 8872 2328
rect 8911 2294 8945 2328
rect 8984 2294 9018 2328
rect 9057 2294 9091 2328
rect 9133 2294 9167 2328
rect 9205 2294 9239 2328
rect 9277 2294 9311 2328
rect 9349 2294 9383 2328
rect 9421 2294 9455 2328
rect 9493 2294 9527 2328
rect 9565 2294 9599 2328
rect 9637 2294 9671 2328
rect 9709 2294 9743 2328
rect 9781 2294 9815 2328
rect 9853 2294 9887 2328
rect 9926 2294 9960 2328
rect 9999 2294 10033 2328
rect 10072 2294 10106 2328
rect 10145 2294 10179 2328
rect 3784 2186 3818 2210
rect 3784 2176 3818 2186
rect 3784 2103 3818 2137
rect 6876 2250 6910 2284
rect 6876 2176 6910 2210
rect 6876 2102 6910 2136
rect 10189 2178 10223 2212
rect 3784 2030 3818 2064
rect 3784 1957 3818 1991
rect 3784 1884 3818 1918
rect 3784 1811 3818 1845
rect 3784 1738 3818 1772
rect 3784 1665 3818 1699
rect 3784 1592 3818 1626
rect 3784 1519 3818 1553
rect 3784 1446 3818 1480
rect 3784 1373 3818 1407
rect 3784 1300 3818 1334
rect 3784 1227 3818 1261
rect 3784 1154 3818 1188
rect 3784 1081 3818 1115
rect 3784 1008 3818 1042
rect 3784 935 3818 969
rect 3784 862 3818 896
rect 3784 788 3818 822
rect 3784 714 3818 748
rect 3784 640 3818 674
rect 3784 566 3818 600
rect 3784 492 3818 526
rect 3784 418 3818 452
rect 3784 344 3818 378
rect 4099 2039 4133 2073
rect 4179 2039 4207 2073
rect 4207 2039 4213 2073
rect 4252 2039 4275 2073
rect 4275 2039 4286 2073
rect 4325 2039 4343 2073
rect 4343 2039 4359 2073
rect 4398 2039 4411 2073
rect 4411 2039 4432 2073
rect 4471 2039 4479 2073
rect 4479 2039 4505 2073
rect 4544 2039 4547 2073
rect 4547 2039 4578 2073
rect 4617 2039 4649 2073
rect 4649 2039 4651 2073
rect 4690 2039 4717 2073
rect 4717 2039 4724 2073
rect 4763 2039 4785 2073
rect 4785 2039 4797 2073
rect 4836 2039 4853 2073
rect 4853 2039 4870 2073
rect 4909 2039 4921 2073
rect 4921 2039 4943 2073
rect 4982 2039 4989 2073
rect 4989 2039 5016 2073
rect 5055 2039 5057 2073
rect 5057 2039 5089 2073
rect 5128 2039 5159 2073
rect 5159 2039 5162 2073
rect 5201 2039 5227 2073
rect 5227 2039 5235 2073
rect 5274 2039 5295 2073
rect 5295 2039 5308 2073
rect 5347 2039 5363 2073
rect 5363 2039 5381 2073
rect 5420 2039 5431 2073
rect 5431 2039 5454 2073
rect 5493 2039 5499 2073
rect 5499 2039 5527 2073
rect 5566 2039 5567 2073
rect 5567 2039 5600 2073
rect 5639 2039 5669 2073
rect 5669 2039 5673 2073
rect 5712 2039 5737 2073
rect 5737 2039 5746 2073
rect 5785 2039 5805 2073
rect 5805 2039 5819 2073
rect 5858 2039 5873 2073
rect 5873 2039 5892 2073
rect 5931 2039 5941 2073
rect 5941 2039 5965 2073
rect 6004 2039 6009 2073
rect 6009 2039 6038 2073
rect 6077 2039 6111 2073
rect 6150 2039 6179 2073
rect 6179 2039 6184 2073
rect 6223 2039 6247 2073
rect 6247 2039 6257 2073
rect 6295 2039 6315 2073
rect 6315 2039 6329 2073
rect 6367 2039 6383 2073
rect 6383 2039 6401 2073
rect 6439 2039 6451 2073
rect 6451 2039 6473 2073
rect 6511 2039 6519 2073
rect 6519 2039 6545 2073
rect 6583 2039 6587 2073
rect 6587 2039 6617 2073
rect 4005 1971 4039 1999
rect 4005 1965 4039 1971
rect 6655 1999 6689 2001
rect 6655 1967 6689 1999
rect 4005 1903 4039 1925
rect 4176 1923 4192 1957
rect 4192 1923 4210 1957
rect 4250 1923 4264 1957
rect 4264 1923 4284 1957
rect 4323 1923 4336 1957
rect 4336 1923 4357 1957
rect 4396 1923 4408 1957
rect 4408 1923 4430 1957
rect 4469 1923 4480 1957
rect 4480 1923 4503 1957
rect 4542 1923 4552 1957
rect 4552 1923 4576 1957
rect 4615 1923 4624 1957
rect 4624 1923 4649 1957
rect 4688 1923 4696 1957
rect 4696 1923 4722 1957
rect 5459 1923 5463 1957
rect 5463 1923 5493 1957
rect 5535 1923 5536 1957
rect 5536 1923 5569 1957
rect 5611 1923 5643 1957
rect 5643 1923 5645 1957
rect 5687 1923 5716 1957
rect 5716 1923 5721 1957
rect 5763 1923 5789 1957
rect 5789 1923 5797 1957
rect 5838 1923 5861 1957
rect 5861 1923 5872 1957
rect 5913 1923 5933 1957
rect 5933 1923 5947 1957
rect 5988 1923 6005 1957
rect 6005 1923 6022 1957
rect 4005 1891 4039 1903
rect 6655 1897 6689 1926
rect 6655 1892 6689 1897
rect 4005 1835 4039 1851
rect 4005 1817 4039 1835
rect 4005 1767 4039 1777
rect 4005 1743 4039 1767
rect 4005 1699 4039 1703
rect 4005 1669 4039 1699
rect 4005 1597 4039 1629
rect 4005 1595 4039 1597
rect 4005 1529 4039 1555
rect 4005 1521 4039 1529
rect 4005 1461 4039 1481
rect 4005 1447 4039 1461
rect 4005 1393 4039 1407
rect 4005 1373 4039 1393
rect 4005 1325 4039 1333
rect 4005 1299 4039 1325
rect 4005 1257 4039 1259
rect 4005 1225 4039 1257
rect 4005 1155 4039 1185
rect 4005 1151 4039 1155
rect 4005 1087 4039 1111
rect 4005 1077 4039 1087
rect 4005 1019 4039 1037
rect 4005 1003 4039 1019
rect 4005 951 4039 963
rect 4005 929 4039 951
rect 4005 883 4039 889
rect 4005 855 4039 883
rect 4005 781 4039 814
rect 4005 780 4039 781
rect 4005 713 4039 739
rect 4005 705 4039 713
rect 4005 645 4039 664
rect 4005 630 4039 645
rect 4005 555 4039 589
rect 4005 486 4039 514
rect 4005 480 4039 486
rect 4131 1839 4165 1873
rect 4131 1779 4165 1801
rect 4131 1767 4165 1779
rect 4131 1711 4165 1729
rect 4131 1695 4165 1711
rect 4131 1643 4165 1657
rect 4131 1623 4165 1643
rect 4131 1575 4165 1585
rect 4131 1551 4165 1575
rect 4131 1507 4165 1513
rect 4131 1479 4165 1507
rect 4131 1439 4165 1441
rect 4131 1407 4165 1439
rect 4131 1337 4165 1369
rect 4131 1335 4165 1337
rect 4131 1269 4165 1297
rect 4131 1263 4165 1269
rect 4131 1201 4165 1225
rect 4131 1191 4165 1201
rect 4131 1133 4165 1153
rect 4131 1119 4165 1133
rect 4131 1065 4165 1081
rect 4131 1047 4165 1065
rect 4131 997 4165 1009
rect 4131 975 4165 997
rect 4131 929 4165 937
rect 4131 903 4165 929
rect 4131 861 4165 865
rect 4131 831 4165 861
rect 4131 759 4165 793
rect 4131 691 4165 721
rect 4131 687 4165 691
rect 4131 623 4165 649
rect 4131 615 4165 623
rect 4131 555 4165 577
rect 4131 543 4165 555
rect 4131 487 4165 505
rect 4131 471 4165 487
rect 4294 1839 4328 1873
rect 4294 1779 4328 1801
rect 4294 1767 4328 1779
rect 4294 1711 4328 1729
rect 4294 1695 4328 1711
rect 4294 1643 4328 1657
rect 4294 1623 4328 1643
rect 4294 1575 4328 1585
rect 4294 1551 4328 1575
rect 4294 1507 4328 1513
rect 4294 1479 4328 1507
rect 4294 1439 4328 1441
rect 4294 1407 4328 1439
rect 4294 1337 4328 1369
rect 4294 1335 4328 1337
rect 4294 1269 4328 1297
rect 4294 1263 4328 1269
rect 4294 1201 4328 1225
rect 4294 1191 4328 1201
rect 4294 1133 4328 1153
rect 4294 1119 4328 1133
rect 4294 1065 4328 1081
rect 4294 1047 4328 1065
rect 4294 997 4328 1009
rect 4294 975 4328 997
rect 4294 929 4328 937
rect 4294 903 4328 929
rect 4294 861 4328 865
rect 4294 831 4328 861
rect 4294 759 4328 793
rect 4294 691 4328 721
rect 4294 687 4328 691
rect 4294 623 4328 649
rect 4294 615 4328 623
rect 4294 555 4328 577
rect 4294 543 4328 555
rect 4294 487 4328 505
rect 4294 471 4328 487
rect 4457 1839 4491 1873
rect 4457 1779 4491 1801
rect 4457 1767 4491 1779
rect 4457 1711 4491 1729
rect 4457 1695 4491 1711
rect 4457 1643 4491 1657
rect 4457 1623 4491 1643
rect 4457 1575 4491 1585
rect 4457 1551 4491 1575
rect 4457 1507 4491 1513
rect 4457 1479 4491 1507
rect 4457 1439 4491 1441
rect 4457 1407 4491 1439
rect 4457 1337 4491 1369
rect 4457 1335 4491 1337
rect 4457 1269 4491 1297
rect 4457 1263 4491 1269
rect 4457 1201 4491 1225
rect 4457 1191 4491 1201
rect 4457 1133 4491 1153
rect 4457 1119 4491 1133
rect 4457 1065 4491 1081
rect 4457 1047 4491 1065
rect 4457 997 4491 1009
rect 4457 975 4491 997
rect 4457 929 4491 937
rect 4457 903 4491 929
rect 4457 861 4491 865
rect 4457 831 4491 861
rect 4457 759 4491 793
rect 4457 691 4491 721
rect 4457 687 4491 691
rect 4457 623 4491 649
rect 4457 615 4491 623
rect 4457 555 4491 577
rect 4457 543 4491 555
rect 4457 487 4491 505
rect 4457 471 4491 487
rect 4620 1839 4654 1873
rect 4620 1779 4654 1801
rect 4620 1767 4654 1779
rect 4620 1711 4654 1729
rect 4620 1695 4654 1711
rect 4620 1643 4654 1657
rect 4620 1623 4654 1643
rect 4620 1575 4654 1585
rect 4620 1551 4654 1575
rect 4620 1507 4654 1513
rect 4620 1479 4654 1507
rect 4620 1439 4654 1441
rect 4620 1407 4654 1439
rect 4620 1337 4654 1369
rect 4620 1335 4654 1337
rect 4620 1269 4654 1297
rect 4620 1263 4654 1269
rect 4620 1201 4654 1225
rect 4620 1191 4654 1201
rect 4620 1133 4654 1153
rect 4620 1119 4654 1133
rect 4620 1065 4654 1081
rect 4620 1047 4654 1065
rect 4620 997 4654 1009
rect 4620 975 4654 997
rect 4620 929 4654 937
rect 4620 903 4654 929
rect 4620 861 4654 865
rect 4620 831 4654 861
rect 4620 759 4654 793
rect 4620 691 4654 721
rect 4620 687 4654 691
rect 4620 623 4654 649
rect 4620 615 4654 623
rect 4620 555 4654 577
rect 4620 543 4654 555
rect 4620 487 4654 505
rect 4620 471 4654 487
rect 4783 1839 4817 1873
rect 4783 1779 4817 1801
rect 4783 1767 4817 1779
rect 4783 1711 4817 1729
rect 4783 1695 4817 1711
rect 4783 1643 4817 1657
rect 4783 1623 4817 1643
rect 4783 1575 4817 1585
rect 4783 1551 4817 1575
rect 4783 1507 4817 1513
rect 4783 1479 4817 1507
rect 4783 1439 4817 1441
rect 4783 1407 4817 1439
rect 4783 1337 4817 1369
rect 4783 1335 4817 1337
rect 4783 1269 4817 1297
rect 4783 1263 4817 1269
rect 4783 1201 4817 1225
rect 4783 1191 4817 1201
rect 4783 1133 4817 1153
rect 4783 1119 4817 1133
rect 4783 1065 4817 1081
rect 4783 1047 4817 1065
rect 4783 997 4817 1009
rect 4783 975 4817 997
rect 4783 929 4817 937
rect 4783 903 4817 929
rect 4783 861 4817 865
rect 4783 831 4817 861
rect 4783 759 4817 793
rect 4783 691 4817 721
rect 4783 687 4817 691
rect 4783 623 4817 649
rect 4783 615 4817 623
rect 4783 555 4817 577
rect 4783 543 4817 555
rect 4783 487 4817 505
rect 4783 471 4817 487
rect 4946 1839 4980 1873
rect 4946 1779 4980 1801
rect 4946 1767 4980 1779
rect 4946 1711 4980 1729
rect 4946 1695 4980 1711
rect 4946 1643 4980 1657
rect 4946 1623 4980 1643
rect 4946 1575 4980 1585
rect 4946 1551 4980 1575
rect 4946 1507 4980 1513
rect 4946 1479 4980 1507
rect 4946 1439 4980 1441
rect 4946 1407 4980 1439
rect 4946 1337 4980 1369
rect 4946 1335 4980 1337
rect 4946 1269 4980 1297
rect 4946 1263 4980 1269
rect 4946 1201 4980 1225
rect 4946 1191 4980 1201
rect 4946 1133 4980 1153
rect 4946 1119 4980 1133
rect 4946 1065 4980 1081
rect 4946 1047 4980 1065
rect 4946 997 4980 1009
rect 4946 975 4980 997
rect 4946 929 4980 937
rect 4946 903 4980 929
rect 4946 861 4980 865
rect 4946 831 4980 861
rect 4946 759 4980 793
rect 4946 691 4980 721
rect 4946 687 4980 691
rect 4946 623 4980 649
rect 4946 615 4980 623
rect 4946 555 4980 577
rect 4946 543 4980 555
rect 4946 487 4980 505
rect 4946 471 4980 487
rect 5109 1839 5143 1873
rect 5109 1779 5143 1801
rect 5109 1767 5143 1779
rect 5109 1711 5143 1729
rect 5109 1695 5143 1711
rect 5109 1643 5143 1657
rect 5109 1623 5143 1643
rect 5109 1575 5143 1585
rect 5109 1551 5143 1575
rect 5109 1507 5143 1513
rect 5109 1479 5143 1507
rect 5109 1439 5143 1441
rect 5109 1407 5143 1439
rect 5109 1337 5143 1369
rect 5109 1335 5143 1337
rect 5109 1269 5143 1297
rect 5109 1263 5143 1269
rect 5109 1201 5143 1225
rect 5109 1191 5143 1201
rect 5109 1133 5143 1153
rect 5109 1119 5143 1133
rect 5109 1065 5143 1081
rect 5109 1047 5143 1065
rect 5109 997 5143 1009
rect 5109 975 5143 997
rect 5109 929 5143 937
rect 5109 903 5143 929
rect 5109 861 5143 865
rect 5109 831 5143 861
rect 5109 759 5143 793
rect 5109 691 5143 721
rect 5109 687 5143 691
rect 5109 623 5143 649
rect 5109 615 5143 623
rect 5109 555 5143 577
rect 5109 543 5143 555
rect 5109 487 5143 505
rect 5109 471 5143 487
rect 5272 1839 5306 1873
rect 5272 1779 5306 1801
rect 5272 1767 5306 1779
rect 5272 1711 5306 1729
rect 5272 1695 5306 1711
rect 5272 1643 5306 1657
rect 5272 1623 5306 1643
rect 5272 1575 5306 1585
rect 5272 1551 5306 1575
rect 5272 1507 5306 1513
rect 5272 1479 5306 1507
rect 5272 1439 5306 1441
rect 5272 1407 5306 1439
rect 5272 1337 5306 1369
rect 5272 1335 5306 1337
rect 5272 1269 5306 1297
rect 5272 1263 5306 1269
rect 5272 1201 5306 1225
rect 5272 1191 5306 1201
rect 5272 1133 5306 1153
rect 5272 1119 5306 1133
rect 5272 1065 5306 1081
rect 5272 1047 5306 1065
rect 5272 997 5306 1009
rect 5272 975 5306 997
rect 5272 929 5306 937
rect 5272 903 5306 929
rect 5272 861 5306 865
rect 5272 831 5306 861
rect 5272 759 5306 793
rect 5272 691 5306 721
rect 5272 687 5306 691
rect 5272 623 5306 649
rect 5272 615 5306 623
rect 5272 555 5306 577
rect 5272 543 5306 555
rect 5272 487 5306 505
rect 5272 471 5306 487
rect 5395 1839 5429 1873
rect 5395 1779 5429 1801
rect 5395 1767 5429 1779
rect 5395 1711 5429 1729
rect 5395 1695 5429 1711
rect 5395 1643 5429 1657
rect 5395 1623 5429 1643
rect 5395 1575 5429 1585
rect 5395 1551 5429 1575
rect 5395 1507 5429 1513
rect 5395 1479 5429 1507
rect 5395 1439 5429 1441
rect 5395 1407 5429 1439
rect 5395 1337 5429 1369
rect 5395 1335 5429 1337
rect 5395 1269 5429 1297
rect 5395 1263 5429 1269
rect 5395 1201 5429 1225
rect 5395 1191 5429 1201
rect 5395 1133 5429 1153
rect 5395 1119 5429 1133
rect 5395 1065 5429 1081
rect 5395 1047 5429 1065
rect 5395 997 5429 1009
rect 5395 975 5429 997
rect 5395 929 5429 937
rect 5395 903 5429 929
rect 5395 861 5429 865
rect 5395 831 5429 861
rect 5395 759 5429 793
rect 5395 691 5429 721
rect 5395 687 5429 691
rect 5395 623 5429 649
rect 5395 615 5429 623
rect 5395 555 5429 577
rect 5395 543 5429 555
rect 5395 487 5429 505
rect 5395 471 5429 487
rect 5558 1839 5592 1873
rect 5558 1779 5592 1801
rect 5558 1767 5592 1779
rect 5558 1711 5592 1729
rect 5558 1695 5592 1711
rect 5558 1643 5592 1657
rect 5558 1623 5592 1643
rect 5558 1575 5592 1585
rect 5558 1551 5592 1575
rect 5558 1507 5592 1513
rect 5558 1479 5592 1507
rect 5558 1439 5592 1441
rect 5558 1407 5592 1439
rect 5558 1337 5592 1369
rect 5558 1335 5592 1337
rect 5558 1269 5592 1297
rect 5558 1263 5592 1269
rect 5558 1201 5592 1225
rect 5558 1191 5592 1201
rect 5558 1133 5592 1153
rect 5558 1119 5592 1133
rect 5558 1065 5592 1081
rect 5558 1047 5592 1065
rect 5558 997 5592 1009
rect 5558 975 5592 997
rect 5558 929 5592 937
rect 5558 903 5592 929
rect 5558 861 5592 865
rect 5558 831 5592 861
rect 5558 759 5592 793
rect 5558 691 5592 721
rect 5558 687 5592 691
rect 5558 623 5592 649
rect 5558 615 5592 623
rect 5558 555 5592 577
rect 5558 543 5592 555
rect 5558 487 5592 505
rect 5558 471 5592 487
rect 5721 1839 5755 1873
rect 5721 1779 5755 1801
rect 5721 1767 5755 1779
rect 5721 1711 5755 1729
rect 5721 1695 5755 1711
rect 5721 1643 5755 1657
rect 5721 1623 5755 1643
rect 5721 1575 5755 1585
rect 5721 1551 5755 1575
rect 5721 1507 5755 1513
rect 5721 1479 5755 1507
rect 5721 1439 5755 1441
rect 5721 1407 5755 1439
rect 5721 1337 5755 1369
rect 5721 1335 5755 1337
rect 5721 1269 5755 1297
rect 5721 1263 5755 1269
rect 5721 1201 5755 1225
rect 5721 1191 5755 1201
rect 5721 1133 5755 1153
rect 5721 1119 5755 1133
rect 5721 1065 5755 1081
rect 5721 1047 5755 1065
rect 5721 997 5755 1009
rect 5721 975 5755 997
rect 5721 929 5755 937
rect 5721 903 5755 929
rect 5721 861 5755 865
rect 5721 831 5755 861
rect 5721 759 5755 793
rect 5721 691 5755 721
rect 5721 687 5755 691
rect 5721 623 5755 649
rect 5721 615 5755 623
rect 5721 555 5755 577
rect 5721 543 5755 555
rect 5721 487 5755 505
rect 5721 471 5755 487
rect 5884 1839 5918 1873
rect 5884 1779 5918 1801
rect 5884 1767 5918 1779
rect 5884 1711 5918 1729
rect 5884 1695 5918 1711
rect 5884 1643 5918 1657
rect 5884 1623 5918 1643
rect 5884 1575 5918 1585
rect 5884 1551 5918 1575
rect 5884 1507 5918 1513
rect 5884 1479 5918 1507
rect 5884 1439 5918 1441
rect 5884 1407 5918 1439
rect 5884 1337 5918 1369
rect 5884 1335 5918 1337
rect 5884 1269 5918 1297
rect 5884 1263 5918 1269
rect 5884 1201 5918 1225
rect 5884 1191 5918 1201
rect 5884 1133 5918 1153
rect 5884 1119 5918 1133
rect 5884 1065 5918 1081
rect 5884 1047 5918 1065
rect 5884 997 5918 1009
rect 5884 975 5918 997
rect 5884 929 5918 937
rect 5884 903 5918 929
rect 5884 861 5918 865
rect 5884 831 5918 861
rect 5884 759 5918 793
rect 5884 691 5918 721
rect 5884 687 5918 691
rect 5884 623 5918 649
rect 5884 615 5918 623
rect 5884 555 5918 577
rect 5884 543 5918 555
rect 5884 487 5918 505
rect 5884 471 5918 487
rect 6047 1839 6081 1873
rect 6047 1779 6081 1801
rect 6047 1767 6081 1779
rect 6047 1711 6081 1729
rect 6047 1695 6081 1711
rect 6047 1643 6081 1657
rect 6047 1623 6081 1643
rect 6047 1575 6081 1585
rect 6047 1551 6081 1575
rect 6047 1507 6081 1513
rect 6047 1479 6081 1507
rect 6047 1439 6081 1441
rect 6047 1407 6081 1439
rect 6047 1337 6081 1369
rect 6047 1335 6081 1337
rect 6047 1269 6081 1297
rect 6047 1263 6081 1269
rect 6047 1201 6081 1225
rect 6047 1191 6081 1201
rect 6047 1133 6081 1153
rect 6047 1119 6081 1133
rect 6047 1065 6081 1081
rect 6047 1047 6081 1065
rect 6047 997 6081 1009
rect 6047 975 6081 997
rect 6047 929 6081 937
rect 6047 903 6081 929
rect 6047 861 6081 865
rect 6047 831 6081 861
rect 6047 759 6081 793
rect 6047 691 6081 721
rect 6047 687 6081 691
rect 6047 623 6081 649
rect 6047 615 6081 623
rect 6047 555 6081 577
rect 6047 543 6081 555
rect 6047 487 6081 505
rect 6047 471 6081 487
rect 6210 1839 6244 1873
rect 6210 1779 6244 1801
rect 6210 1767 6244 1779
rect 6210 1711 6244 1729
rect 6210 1695 6244 1711
rect 6210 1643 6244 1657
rect 6210 1623 6244 1643
rect 6210 1575 6244 1585
rect 6210 1551 6244 1575
rect 6210 1507 6244 1513
rect 6210 1479 6244 1507
rect 6210 1439 6244 1441
rect 6210 1407 6244 1439
rect 6210 1337 6244 1369
rect 6210 1335 6244 1337
rect 6210 1269 6244 1297
rect 6210 1263 6244 1269
rect 6210 1201 6244 1225
rect 6210 1191 6244 1201
rect 6210 1133 6244 1153
rect 6210 1119 6244 1133
rect 6210 1065 6244 1081
rect 6210 1047 6244 1065
rect 6210 997 6244 1009
rect 6210 975 6244 997
rect 6210 929 6244 937
rect 6210 903 6244 929
rect 6210 861 6244 865
rect 6210 831 6244 861
rect 6210 759 6244 793
rect 6210 691 6244 721
rect 6210 687 6244 691
rect 6210 623 6244 649
rect 6210 615 6244 623
rect 6210 555 6244 577
rect 6210 543 6244 555
rect 6210 487 6244 505
rect 6210 471 6244 487
rect 6373 1839 6407 1873
rect 6373 1779 6407 1801
rect 6373 1767 6407 1779
rect 6373 1711 6407 1729
rect 6373 1695 6407 1711
rect 6373 1643 6407 1657
rect 6373 1623 6407 1643
rect 6373 1575 6407 1585
rect 6373 1551 6407 1575
rect 6373 1507 6407 1513
rect 6373 1479 6407 1507
rect 6373 1439 6407 1441
rect 6373 1407 6407 1439
rect 6373 1337 6407 1369
rect 6373 1335 6407 1337
rect 6373 1269 6407 1297
rect 6373 1263 6407 1269
rect 6373 1201 6407 1225
rect 6373 1191 6407 1201
rect 6373 1133 6407 1153
rect 6373 1119 6407 1133
rect 6373 1065 6407 1081
rect 6373 1047 6407 1065
rect 6373 997 6407 1009
rect 6373 975 6407 997
rect 6373 929 6407 937
rect 6373 903 6407 929
rect 6373 861 6407 865
rect 6373 831 6407 861
rect 6373 759 6407 793
rect 6373 691 6407 721
rect 6373 687 6407 691
rect 6373 623 6407 649
rect 6373 615 6407 623
rect 6373 555 6407 577
rect 6373 543 6407 555
rect 6373 487 6407 505
rect 6373 471 6407 487
rect 6536 1839 6570 1873
rect 6536 1779 6570 1801
rect 6536 1767 6570 1779
rect 6536 1711 6570 1729
rect 6536 1695 6570 1711
rect 6536 1643 6570 1657
rect 6536 1623 6570 1643
rect 6536 1575 6570 1585
rect 6536 1551 6570 1575
rect 6536 1507 6570 1513
rect 6536 1479 6570 1507
rect 6536 1439 6570 1441
rect 6536 1407 6570 1439
rect 6536 1337 6570 1369
rect 6536 1335 6570 1337
rect 6536 1269 6570 1297
rect 6536 1263 6570 1269
rect 6536 1201 6570 1225
rect 6536 1191 6570 1201
rect 6536 1133 6570 1153
rect 6536 1119 6570 1133
rect 6536 1065 6570 1081
rect 6536 1047 6570 1065
rect 6536 997 6570 1009
rect 6536 975 6570 997
rect 6536 929 6570 937
rect 6536 903 6570 929
rect 6536 861 6570 865
rect 6536 831 6570 861
rect 6536 759 6570 793
rect 6536 691 6570 721
rect 6536 687 6570 691
rect 6536 623 6570 649
rect 6536 615 6570 623
rect 6536 555 6570 577
rect 6536 543 6570 555
rect 6536 487 6570 505
rect 6536 471 6570 487
rect 6655 1829 6689 1851
rect 6655 1817 6689 1829
rect 6655 1761 6689 1776
rect 6655 1742 6689 1761
rect 6655 1693 6689 1701
rect 6655 1667 6689 1693
rect 6655 1625 6689 1626
rect 6655 1592 6689 1625
rect 6655 1523 6689 1551
rect 6655 1517 6689 1523
rect 6655 1455 6689 1477
rect 6655 1443 6689 1455
rect 6655 1387 6689 1403
rect 6655 1369 6689 1387
rect 6655 1319 6689 1329
rect 6655 1295 6689 1319
rect 6655 1251 6689 1255
rect 6655 1221 6689 1251
rect 6655 1149 6689 1181
rect 6655 1147 6689 1149
rect 6655 1081 6689 1107
rect 6655 1073 6689 1081
rect 6655 1013 6689 1033
rect 6655 999 6689 1013
rect 6655 945 6689 959
rect 6655 925 6689 945
rect 6655 877 6689 885
rect 6655 851 6689 877
rect 6655 809 6689 811
rect 6655 777 6689 809
rect 6655 707 6689 737
rect 6655 703 6689 707
rect 6655 639 6689 663
rect 6655 629 6689 639
rect 6655 571 6689 589
rect 6655 555 6689 571
rect 6655 503 6689 515
rect 6655 481 6689 503
rect 4005 405 4039 439
rect 6655 435 6689 441
rect 6655 407 6689 435
rect 4078 333 4107 367
rect 4107 333 4112 367
rect 4151 333 4175 367
rect 4175 333 4185 367
rect 4224 333 4243 367
rect 4243 333 4258 367
rect 4297 333 4311 367
rect 4311 333 4331 367
rect 4370 333 4379 367
rect 4379 333 4404 367
rect 4443 333 4447 367
rect 4447 333 4477 367
rect 4516 333 4549 367
rect 4549 333 4550 367
rect 4589 333 4617 367
rect 4617 333 4623 367
rect 4662 333 4685 367
rect 4685 333 4696 367
rect 4735 333 4753 367
rect 4753 333 4769 367
rect 4808 333 4821 367
rect 4821 333 4842 367
rect 4881 333 4889 367
rect 4889 333 4915 367
rect 4955 333 4957 367
rect 4957 333 4989 367
rect 5029 333 5059 367
rect 5059 333 5063 367
rect 5103 333 5127 367
rect 5127 333 5137 367
rect 5177 333 5195 367
rect 5195 333 5211 367
rect 5251 333 5263 367
rect 5263 333 5285 367
rect 5325 333 5331 367
rect 5331 333 5359 367
rect 5399 333 5433 367
rect 5473 333 5501 367
rect 5501 333 5507 367
rect 5547 333 5569 367
rect 5569 333 5581 367
rect 5621 333 5637 367
rect 5637 333 5655 367
rect 5695 333 5705 367
rect 5705 333 5729 367
rect 5769 333 5773 367
rect 5773 333 5803 367
rect 5843 333 5875 367
rect 5875 333 5877 367
rect 5917 333 5943 367
rect 5943 333 5951 367
rect 5991 333 6011 367
rect 6011 333 6025 367
rect 6065 333 6079 367
rect 6079 333 6099 367
rect 6139 333 6147 367
rect 6147 333 6173 367
rect 6213 333 6215 367
rect 6215 333 6247 367
rect 6287 333 6317 367
rect 6317 333 6321 367
rect 6361 333 6385 367
rect 6385 333 6395 367
rect 6435 333 6453 367
rect 6453 333 6469 367
rect 6509 333 6521 367
rect 6521 333 6543 367
rect 6583 333 6617 367
rect 6876 2028 6910 2062
rect 6876 1954 6910 1988
rect 6876 1880 6910 1914
rect 6876 1806 6910 1840
rect 6876 1732 6910 1766
rect 6876 1658 6910 1692
rect 6876 1584 6910 1618
rect 6876 1510 6910 1544
rect 6876 1437 6910 1471
rect 6876 1364 6910 1398
rect 6876 1291 6910 1325
rect 6876 1218 6910 1252
rect 6876 1145 6910 1179
rect 6876 1072 6910 1106
rect 6876 999 6910 1033
rect 6876 926 6910 960
rect 6876 853 6910 887
rect 6876 780 6910 814
rect 6876 707 6910 741
rect 6876 634 6910 668
rect 6876 561 6910 595
rect 6876 488 6910 522
rect 6876 415 6910 449
rect 7170 2073 7175 2107
rect 7175 2073 7204 2107
rect 7243 2073 7277 2107
rect 7316 2073 7345 2107
rect 7345 2073 7350 2107
rect 7389 2073 7413 2107
rect 7413 2073 7423 2107
rect 7463 2073 7481 2107
rect 7481 2073 7497 2107
rect 7537 2073 7549 2107
rect 7549 2073 7571 2107
rect 7611 2073 7617 2107
rect 7617 2073 7645 2107
rect 7685 2073 7719 2107
rect 7759 2073 7787 2107
rect 7787 2073 7793 2107
rect 7833 2073 7855 2107
rect 7855 2073 7867 2107
rect 7907 2073 7923 2107
rect 7923 2073 7941 2107
rect 7981 2073 7991 2107
rect 7991 2073 8015 2107
rect 8055 2073 8059 2107
rect 8059 2073 8089 2107
rect 8129 2073 8161 2107
rect 8161 2073 8163 2107
rect 8203 2073 8229 2107
rect 8229 2073 8237 2107
rect 8277 2073 8297 2107
rect 8297 2073 8311 2107
rect 8351 2073 8365 2107
rect 8365 2073 8385 2107
rect 8425 2073 8433 2107
rect 8433 2073 8459 2107
rect 8499 2073 8501 2107
rect 8501 2073 8533 2107
rect 8573 2073 8603 2107
rect 8603 2073 8607 2107
rect 8647 2073 8671 2107
rect 8671 2073 8681 2107
rect 8721 2073 8739 2107
rect 8739 2073 8755 2107
rect 8795 2073 8807 2107
rect 8807 2073 8829 2107
rect 8869 2073 8875 2107
rect 8875 2073 8903 2107
rect 8943 2073 8977 2107
rect 9017 2073 9045 2107
rect 9045 2073 9051 2107
rect 9091 2073 9113 2107
rect 9113 2073 9125 2107
rect 9165 2073 9181 2107
rect 9181 2073 9199 2107
rect 9239 2073 9249 2107
rect 9249 2073 9273 2107
rect 9313 2073 9317 2107
rect 9317 2073 9347 2107
rect 9387 2073 9419 2107
rect 9419 2073 9421 2107
rect 9461 2073 9487 2107
rect 9487 2073 9495 2107
rect 9535 2073 9555 2107
rect 9555 2073 9569 2107
rect 9645 2073 9657 2107
rect 9657 2073 9679 2107
rect 9727 2073 9759 2107
rect 9759 2073 9761 2107
rect 9809 2073 9827 2107
rect 9827 2073 9843 2107
rect 9891 2073 9895 2107
rect 9895 2073 9925 2107
rect 7097 2005 7131 2035
rect 7097 2001 7131 2005
rect 7273 1991 7277 2025
rect 7277 1991 7307 2025
rect 7346 1991 7350 2025
rect 7350 1991 7380 2025
rect 7419 1991 7423 2025
rect 7423 1991 7453 2025
rect 7492 1991 7496 2025
rect 7496 1991 7526 2025
rect 7565 1991 7569 2025
rect 7569 1991 7599 2025
rect 7638 1991 7641 2025
rect 7641 1991 7672 2025
rect 7711 1991 7713 2025
rect 7713 1991 7745 2025
rect 7784 1991 7785 2025
rect 7785 1991 7818 2025
rect 7857 1991 7891 2025
rect 7930 1991 7963 2025
rect 7963 1991 7964 2025
rect 8003 1991 8035 2025
rect 8035 1991 8037 2025
rect 8075 1991 8107 2025
rect 8107 1991 8109 2025
rect 8147 1991 8179 2025
rect 8179 1991 8181 2025
rect 8544 1991 8548 2025
rect 8548 1991 8578 2025
rect 8619 1991 8651 2025
rect 8651 1991 8653 2025
rect 8694 1991 8720 2025
rect 8720 1991 8728 2025
rect 8769 1991 8789 2025
rect 8789 1991 8803 2025
rect 8844 1991 8858 2025
rect 8858 1991 8878 2025
rect 8918 1991 8927 2025
rect 8927 1991 8952 2025
rect 8992 1991 8996 2025
rect 8996 1991 9026 2025
rect 9066 1991 9100 2025
rect 9140 1991 9169 2025
rect 9169 1991 9174 2025
rect 9214 1991 9238 2025
rect 9238 1991 9248 2025
rect 9288 1991 9307 2025
rect 9307 1991 9322 2025
rect 9362 1991 9376 2025
rect 9376 1991 9396 2025
rect 9436 1991 9444 2025
rect 9444 1991 9470 2025
rect 9510 1991 9512 2025
rect 9512 1991 9544 2025
rect 9584 1991 9614 2025
rect 9614 1991 9618 2025
rect 9658 1991 9682 2025
rect 9682 1991 9692 2025
rect 9732 1991 9750 2025
rect 9750 1991 9766 2025
rect 9963 1999 9997 2033
rect 7097 1937 7131 1960
rect 7097 1926 7131 1937
rect 7097 1869 7131 1885
rect 7097 1851 7131 1869
rect 7097 1801 7131 1810
rect 7097 1776 7131 1801
rect 7097 1733 7131 1735
rect 7097 1701 7131 1733
rect 7097 1631 7131 1660
rect 7097 1626 7131 1631
rect 7097 1563 7131 1585
rect 7097 1551 7131 1563
rect 7097 1495 7131 1510
rect 7097 1476 7131 1495
rect 7097 1427 7131 1435
rect 7097 1401 7131 1427
rect 7097 1359 7131 1360
rect 7097 1326 7131 1359
rect 7097 1257 7131 1285
rect 7097 1251 7131 1257
rect 7097 1189 7131 1210
rect 7097 1176 7131 1189
rect 7097 1121 7131 1135
rect 7097 1101 7131 1121
rect 7097 1053 7131 1061
rect 7097 1027 7131 1053
rect 7097 985 7131 987
rect 7097 953 7131 985
rect 7097 883 7131 913
rect 7097 879 7131 883
rect 7097 815 7131 839
rect 7097 805 7131 815
rect 7097 747 7131 765
rect 7097 731 7131 747
rect 7097 679 7131 691
rect 7097 657 7131 679
rect 7097 583 7131 617
rect 7097 520 7131 543
rect 7097 509 7131 520
rect 7216 1907 7250 1941
rect 7216 1847 7250 1869
rect 7216 1835 7250 1847
rect 7216 1779 7250 1797
rect 7216 1763 7250 1779
rect 7216 1711 7250 1725
rect 7216 1691 7250 1711
rect 7216 1643 7250 1653
rect 7216 1619 7250 1643
rect 7216 1575 7250 1581
rect 7216 1547 7250 1575
rect 7216 1507 7250 1509
rect 7216 1475 7250 1507
rect 7216 1405 7250 1437
rect 7216 1403 7250 1405
rect 7216 1337 7250 1365
rect 7216 1331 7250 1337
rect 7216 1269 7250 1293
rect 7216 1259 7250 1269
rect 7216 1201 7250 1221
rect 7216 1187 7250 1201
rect 7216 1133 7250 1149
rect 7216 1115 7250 1133
rect 7216 1065 7250 1077
rect 7216 1043 7250 1065
rect 7216 997 7250 1005
rect 7216 971 7250 997
rect 7216 929 7250 933
rect 7216 899 7250 929
rect 7216 827 7250 861
rect 7216 759 7250 789
rect 7216 755 7250 759
rect 7216 691 7250 717
rect 7216 683 7250 691
rect 7216 623 7250 645
rect 7216 611 7250 623
rect 7216 555 7250 573
rect 7216 539 7250 555
rect 7379 1907 7413 1941
rect 7379 1847 7413 1869
rect 7379 1835 7413 1847
rect 7379 1779 7413 1797
rect 7379 1763 7413 1779
rect 7379 1711 7413 1725
rect 7379 1691 7413 1711
rect 7379 1643 7413 1653
rect 7379 1619 7413 1643
rect 7379 1575 7413 1581
rect 7379 1547 7413 1575
rect 7379 1507 7413 1509
rect 7379 1475 7413 1507
rect 7379 1405 7413 1437
rect 7379 1403 7413 1405
rect 7379 1337 7413 1365
rect 7379 1331 7413 1337
rect 7379 1269 7413 1293
rect 7379 1259 7413 1269
rect 7379 1201 7413 1221
rect 7379 1187 7413 1201
rect 7379 1133 7413 1149
rect 7379 1115 7413 1133
rect 7379 1065 7413 1077
rect 7379 1043 7413 1065
rect 7379 997 7413 1005
rect 7379 971 7413 997
rect 7379 929 7413 933
rect 7379 899 7413 929
rect 7379 827 7413 861
rect 7379 759 7413 789
rect 7379 755 7413 759
rect 7379 691 7413 717
rect 7379 683 7413 691
rect 7379 623 7413 645
rect 7379 611 7413 623
rect 7379 555 7413 573
rect 7379 539 7413 555
rect 7542 1907 7576 1941
rect 7542 1847 7576 1869
rect 7542 1835 7576 1847
rect 7542 1779 7576 1797
rect 7542 1763 7576 1779
rect 7542 1711 7576 1725
rect 7542 1691 7576 1711
rect 7542 1643 7576 1653
rect 7542 1619 7576 1643
rect 7542 1575 7576 1581
rect 7542 1547 7576 1575
rect 7542 1507 7576 1509
rect 7542 1475 7576 1507
rect 7542 1405 7576 1437
rect 7542 1403 7576 1405
rect 7542 1337 7576 1365
rect 7542 1331 7576 1337
rect 7542 1269 7576 1293
rect 7542 1259 7576 1269
rect 7542 1201 7576 1221
rect 7542 1187 7576 1201
rect 7542 1133 7576 1149
rect 7542 1115 7576 1133
rect 7542 1065 7576 1077
rect 7542 1043 7576 1065
rect 7542 997 7576 1005
rect 7542 971 7576 997
rect 7542 929 7576 933
rect 7542 899 7576 929
rect 7542 827 7576 861
rect 7542 759 7576 789
rect 7542 755 7576 759
rect 7542 691 7576 717
rect 7542 683 7576 691
rect 7542 623 7576 645
rect 7542 611 7576 623
rect 7542 555 7576 573
rect 7542 539 7576 555
rect 7705 1907 7739 1941
rect 7705 1847 7739 1869
rect 7705 1835 7739 1847
rect 7705 1779 7739 1797
rect 7705 1763 7739 1779
rect 7705 1711 7739 1725
rect 7705 1691 7739 1711
rect 7705 1643 7739 1653
rect 7705 1619 7739 1643
rect 7705 1575 7739 1581
rect 7705 1547 7739 1575
rect 7705 1507 7739 1509
rect 7705 1475 7739 1507
rect 7705 1405 7739 1437
rect 7705 1403 7739 1405
rect 7705 1337 7739 1365
rect 7705 1331 7739 1337
rect 7705 1269 7739 1293
rect 7705 1259 7739 1269
rect 7705 1201 7739 1221
rect 7705 1187 7739 1201
rect 7705 1133 7739 1149
rect 7705 1115 7739 1133
rect 7705 1065 7739 1077
rect 7705 1043 7739 1065
rect 7705 997 7739 1005
rect 7705 971 7739 997
rect 7705 929 7739 933
rect 7705 899 7739 929
rect 7705 827 7739 861
rect 7705 759 7739 789
rect 7705 755 7739 759
rect 7705 691 7739 717
rect 7705 683 7739 691
rect 7705 623 7739 645
rect 7705 611 7739 623
rect 7705 555 7739 573
rect 7705 539 7739 555
rect 7868 1907 7902 1941
rect 7868 1847 7902 1869
rect 7868 1835 7902 1847
rect 7868 1779 7902 1797
rect 7868 1763 7902 1779
rect 7868 1711 7902 1725
rect 7868 1691 7902 1711
rect 7868 1643 7902 1653
rect 7868 1619 7902 1643
rect 7868 1575 7902 1581
rect 7868 1547 7902 1575
rect 7868 1507 7902 1509
rect 7868 1475 7902 1507
rect 7868 1405 7902 1437
rect 7868 1403 7902 1405
rect 7868 1337 7902 1365
rect 7868 1331 7902 1337
rect 7868 1269 7902 1293
rect 7868 1259 7902 1269
rect 7868 1201 7902 1221
rect 7868 1187 7902 1201
rect 7868 1133 7902 1149
rect 7868 1115 7902 1133
rect 7868 1065 7902 1077
rect 7868 1043 7902 1065
rect 7868 997 7902 1005
rect 7868 971 7902 997
rect 7868 929 7902 933
rect 7868 899 7902 929
rect 7868 827 7902 861
rect 7868 759 7902 789
rect 7868 755 7902 759
rect 7868 691 7902 717
rect 7868 683 7902 691
rect 7868 623 7902 645
rect 7868 611 7902 623
rect 7868 555 7902 573
rect 7868 539 7902 555
rect 8031 1907 8065 1941
rect 8031 1847 8065 1869
rect 8031 1835 8065 1847
rect 8031 1779 8065 1797
rect 8031 1763 8065 1779
rect 8031 1711 8065 1725
rect 8031 1691 8065 1711
rect 8031 1643 8065 1653
rect 8031 1619 8065 1643
rect 8031 1575 8065 1581
rect 8031 1547 8065 1575
rect 8031 1507 8065 1509
rect 8031 1475 8065 1507
rect 8031 1405 8065 1437
rect 8031 1403 8065 1405
rect 8031 1337 8065 1365
rect 8031 1331 8065 1337
rect 8031 1269 8065 1293
rect 8031 1259 8065 1269
rect 8031 1201 8065 1221
rect 8031 1187 8065 1201
rect 8031 1133 8065 1149
rect 8031 1115 8065 1133
rect 8031 1065 8065 1077
rect 8031 1043 8065 1065
rect 8031 997 8065 1005
rect 8031 971 8065 997
rect 8031 929 8065 933
rect 8031 899 8065 929
rect 8031 827 8065 861
rect 8031 759 8065 789
rect 8031 755 8065 759
rect 8031 691 8065 717
rect 8031 683 8065 691
rect 8031 623 8065 645
rect 8031 611 8065 623
rect 8031 555 8065 573
rect 8031 539 8065 555
rect 8194 1907 8228 1941
rect 8194 1847 8228 1869
rect 8194 1835 8228 1847
rect 8194 1779 8228 1797
rect 8194 1763 8228 1779
rect 8194 1711 8228 1725
rect 8194 1691 8228 1711
rect 8194 1643 8228 1653
rect 8194 1619 8228 1643
rect 8194 1575 8228 1581
rect 8194 1547 8228 1575
rect 8194 1507 8228 1509
rect 8194 1475 8228 1507
rect 8194 1405 8228 1437
rect 8194 1403 8228 1405
rect 8194 1337 8228 1365
rect 8194 1331 8228 1337
rect 8194 1269 8228 1293
rect 8194 1259 8228 1269
rect 8194 1201 8228 1221
rect 8194 1187 8228 1201
rect 8194 1133 8228 1149
rect 8194 1115 8228 1133
rect 8194 1065 8228 1077
rect 8194 1043 8228 1065
rect 8194 997 8228 1005
rect 8194 971 8228 997
rect 8194 929 8228 933
rect 8194 899 8228 929
rect 8194 827 8228 861
rect 8194 759 8228 789
rect 8194 755 8228 759
rect 8194 691 8228 717
rect 8194 683 8228 691
rect 8194 623 8228 645
rect 8194 611 8228 623
rect 8194 555 8228 573
rect 8194 539 8228 555
rect 8357 1907 8391 1941
rect 9963 1931 9997 1959
rect 9963 1925 9997 1931
rect 8357 1847 8391 1869
rect 8357 1835 8391 1847
rect 8357 1779 8391 1797
rect 8357 1763 8391 1779
rect 8357 1711 8391 1725
rect 8357 1691 8391 1711
rect 8357 1643 8391 1653
rect 8357 1619 8391 1643
rect 8357 1575 8391 1581
rect 8357 1547 8391 1575
rect 8357 1507 8391 1509
rect 8357 1475 8391 1507
rect 8357 1405 8391 1437
rect 8357 1403 8391 1405
rect 8357 1337 8391 1365
rect 8357 1331 8391 1337
rect 8357 1269 8391 1293
rect 8357 1259 8391 1269
rect 8357 1201 8391 1221
rect 8357 1187 8391 1201
rect 8357 1133 8391 1149
rect 8357 1115 8391 1133
rect 8357 1065 8391 1077
rect 8357 1043 8391 1065
rect 8357 997 8391 1005
rect 8357 971 8391 997
rect 8357 929 8391 933
rect 8357 899 8391 929
rect 8357 827 8391 861
rect 8357 759 8391 789
rect 8357 755 8391 759
rect 8357 691 8391 717
rect 8357 683 8391 691
rect 8357 623 8391 645
rect 8357 611 8391 623
rect 8357 555 8391 573
rect 8357 539 8391 555
rect 8480 1881 8514 1899
rect 8480 1865 8514 1881
rect 8480 1813 8514 1824
rect 8480 1790 8514 1813
rect 8480 1745 8514 1749
rect 8480 1715 8514 1745
rect 8480 1643 8514 1674
rect 8480 1640 8514 1643
rect 8480 1575 8514 1599
rect 8480 1565 8514 1575
rect 8480 1507 8514 1524
rect 8480 1490 8514 1507
rect 8480 1439 8514 1449
rect 8480 1415 8514 1439
rect 8480 1371 8514 1374
rect 8480 1340 8514 1371
rect 8480 1269 8514 1299
rect 8480 1265 8514 1269
rect 8480 1201 8514 1224
rect 8480 1190 8514 1201
rect 8480 1133 8514 1149
rect 8480 1115 8514 1133
rect 8480 1065 8514 1073
rect 8480 1039 8514 1065
rect 8480 963 8514 997
rect 8480 895 8514 921
rect 8480 887 8514 895
rect 8480 827 8514 845
rect 8480 811 8514 827
rect 8480 759 8514 769
rect 8480 735 8514 759
rect 8480 691 8514 693
rect 8480 659 8514 691
rect 8480 589 8514 617
rect 8480 583 8514 589
rect 8480 507 8514 541
rect 8643 1881 8677 1897
rect 8643 1863 8677 1881
rect 8643 1813 8677 1824
rect 8643 1790 8677 1813
rect 8643 1745 8677 1751
rect 8643 1717 8677 1745
rect 8643 1677 8677 1678
rect 8643 1644 8677 1677
rect 8643 1575 8677 1605
rect 8643 1571 8677 1575
rect 8643 1507 8677 1531
rect 8643 1497 8677 1507
rect 8643 1439 8677 1457
rect 8643 1423 8677 1439
rect 8643 1371 8677 1383
rect 8643 1349 8677 1371
rect 8806 1065 8840 1087
rect 8806 1053 8840 1065
rect 8806 997 8840 1009
rect 8806 975 8840 997
rect 8806 929 8840 931
rect 8806 897 8840 929
rect 8806 827 8840 853
rect 8806 819 8840 827
rect 8806 759 8840 775
rect 8806 741 8840 759
rect 8806 691 8840 697
rect 8806 663 8840 691
rect 8806 589 8840 619
rect 8806 585 8840 589
rect 8806 507 8840 541
rect 8969 1881 9003 1897
rect 8969 1863 9003 1881
rect 8969 1813 9003 1824
rect 8969 1790 9003 1813
rect 8969 1745 9003 1751
rect 8969 1717 9003 1745
rect 8969 1677 9003 1678
rect 8969 1644 9003 1677
rect 8969 1575 9003 1605
rect 8969 1571 9003 1575
rect 8969 1507 9003 1531
rect 8969 1497 9003 1507
rect 8969 1439 9003 1457
rect 8969 1423 9003 1439
rect 8969 1371 9003 1383
rect 8969 1349 9003 1371
rect 9132 1065 9166 1087
rect 9132 1053 9166 1065
rect 9132 997 9166 1009
rect 9132 975 9166 997
rect 9132 929 9166 931
rect 9132 897 9166 929
rect 9132 827 9166 853
rect 9132 819 9166 827
rect 9132 759 9166 775
rect 9132 741 9166 759
rect 9132 691 9166 697
rect 9132 663 9166 691
rect 9132 589 9166 619
rect 9132 585 9166 589
rect 9132 507 9166 541
rect 9295 1881 9329 1897
rect 9295 1863 9329 1881
rect 9295 1813 9329 1824
rect 9295 1790 9329 1813
rect 9295 1745 9329 1751
rect 9295 1717 9329 1745
rect 9295 1677 9329 1678
rect 9295 1644 9329 1677
rect 9295 1575 9329 1605
rect 9295 1571 9329 1575
rect 9295 1507 9329 1531
rect 9295 1497 9329 1507
rect 9295 1439 9329 1457
rect 9295 1423 9329 1439
rect 9295 1371 9329 1383
rect 9295 1349 9329 1371
rect 9458 1065 9492 1087
rect 9458 1053 9492 1065
rect 9458 997 9492 1009
rect 9458 975 9492 997
rect 9458 929 9492 931
rect 9458 897 9492 929
rect 9458 827 9492 853
rect 9458 819 9492 827
rect 9458 759 9492 775
rect 9458 741 9492 759
rect 9458 691 9492 697
rect 9458 663 9492 691
rect 9458 589 9492 619
rect 9458 585 9492 589
rect 9458 507 9492 541
rect 9621 1881 9655 1897
rect 9621 1863 9655 1881
rect 9621 1813 9655 1824
rect 9621 1790 9655 1813
rect 9621 1745 9655 1751
rect 9621 1717 9655 1745
rect 9621 1677 9655 1678
rect 9621 1644 9655 1677
rect 9621 1575 9655 1605
rect 9621 1571 9655 1575
rect 9621 1507 9655 1531
rect 9621 1497 9655 1507
rect 9621 1439 9655 1457
rect 9621 1423 9655 1439
rect 9621 1371 9655 1383
rect 9621 1349 9655 1371
rect 9784 1065 9818 1087
rect 9784 1053 9818 1065
rect 9784 997 9818 1009
rect 9784 975 9818 997
rect 9784 929 9818 931
rect 9784 897 9818 929
rect 9784 827 9818 853
rect 9784 819 9818 827
rect 9784 759 9818 775
rect 9784 741 9818 759
rect 9784 691 9818 697
rect 9784 663 9818 691
rect 9784 589 9818 619
rect 9784 585 9818 589
rect 9784 507 9818 541
rect 9963 1863 9997 1885
rect 9963 1851 9997 1863
rect 9963 1795 9997 1811
rect 9963 1777 9997 1795
rect 9963 1727 9997 1737
rect 9963 1703 9997 1727
rect 9963 1659 9997 1663
rect 9963 1629 9997 1659
rect 9963 1557 9997 1589
rect 9963 1555 9997 1557
rect 9963 1489 9997 1515
rect 9963 1481 9997 1489
rect 9963 1421 9997 1441
rect 9963 1407 9997 1421
rect 9963 1353 9997 1366
rect 9963 1332 9997 1353
rect 9963 1285 9997 1291
rect 9963 1257 9997 1285
rect 9963 1183 9997 1216
rect 9963 1182 9997 1183
rect 9963 1115 9997 1141
rect 9963 1107 9997 1115
rect 9963 1047 9997 1066
rect 9963 1032 9997 1047
rect 9963 979 9997 991
rect 9963 957 9997 979
rect 9963 911 9997 916
rect 9963 882 9997 911
rect 9963 809 9997 841
rect 9963 807 9997 809
rect 9963 741 9997 766
rect 9963 732 9997 741
rect 9963 673 9997 691
rect 9963 657 9997 673
rect 9963 605 9997 616
rect 9963 582 9997 605
rect 9963 537 9997 541
rect 9963 507 9997 537
rect 7169 447 7199 469
rect 7169 435 7199 447
rect 7199 435 7203 469
rect 7243 447 7267 469
rect 7243 435 7267 447
rect 7267 435 7277 469
rect 7317 447 7335 469
rect 7317 435 7335 447
rect 7335 435 7351 469
rect 7391 447 7403 469
rect 7391 435 7403 447
rect 7403 435 7425 469
rect 7465 447 7471 469
rect 7465 435 7471 447
rect 7471 435 7499 469
rect 7539 435 7573 469
rect 7613 435 7641 469
rect 7641 447 7647 469
rect 7641 435 7647 447
rect 7687 435 7709 469
rect 7709 447 7721 469
rect 7709 435 7721 447
rect 7761 435 7777 469
rect 7777 447 7795 469
rect 7777 435 7795 447
rect 7835 435 7845 469
rect 7845 447 7869 469
rect 7845 435 7869 447
rect 7909 435 7913 469
rect 7913 447 7943 469
rect 7913 435 7943 447
rect 7983 447 8015 469
rect 7983 435 8015 447
rect 8015 435 8017 469
rect 8057 447 8083 469
rect 8057 435 8083 447
rect 8083 435 8091 469
rect 8131 447 8151 469
rect 8131 435 8151 447
rect 8151 435 8165 469
rect 8205 447 8219 469
rect 8205 435 8219 447
rect 8219 435 8239 469
rect 8279 447 8287 469
rect 8279 435 8287 447
rect 8287 435 8313 469
rect 8353 447 8355 469
rect 8353 435 8355 447
rect 8355 435 8387 469
rect 8427 435 8457 469
rect 8457 447 8461 469
rect 8457 435 8461 447
rect 8501 435 8525 469
rect 8525 447 8535 469
rect 8525 435 8535 447
rect 8575 435 8593 469
rect 8593 447 8609 469
rect 8593 435 8609 447
rect 8649 435 8661 469
rect 8661 447 8683 469
rect 8661 435 8683 447
rect 8722 435 8729 469
rect 8729 447 8756 469
rect 8729 435 8756 447
rect 8795 435 8797 469
rect 8797 447 8829 469
rect 8797 435 8829 447
rect 8868 447 8899 469
rect 8868 435 8899 447
rect 8899 435 8902 469
rect 8941 447 8967 469
rect 8941 435 8967 447
rect 8967 435 8975 469
rect 9014 447 9035 469
rect 9014 435 9035 447
rect 9035 435 9048 469
rect 9087 447 9103 469
rect 9087 435 9103 447
rect 9103 435 9121 469
rect 9160 447 9171 469
rect 9160 435 9171 447
rect 9171 435 9194 469
rect 9233 447 9239 469
rect 9233 435 9239 447
rect 9239 435 9267 469
rect 9306 447 9307 469
rect 9306 435 9307 447
rect 9307 435 9340 469
rect 9379 435 9409 469
rect 9409 447 9413 469
rect 9409 435 9413 447
rect 9452 435 9477 469
rect 9477 447 9486 469
rect 9477 435 9486 447
rect 9525 435 9545 469
rect 9545 447 9559 469
rect 9545 435 9559 447
rect 9598 435 9613 469
rect 9613 447 9632 469
rect 9613 435 9632 447
rect 9671 435 9681 469
rect 9681 447 9705 469
rect 9681 435 9705 447
rect 9744 435 9749 469
rect 9749 447 9778 469
rect 9749 435 9778 447
rect 9817 447 9851 469
rect 9817 435 9851 447
rect 9890 447 9919 469
rect 9890 435 9919 447
rect 9919 435 9924 469
rect 10189 2106 10223 2140
rect 10189 2034 10223 2068
rect 10189 1962 10223 1996
rect 10189 1890 10223 1924
rect 10189 1818 10223 1852
rect 10189 1746 10223 1780
rect 10189 1674 10223 1708
rect 10189 1602 10223 1636
rect 10189 1530 10223 1564
rect 10189 1458 10223 1492
rect 10189 1386 10223 1420
rect 10189 1314 10223 1348
rect 10189 1242 10223 1276
rect 10189 1170 10223 1204
rect 10189 1098 10223 1132
rect 10189 1026 10223 1060
rect 10189 954 10223 988
rect 10189 881 10223 915
rect 10189 808 10223 842
rect 10189 735 10223 769
rect 10189 662 10223 696
rect 10189 589 10223 623
rect 10189 516 10223 550
rect 10189 472 10223 477
rect 10189 443 10223 472
rect 6876 342 6910 376
rect 3784 270 3818 304
rect 3784 196 3818 230
rect 3784 122 3818 156
rect 6876 269 6910 303
rect 10189 370 10223 404
rect 10189 297 10223 331
rect 10189 248 10223 258
rect 6876 196 6910 230
rect 10189 224 10194 248
rect 10194 224 10223 248
rect 6956 180 6990 214
rect 7029 180 7032 214
rect 7032 180 7063 214
rect 7102 180 7136 214
rect 7175 180 7209 214
rect 7248 180 7282 214
rect 7321 180 7355 214
rect 7394 180 7428 214
rect 7467 180 7501 214
rect 7540 180 7574 214
rect 7613 180 7647 214
rect 7686 180 7720 214
rect 7759 180 7793 214
rect 7832 180 7866 214
rect 7905 180 7939 214
rect 7978 180 8012 214
rect 8051 180 8085 214
rect 8124 180 8158 214
rect 8197 180 8231 214
rect 8270 180 8304 214
rect 8343 180 8377 214
rect 8416 180 8450 214
rect 8489 180 8523 214
rect 8561 180 8595 214
rect 8633 180 8667 214
rect 8705 180 8739 214
rect 8777 180 8811 214
rect 8849 180 8883 214
rect 8921 180 8955 214
rect 8993 180 9027 214
rect 9065 180 9099 214
rect 9137 180 9171 214
rect 9209 180 9243 214
rect 9281 180 9315 214
rect 9353 180 9387 214
rect 9425 180 9459 214
rect 9497 180 9531 214
rect 9569 180 9603 214
rect 9641 180 9675 214
rect 9713 180 9747 214
rect 9785 180 9819 214
rect 9857 180 9891 214
rect 9929 180 9963 214
rect 10001 180 10035 214
rect 10073 180 10107 214
rect 3902 78 3918 112
rect 3918 78 3936 112
rect 3975 78 4009 112
rect 4048 78 4082 112
rect 4121 78 4155 112
rect 4194 78 4228 112
rect 4267 78 4301 112
rect 4340 78 4374 112
rect 4413 78 4447 112
rect 4486 78 4520 112
rect 4559 78 4593 112
rect 4632 78 4666 112
rect 4705 78 4739 112
rect 4778 78 4812 112
rect 4851 78 4885 112
rect 4924 78 4958 112
rect 4997 78 5031 112
rect 5070 78 5104 112
rect 5143 78 5177 112
rect 5216 78 5250 112
rect 5289 78 5323 112
rect 5362 78 5396 112
rect 5435 78 5469 112
rect 5508 78 5542 112
rect 5581 78 5615 112
rect 5654 78 5688 112
rect 5727 78 5761 112
rect 5800 78 5834 112
rect 5873 78 5907 112
rect 5946 78 5980 112
rect 6019 78 6053 112
rect 6092 78 6126 112
rect 6166 78 6200 112
rect 6240 78 6274 112
rect 6314 78 6348 112
rect 6388 78 6422 112
rect 6462 78 6496 112
rect 6536 78 6570 112
rect 6610 78 6644 112
rect 6684 78 6718 112
rect 6758 78 6792 112
rect 6832 78 6866 112
<< metal1 >>
rect -24 2328 3537 2362
rect -24 2294 54 2328
rect 88 2294 148 2328
rect 182 2294 241 2328
rect 275 2294 334 2328
rect 368 2294 410 2328
rect 444 2294 484 2328
rect 518 2294 558 2328
rect 592 2294 632 2328
rect 666 2294 706 2328
rect 740 2294 780 2328
rect 814 2294 854 2328
rect 888 2294 928 2328
rect 962 2294 1002 2328
rect 1036 2294 1076 2328
rect 1110 2294 1150 2328
rect 1184 2294 1224 2328
rect 1258 2294 1298 2328
rect 1332 2294 1372 2328
rect 1406 2294 1446 2328
rect 1480 2294 1520 2328
rect 1554 2294 1594 2328
rect 1628 2294 1668 2328
rect 1702 2294 1742 2328
rect 1776 2294 1816 2328
rect 1850 2294 1890 2328
rect 1924 2294 1964 2328
rect 1998 2294 2037 2328
rect 2071 2294 2110 2328
rect 2144 2294 2183 2328
rect 2217 2294 2256 2328
rect 2290 2294 2329 2328
rect 2363 2294 2402 2328
rect 2436 2294 2475 2328
rect 2509 2294 2548 2328
rect 2582 2294 2621 2328
rect 2655 2294 2694 2328
rect 2728 2294 2767 2328
rect 2801 2294 2840 2328
rect 2874 2294 2913 2328
rect 2947 2294 2986 2328
rect 3020 2294 3059 2328
rect 3093 2294 3132 2328
rect 3166 2294 3205 2328
rect 3239 2294 3278 2328
rect 3312 2294 3351 2328
rect 3385 2294 3537 2328
rect -24 2284 3537 2294
rect -24 2260 3469 2284
rect -24 2250 102 2260
tri 102 2250 112 2260 nw
tri 1550 2250 1560 2260 ne
rect 1560 2250 1994 2260
tri 1994 2250 2004 2260 nw
tri 3401 2250 3411 2260 ne
rect 3411 2250 3469 2260
rect 3503 2250 3537 2284
rect -24 2228 80 2250
tri 80 2228 102 2250 nw
tri 1560 2228 1582 2250 ne
rect 1582 2228 1956 2250
rect -24 2210 78 2228
tri 78 2226 80 2228 nw
tri 1582 2226 1584 2228 ne
rect 1584 2226 1648 2228
rect -24 2176 10 2210
rect 44 2176 78 2210
rect -24 2137 78 2176
tri 1584 2169 1641 2226 ne
rect -24 2103 10 2137
rect 44 2103 78 2137
rect -24 2064 78 2103
rect -24 2030 10 2064
rect 44 2030 78 2064
rect -24 1991 78 2030
rect -24 1957 10 1991
rect 44 1957 78 1991
rect -24 1918 78 1957
rect -24 1884 10 1918
rect 44 1884 78 1918
rect -24 1845 78 1884
rect -24 1811 10 1845
rect 44 1811 78 1845
rect -24 1772 78 1811
rect -24 1738 10 1772
rect 44 1738 78 1772
rect -24 1699 78 1738
rect -24 1665 10 1699
rect 44 1665 78 1699
rect -24 1626 78 1665
rect -24 1592 10 1626
rect 44 1592 78 1626
rect -24 1553 78 1592
rect -24 1519 10 1553
rect 44 1519 78 1553
rect -24 1480 78 1519
rect -24 1446 10 1480
rect 44 1446 78 1480
rect -24 1406 78 1446
rect -24 1372 10 1406
rect 44 1372 78 1406
rect -24 1332 78 1372
rect -24 1298 10 1332
rect 44 1298 78 1332
rect -24 1258 78 1298
rect -24 1224 10 1258
rect 44 1224 78 1258
rect -24 1184 78 1224
rect -24 1150 10 1184
rect 44 1150 78 1184
rect -24 1110 78 1150
rect -24 1076 10 1110
rect 44 1076 78 1110
rect -24 1036 78 1076
rect -24 1002 10 1036
rect 44 1002 78 1036
rect -24 962 78 1002
rect -24 928 10 962
rect 44 928 78 962
rect -24 888 78 928
rect -24 854 10 888
rect 44 854 78 888
rect -24 814 78 854
rect -24 780 10 814
rect 44 780 78 814
rect -24 740 78 780
rect -24 706 10 740
rect 44 706 78 740
rect -24 666 78 706
rect -24 632 10 666
rect 44 632 78 666
rect -24 592 78 632
rect -24 558 10 592
rect 44 558 78 592
rect -24 518 78 558
rect -24 484 10 518
rect 44 484 78 518
rect -24 444 78 484
rect -24 410 10 444
rect 44 410 78 444
rect -24 370 78 410
rect -24 336 10 370
rect 44 336 78 370
rect -24 296 78 336
rect 175 2073 1555 2107
rect 175 2039 329 2073
rect 363 2039 403 2073
rect 437 2039 477 2073
rect 511 2039 551 2073
rect 585 2039 625 2073
rect 659 2039 699 2073
rect 733 2039 773 2073
rect 807 2039 847 2073
rect 881 2039 921 2073
rect 955 2039 995 2073
rect 1029 2039 1069 2073
rect 1103 2039 1143 2073
rect 1177 2039 1218 2073
rect 1252 2039 1293 2073
rect 1327 2039 1368 2073
rect 1402 2039 1443 2073
rect 1477 2039 1555 2073
rect 175 2029 1555 2039
rect 175 1995 209 2029
rect 243 2005 1555 2029
rect 243 1995 280 2005
rect 175 1966 280 1995
tri 280 1966 319 2005 nw
tri 1411 1966 1450 2005 ne
rect 1450 1966 1555 2005
rect 175 1955 277 1966
tri 277 1963 280 1966 nw
rect 175 1921 209 1955
rect 243 1921 277 1955
rect 175 1881 277 1921
rect 415 1914 421 1966
rect 473 1914 485 1966
rect 537 1957 1337 1966
tri 1450 1963 1453 1966 ne
rect 540 1923 585 1957
rect 619 1923 664 1957
rect 698 1923 742 1957
rect 776 1923 820 1957
rect 854 1923 898 1957
rect 932 1923 976 1957
rect 1010 1923 1054 1957
rect 1088 1923 1132 1957
rect 1166 1923 1210 1957
rect 1244 1923 1288 1957
rect 1322 1923 1337 1957
rect 537 1914 1337 1923
rect 1453 1955 1555 1966
rect 1453 1921 1487 1955
rect 1521 1921 1555 1955
rect 175 1847 209 1881
rect 243 1847 277 1881
rect 175 1807 277 1847
rect 175 1773 209 1807
rect 243 1773 277 1807
rect 175 1733 277 1773
rect 175 1699 209 1733
rect 243 1699 277 1733
rect 175 1659 277 1699
rect 175 1625 209 1659
rect 243 1625 277 1659
rect 175 1585 277 1625
rect 175 1551 209 1585
rect 243 1551 277 1585
rect 175 1511 277 1551
rect 175 1477 209 1511
rect 243 1477 277 1511
rect 175 1437 277 1477
rect 175 1403 209 1437
rect 243 1403 277 1437
rect 175 1363 277 1403
tri 353 1879 356 1882 se
rect 356 1879 402 1885
tri 402 1879 405 1882 sw
rect 353 1873 405 1879
rect 353 1801 405 1821
rect 353 1800 362 1801
rect 396 1800 405 1801
rect 353 1729 405 1748
rect 353 1726 362 1729
rect 396 1726 405 1729
rect 353 1657 405 1674
rect 353 1652 362 1657
rect 396 1652 405 1657
rect 353 1585 405 1600
rect 353 1578 362 1585
rect 396 1578 405 1585
rect 353 1513 405 1526
rect 353 1504 362 1513
rect 396 1504 405 1513
rect 353 1441 405 1452
rect 353 1430 362 1441
rect 396 1430 405 1441
rect 353 1372 405 1378
tri 353 1371 354 1372 ne
rect 354 1371 404 1372
tri 404 1371 405 1372 nw
rect 519 1873 565 1885
rect 519 1839 525 1873
rect 559 1839 565 1873
rect 519 1801 565 1839
rect 519 1767 525 1801
rect 559 1767 565 1801
rect 519 1729 565 1767
rect 519 1695 525 1729
rect 559 1695 565 1729
rect 519 1657 565 1695
rect 519 1623 525 1657
rect 559 1623 565 1657
rect 519 1585 565 1623
rect 519 1551 525 1585
rect 559 1551 565 1585
rect 519 1513 565 1551
rect 519 1479 525 1513
rect 559 1479 565 1513
rect 519 1441 565 1479
rect 519 1407 525 1441
rect 559 1407 565 1441
tri 354 1369 356 1371 ne
rect 356 1369 402 1371
tri 402 1369 404 1371 nw
rect 519 1369 565 1407
tri 679 1879 682 1882 se
rect 682 1879 728 1885
tri 728 1879 731 1882 sw
rect 679 1873 731 1879
rect 679 1801 731 1821
rect 679 1800 688 1801
rect 722 1800 731 1801
rect 679 1729 731 1748
rect 679 1726 688 1729
rect 722 1726 731 1729
rect 679 1657 731 1674
rect 679 1652 688 1657
rect 722 1652 731 1657
rect 679 1585 731 1600
rect 679 1578 688 1585
rect 722 1578 731 1585
rect 679 1513 731 1526
rect 679 1504 688 1513
rect 722 1504 731 1513
rect 679 1441 731 1452
rect 679 1430 688 1441
rect 722 1430 731 1441
rect 679 1372 731 1378
tri 679 1371 680 1372 ne
rect 680 1371 730 1372
tri 730 1371 731 1372 nw
rect 845 1873 891 1885
rect 845 1839 851 1873
rect 885 1839 891 1873
rect 1008 1873 1054 1885
rect 845 1801 891 1839
rect 845 1767 851 1801
rect 885 1767 891 1801
rect 845 1729 891 1767
rect 845 1695 851 1729
rect 885 1695 891 1729
rect 845 1657 891 1695
rect 845 1623 851 1657
rect 885 1623 891 1657
rect 845 1585 891 1623
rect 845 1551 851 1585
rect 885 1551 891 1585
rect 845 1513 891 1551
rect 845 1479 851 1513
rect 885 1479 891 1513
tri 1005 1859 1008 1862 se
rect 1008 1859 1014 1873
rect 1005 1853 1014 1859
rect 1048 1859 1054 1873
rect 1171 1873 1217 1885
tri 1054 1859 1057 1862 sw
rect 1048 1853 1057 1859
rect 1005 1775 1014 1801
rect 1048 1775 1057 1801
rect 1005 1696 1014 1723
rect 1048 1696 1057 1723
rect 1005 1623 1014 1644
rect 1048 1623 1057 1644
rect 1005 1617 1057 1623
rect 1005 1551 1014 1565
rect 1048 1551 1057 1565
rect 1005 1538 1057 1551
rect 1005 1480 1014 1486
tri 1005 1479 1006 1480 ne
rect 1006 1479 1014 1480
rect 1048 1480 1057 1486
rect 1048 1479 1056 1480
tri 1056 1479 1057 1480 nw
rect 1171 1839 1177 1873
rect 1211 1839 1217 1873
rect 1334 1873 1380 1885
rect 1171 1801 1217 1839
rect 1171 1767 1177 1801
rect 1211 1767 1217 1801
rect 1171 1729 1217 1767
rect 1171 1695 1177 1729
rect 1211 1695 1217 1729
rect 1171 1657 1217 1695
rect 1171 1623 1177 1657
rect 1211 1623 1217 1657
rect 1171 1585 1217 1623
rect 1171 1551 1177 1585
rect 1211 1551 1217 1585
rect 1171 1513 1217 1551
rect 1171 1479 1177 1513
rect 1211 1479 1217 1513
tri 1331 1859 1334 1862 se
rect 1334 1859 1340 1873
rect 1331 1853 1340 1859
rect 1374 1859 1380 1873
rect 1453 1882 1555 1921
tri 1380 1859 1383 1862 sw
rect 1374 1853 1383 1859
rect 1331 1775 1340 1801
rect 1374 1775 1383 1801
rect 1331 1696 1340 1723
rect 1374 1696 1383 1723
rect 1331 1623 1340 1644
rect 1374 1623 1383 1644
rect 1331 1617 1383 1623
rect 1331 1551 1340 1565
rect 1374 1551 1383 1565
rect 1331 1538 1383 1551
rect 1331 1480 1340 1486
tri 1331 1479 1332 1480 ne
rect 1332 1479 1340 1480
rect 1374 1480 1383 1486
rect 1374 1479 1380 1480
rect 845 1441 891 1479
tri 1006 1477 1008 1479 ne
rect 845 1407 851 1441
rect 885 1407 891 1441
tri 680 1369 682 1371 ne
rect 682 1369 728 1371
tri 728 1369 730 1371 nw
rect 845 1369 891 1407
rect 175 1329 209 1363
rect 243 1329 277 1363
rect 175 1289 277 1329
rect 175 1255 209 1289
rect 243 1255 277 1289
rect 175 1215 277 1255
rect 175 1181 209 1215
rect 243 1181 277 1215
rect 175 1142 277 1181
rect 175 1108 209 1142
rect 243 1108 277 1142
rect 175 1069 277 1108
rect 175 1035 209 1069
rect 243 1035 277 1069
rect 175 996 277 1035
rect 175 962 209 996
rect 243 962 277 996
rect 175 923 277 962
rect 175 889 209 923
rect 243 889 277 923
rect 175 850 277 889
rect 175 816 209 850
rect 243 816 277 850
rect 175 777 277 816
rect 175 743 209 777
rect 243 743 277 777
rect 175 704 277 743
rect 175 670 209 704
rect 243 670 277 704
rect 175 631 277 670
rect 175 597 209 631
rect 243 597 277 631
rect 175 558 277 597
rect 175 524 209 558
rect 243 524 277 558
rect 175 485 277 524
rect 175 451 209 485
rect 243 451 277 485
rect 356 1335 362 1369
rect 396 1335 402 1369
rect 356 1297 402 1335
rect 356 1263 362 1297
rect 396 1263 402 1297
rect 356 1225 402 1263
rect 356 1191 362 1225
rect 396 1191 402 1225
rect 356 1153 402 1191
rect 356 1119 362 1153
rect 396 1119 402 1153
rect 356 1081 402 1119
rect 356 1047 362 1081
rect 396 1047 402 1081
rect 356 1009 402 1047
rect 356 975 362 1009
rect 396 975 402 1009
rect 356 937 402 975
rect 356 903 362 937
rect 396 903 402 937
rect 356 865 402 903
rect 356 831 362 865
rect 396 831 402 865
rect 356 793 402 831
rect 519 1335 525 1369
rect 559 1335 565 1369
rect 519 1297 565 1335
rect 519 1263 525 1297
rect 559 1263 565 1297
rect 519 1225 565 1263
rect 519 1191 525 1225
rect 559 1191 565 1225
rect 519 1153 565 1191
rect 519 1119 525 1153
rect 559 1119 565 1153
rect 519 1081 565 1119
rect 519 1047 525 1081
rect 559 1047 565 1081
rect 519 1009 565 1047
rect 519 975 525 1009
rect 559 975 565 1009
rect 519 937 565 975
rect 519 903 525 937
rect 559 903 565 937
rect 519 865 565 903
rect 519 831 525 865
rect 559 831 565 865
rect 356 759 362 793
rect 396 759 402 793
rect 356 721 402 759
rect 356 687 362 721
rect 396 687 402 721
rect 356 649 402 687
rect 356 615 362 649
rect 396 615 402 649
rect 356 577 402 615
rect 356 543 362 577
rect 396 543 402 577
rect 356 505 402 543
rect 356 471 362 505
rect 396 471 402 505
rect 356 459 402 471
tri 516 809 519 812 se
rect 519 809 565 831
rect 682 1335 688 1369
rect 722 1335 728 1369
rect 682 1297 728 1335
rect 682 1263 688 1297
rect 722 1263 728 1297
rect 682 1225 728 1263
rect 682 1191 688 1225
rect 722 1191 728 1225
rect 682 1153 728 1191
rect 682 1119 688 1153
rect 722 1119 728 1153
rect 682 1081 728 1119
rect 682 1047 688 1081
rect 722 1047 728 1081
rect 682 1009 728 1047
rect 682 975 688 1009
rect 722 975 728 1009
rect 682 937 728 975
rect 682 903 688 937
rect 722 903 728 937
rect 682 865 728 903
rect 682 831 688 865
rect 722 831 728 865
tri 565 809 568 812 sw
rect 516 803 568 809
rect 516 735 568 751
rect 516 666 568 683
rect 516 597 568 614
rect 516 543 525 545
rect 559 543 568 545
rect 516 528 568 543
rect 516 471 525 476
rect 559 471 568 476
rect 516 470 568 471
tri 516 467 519 470 ne
rect 519 459 565 470
tri 565 467 568 470 nw
rect 682 793 728 831
rect 845 1335 851 1369
rect 885 1335 891 1369
rect 845 1297 891 1335
rect 845 1263 851 1297
rect 885 1263 891 1297
rect 845 1225 891 1263
rect 845 1191 851 1225
rect 885 1191 891 1225
rect 845 1153 891 1191
rect 845 1119 851 1153
rect 885 1119 891 1153
rect 845 1081 891 1119
rect 845 1047 851 1081
rect 885 1047 891 1081
rect 845 1009 891 1047
rect 845 975 851 1009
rect 885 975 891 1009
rect 845 937 891 975
rect 845 903 851 937
rect 885 903 891 937
rect 845 865 891 903
rect 845 831 851 865
rect 885 831 891 865
rect 682 759 688 793
rect 722 759 728 793
rect 682 721 728 759
rect 682 687 688 721
rect 722 687 728 721
rect 682 649 728 687
rect 682 615 688 649
rect 722 615 728 649
rect 682 577 728 615
rect 682 543 688 577
rect 722 543 728 577
rect 682 505 728 543
rect 682 471 688 505
rect 722 471 728 505
rect 682 459 728 471
tri 842 809 845 812 se
rect 845 809 891 831
rect 1008 1441 1054 1479
tri 1054 1477 1056 1479 nw
rect 1008 1407 1014 1441
rect 1048 1407 1054 1441
rect 1008 1369 1054 1407
rect 1008 1335 1014 1369
rect 1048 1335 1054 1369
rect 1008 1297 1054 1335
rect 1008 1263 1014 1297
rect 1048 1263 1054 1297
rect 1008 1225 1054 1263
rect 1008 1191 1014 1225
rect 1048 1191 1054 1225
rect 1008 1153 1054 1191
rect 1008 1119 1014 1153
rect 1048 1119 1054 1153
rect 1008 1081 1054 1119
rect 1008 1047 1014 1081
rect 1048 1047 1054 1081
rect 1008 1009 1054 1047
rect 1008 975 1014 1009
rect 1048 975 1054 1009
rect 1008 937 1054 975
rect 1008 903 1014 937
rect 1048 903 1054 937
rect 1008 865 1054 903
rect 1008 831 1014 865
rect 1048 831 1054 865
tri 891 809 894 812 sw
rect 842 803 894 809
rect 842 735 894 751
rect 842 666 894 683
rect 842 597 894 614
rect 842 543 851 545
rect 885 543 894 545
rect 842 528 894 543
rect 842 471 851 476
rect 885 471 894 476
rect 842 470 894 471
tri 842 467 845 470 ne
rect 845 459 891 470
tri 891 467 894 470 nw
rect 1008 793 1054 831
rect 1171 1441 1217 1479
tri 1332 1477 1334 1479 ne
rect 1171 1407 1177 1441
rect 1211 1407 1217 1441
rect 1171 1369 1217 1407
rect 1171 1335 1177 1369
rect 1211 1335 1217 1369
rect 1171 1297 1217 1335
rect 1171 1263 1177 1297
rect 1211 1263 1217 1297
rect 1171 1225 1217 1263
rect 1171 1191 1177 1225
rect 1211 1191 1217 1225
rect 1171 1153 1217 1191
rect 1171 1119 1177 1153
rect 1211 1119 1217 1153
rect 1171 1081 1217 1119
rect 1171 1047 1177 1081
rect 1211 1047 1217 1081
rect 1171 1009 1217 1047
rect 1171 975 1177 1009
rect 1211 975 1217 1009
rect 1171 937 1217 975
rect 1171 903 1177 937
rect 1211 903 1217 937
rect 1171 865 1217 903
rect 1171 831 1177 865
rect 1211 831 1217 865
rect 1008 759 1014 793
rect 1048 759 1054 793
rect 1008 721 1054 759
rect 1008 687 1014 721
rect 1048 687 1054 721
rect 1008 649 1054 687
rect 1008 615 1014 649
rect 1048 615 1054 649
rect 1008 577 1054 615
rect 1008 543 1014 577
rect 1048 543 1054 577
rect 1008 505 1054 543
rect 1008 471 1014 505
rect 1048 471 1054 505
rect 1008 459 1054 471
tri 1168 809 1171 812 se
rect 1171 809 1217 831
rect 1334 1441 1380 1479
tri 1380 1477 1383 1480 nw
rect 1453 1848 1487 1882
rect 1521 1848 1555 1882
rect 1453 1809 1555 1848
rect 1453 1775 1487 1809
rect 1521 1775 1555 1809
rect 1453 1736 1555 1775
rect 1453 1702 1487 1736
rect 1521 1702 1555 1736
rect 1453 1663 1555 1702
rect 1453 1629 1487 1663
rect 1521 1629 1555 1663
rect 1453 1590 1555 1629
rect 1453 1556 1487 1590
rect 1521 1556 1555 1590
rect 1453 1517 1555 1556
rect 1453 1483 1487 1517
rect 1521 1483 1555 1517
rect 1334 1407 1340 1441
rect 1374 1407 1380 1441
rect 1334 1369 1380 1407
rect 1334 1335 1340 1369
rect 1374 1335 1380 1369
rect 1334 1297 1380 1335
rect 1334 1263 1340 1297
rect 1374 1263 1380 1297
rect 1334 1225 1380 1263
rect 1334 1191 1340 1225
rect 1374 1191 1380 1225
rect 1334 1153 1380 1191
rect 1334 1119 1340 1153
rect 1374 1119 1380 1153
rect 1334 1081 1380 1119
rect 1334 1047 1340 1081
rect 1374 1047 1380 1081
rect 1334 1009 1380 1047
rect 1334 975 1340 1009
rect 1374 975 1380 1009
rect 1334 937 1380 975
rect 1334 903 1340 937
rect 1374 903 1380 937
rect 1334 865 1380 903
rect 1334 831 1340 865
rect 1374 831 1380 865
tri 1217 809 1220 812 sw
rect 1168 803 1220 809
rect 1168 735 1220 751
rect 1168 666 1220 683
rect 1168 597 1220 614
rect 1168 543 1177 545
rect 1211 543 1220 545
rect 1168 528 1220 543
rect 1168 471 1177 476
rect 1211 471 1220 476
rect 1168 470 1220 471
tri 1168 467 1171 470 ne
rect 1171 459 1217 470
tri 1217 467 1220 470 nw
rect 1334 793 1380 831
rect 1334 759 1340 793
rect 1374 759 1380 793
rect 1334 721 1380 759
rect 1334 687 1340 721
rect 1374 687 1380 721
rect 1334 649 1380 687
rect 1334 615 1340 649
rect 1374 615 1380 649
rect 1334 577 1380 615
rect 1334 543 1340 577
rect 1374 543 1380 577
rect 1334 505 1380 543
rect 1334 471 1340 505
rect 1374 471 1380 505
rect 1334 459 1380 471
rect 1453 1444 1555 1483
rect 1453 1410 1487 1444
rect 1521 1410 1555 1444
rect 1453 1371 1555 1410
rect 1453 1337 1487 1371
rect 1521 1337 1555 1371
rect 1453 1298 1555 1337
rect 1453 1264 1487 1298
rect 1521 1264 1555 1298
rect 1453 1225 1555 1264
rect 1453 1191 1487 1225
rect 1521 1191 1555 1225
rect 1453 1151 1555 1191
rect 1453 1117 1487 1151
rect 1521 1117 1555 1151
rect 1453 1077 1555 1117
rect 1453 1043 1487 1077
rect 1521 1043 1555 1077
rect 1453 1003 1555 1043
rect 1453 969 1487 1003
rect 1521 969 1555 1003
rect 1453 929 1555 969
rect 1453 895 1487 929
rect 1521 895 1555 929
rect 1453 855 1555 895
rect 1453 821 1487 855
rect 1521 821 1555 855
rect 1453 781 1555 821
rect 1453 747 1487 781
rect 1521 747 1555 781
rect 1453 707 1555 747
rect 1453 673 1487 707
rect 1521 673 1555 707
rect 1453 633 1555 673
rect 1453 599 1487 633
rect 1521 599 1555 633
rect 1453 559 1555 599
rect 1453 525 1487 559
rect 1521 525 1555 559
rect 1453 485 1555 525
rect 175 423 277 451
rect 1453 451 1487 485
rect 1521 451 1555 485
tri 1450 441 1453 444 se
rect 1453 441 1555 451
tri 1444 435 1450 441 se
rect 1450 435 1555 441
tri 277 423 289 435 sw
tri 1432 423 1444 435 se
rect 1444 423 1555 435
rect 175 411 289 423
tri 289 411 301 423 sw
tri 1420 411 1432 423 se
rect 1432 411 1555 423
rect 175 401 301 411
tri 301 401 311 411 sw
tri 1410 401 1420 411 se
rect 1420 401 1487 411
rect 175 377 1487 401
rect 1521 377 1555 411
rect 175 367 1555 377
rect 175 333 253 367
rect 287 333 347 367
rect 381 333 440 367
rect 474 333 533 367
rect 567 333 609 367
rect 643 333 685 367
rect 719 333 761 367
rect 795 333 837 367
rect 871 333 913 367
rect 947 333 989 367
rect 1023 333 1065 367
rect 1099 333 1140 367
rect 1174 333 1215 367
rect 1249 333 1290 367
rect 1324 333 1365 367
rect 1399 333 1555 367
rect 175 299 1555 333
rect 1641 754 1648 2226
rect 1898 2212 1956 2228
tri 1956 2212 1994 2250 nw
tri 3411 2226 3435 2250 ne
rect 1898 2210 1954 2212
tri 1954 2210 1956 2212 nw
rect 3435 2210 3537 2250
rect 1898 2176 1920 2210
tri 1920 2176 1954 2210 nw
rect 3435 2176 3469 2210
rect 3503 2176 3537 2210
rect 1898 754 1905 2176
tri 1905 2161 1920 2176 nw
rect 3435 2136 3537 2176
rect 1641 715 1905 754
rect 1641 681 1648 715
rect 1682 681 1720 715
rect 1754 681 1792 715
rect 1826 681 1864 715
rect 1898 681 1905 715
rect 1641 642 1905 681
rect 1641 608 1648 642
rect 1682 608 1720 642
rect 1754 608 1792 642
rect 1826 608 1864 642
rect 1898 608 1905 642
rect 1641 569 1905 608
rect 1641 535 1648 569
rect 1682 535 1720 569
rect 1754 535 1792 569
rect 1826 535 1864 569
rect 1898 535 1905 569
rect 1641 496 1905 535
rect 1641 462 1648 496
rect 1682 462 1720 496
rect 1754 462 1792 496
rect 1826 462 1864 496
rect 1898 462 1905 496
rect 1641 423 1905 462
rect 1641 389 1648 423
rect 1682 389 1720 423
rect 1754 389 1792 423
rect 1826 389 1864 423
rect 1898 389 1905 423
rect 1641 350 1905 389
rect 1641 316 1648 350
rect 1682 316 1720 350
rect 1754 316 1792 350
rect 1826 316 1864 350
rect 1898 316 1905 350
rect -24 262 10 296
rect 44 262 78 296
rect -24 222 78 262
rect -24 188 10 222
rect 44 188 78 222
rect 1641 277 1905 316
rect 2058 2073 3288 2107
rect 2058 2039 2212 2073
rect 2246 2039 2286 2073
rect 2320 2039 2360 2073
rect 2394 2039 2434 2073
rect 2468 2039 2508 2073
rect 2542 2039 2582 2073
rect 2616 2039 2656 2073
rect 2690 2039 2730 2073
rect 2764 2039 2804 2073
rect 2838 2039 2878 2073
rect 2912 2039 2952 2073
rect 2986 2039 3026 2073
rect 3060 2039 3101 2073
rect 3135 2039 3176 2073
rect 3210 2039 3288 2073
rect 2058 2029 3288 2039
rect 2058 1995 2092 2029
rect 2126 2005 3288 2029
rect 2126 2001 2201 2005
tri 2201 2001 2205 2005 nw
rect 2126 1999 2199 2001
tri 2199 1999 2201 2001 nw
rect 2126 1995 2191 1999
rect 2058 1991 2191 1995
tri 2191 1991 2199 1999 nw
rect 2058 1988 2188 1991
tri 2188 1988 2191 1991 nw
rect 2058 1963 2163 1988
tri 2163 1963 2188 1988 nw
rect 2058 1955 2160 1963
tri 2160 1960 2163 1963 nw
rect 2058 1921 2092 1955
rect 2126 1921 2160 1955
rect 2058 1881 2160 1921
rect 2291 1914 2297 1966
rect 2349 1914 2361 1966
rect 2413 1957 3055 1966
rect 2416 1923 2461 1957
rect 2495 1923 2540 1957
rect 2574 1923 2619 1957
rect 2653 1923 2697 1957
rect 2731 1923 2775 1957
rect 2809 1923 2853 1957
rect 2887 1923 2931 1957
rect 2965 1923 3009 1957
rect 3043 1923 3055 1957
rect 2413 1914 3055 1923
rect 3186 1953 3211 2005
rect 3263 1953 3288 2005
rect 3186 1921 3220 1953
rect 3254 1921 3288 1953
rect 3186 1920 3288 1921
rect 2058 1847 2092 1881
rect 2126 1847 2160 1881
rect 2058 1807 2160 1847
rect 2058 1773 2092 1807
rect 2126 1773 2160 1807
rect 2058 1733 2160 1773
rect 2058 1699 2092 1733
rect 2126 1699 2160 1733
rect 2058 1659 2160 1699
rect 2058 1625 2092 1659
rect 2126 1625 2160 1659
rect 2058 1585 2160 1625
rect 2058 1551 2092 1585
rect 2126 1551 2160 1585
rect 2058 1511 2160 1551
rect 2058 1477 2092 1511
rect 2126 1477 2160 1511
rect 2058 1437 2160 1477
rect 2058 1403 2092 1437
rect 2126 1403 2160 1437
rect 2058 1363 2160 1403
rect 2058 1329 2092 1363
rect 2126 1329 2160 1363
rect 2058 1289 2160 1329
rect 2058 1255 2092 1289
rect 2126 1255 2160 1289
rect 2058 1215 2160 1255
rect 2240 1873 2286 1885
rect 2240 1839 2246 1873
rect 2280 1839 2286 1873
rect 2240 1801 2286 1839
rect 2240 1767 2246 1801
rect 2280 1767 2286 1801
rect 2240 1729 2286 1767
rect 2240 1695 2246 1729
rect 2280 1695 2286 1729
rect 2240 1657 2286 1695
rect 2240 1623 2246 1657
rect 2280 1623 2286 1657
rect 2240 1585 2286 1623
rect 2240 1551 2246 1585
rect 2280 1551 2286 1585
rect 2240 1513 2286 1551
rect 2240 1479 2246 1513
rect 2280 1479 2286 1513
rect 2240 1441 2286 1479
rect 2240 1407 2246 1441
rect 2280 1407 2286 1441
rect 2240 1369 2286 1407
rect 2240 1335 2246 1369
rect 2280 1335 2286 1369
rect 2240 1297 2286 1335
rect 2240 1263 2246 1297
rect 2280 1263 2286 1297
rect 2058 1181 2092 1215
rect 2126 1181 2160 1215
rect 2058 1142 2160 1181
rect 2058 1108 2092 1142
rect 2126 1108 2160 1142
rect 2058 1069 2160 1108
rect 2058 1035 2092 1069
rect 2126 1035 2160 1069
rect 2058 996 2160 1035
rect 2058 962 2092 996
rect 2126 962 2160 996
rect 2058 923 2160 962
rect 2058 889 2092 923
rect 2126 889 2160 923
tri 2237 1232 2240 1235 se
rect 2240 1232 2286 1263
rect 2403 1873 2449 1885
rect 2403 1839 2409 1873
rect 2443 1839 2449 1873
rect 2403 1801 2449 1839
rect 2403 1767 2409 1801
rect 2443 1767 2449 1801
rect 2403 1729 2449 1767
rect 2403 1695 2409 1729
rect 2443 1695 2449 1729
rect 2403 1657 2449 1695
rect 2403 1623 2409 1657
rect 2443 1623 2449 1657
rect 2403 1585 2449 1623
rect 2403 1551 2409 1585
rect 2443 1551 2449 1585
rect 2403 1513 2449 1551
rect 2403 1479 2409 1513
rect 2443 1479 2449 1513
rect 2403 1441 2449 1479
rect 2403 1407 2409 1441
rect 2443 1407 2449 1441
rect 2403 1369 2449 1407
rect 2403 1335 2409 1369
rect 2443 1335 2449 1369
rect 2403 1297 2449 1335
rect 2403 1263 2409 1297
rect 2443 1263 2449 1297
tri 2286 1232 2289 1235 sw
rect 2237 1226 2289 1232
rect 2237 1157 2289 1174
rect 2237 1088 2289 1105
rect 2237 1019 2289 1036
rect 2237 950 2289 967
rect 2237 892 2289 898
tri 2237 889 2240 892 ne
rect 2058 850 2160 889
rect 2058 816 2092 850
rect 2126 816 2160 850
rect 2058 777 2160 816
rect 2058 743 2092 777
rect 2126 743 2160 777
rect 2058 704 2160 743
rect 2058 670 2092 704
rect 2126 670 2160 704
rect 2058 631 2160 670
rect 2058 597 2092 631
rect 2126 597 2160 631
rect 2058 558 2160 597
rect 2058 524 2092 558
rect 2126 524 2160 558
rect 2058 485 2160 524
rect 2058 451 2092 485
rect 2126 451 2160 485
rect 2240 865 2286 892
tri 2286 889 2289 892 nw
rect 2403 1225 2449 1263
rect 2566 1873 2612 1885
rect 2566 1839 2572 1873
rect 2606 1839 2612 1873
rect 2566 1801 2612 1839
rect 2566 1767 2572 1801
rect 2606 1767 2612 1801
rect 2566 1729 2612 1767
rect 2566 1695 2572 1729
rect 2606 1695 2612 1729
rect 2566 1657 2612 1695
rect 2566 1623 2572 1657
rect 2606 1623 2612 1657
rect 2566 1585 2612 1623
rect 2566 1551 2572 1585
rect 2606 1551 2612 1585
rect 2566 1513 2612 1551
rect 2566 1479 2572 1513
rect 2606 1479 2612 1513
rect 2566 1441 2612 1479
rect 2566 1407 2572 1441
rect 2606 1407 2612 1441
rect 2566 1369 2612 1407
rect 2566 1335 2572 1369
rect 2606 1335 2612 1369
rect 2566 1297 2612 1335
rect 2566 1263 2572 1297
rect 2606 1263 2612 1297
rect 2403 1191 2409 1225
rect 2443 1191 2449 1225
rect 2403 1153 2449 1191
rect 2403 1119 2409 1153
rect 2443 1119 2449 1153
rect 2403 1081 2449 1119
rect 2403 1047 2409 1081
rect 2443 1047 2449 1081
rect 2403 1009 2449 1047
rect 2403 975 2409 1009
rect 2443 975 2449 1009
rect 2403 937 2449 975
rect 2403 903 2409 937
rect 2443 903 2449 937
rect 2240 831 2246 865
rect 2280 831 2286 865
rect 2240 793 2286 831
rect 2403 865 2449 903
tri 2563 1232 2566 1235 se
rect 2566 1232 2612 1263
rect 2729 1873 2775 1885
rect 2729 1839 2735 1873
rect 2769 1839 2775 1873
rect 2729 1801 2775 1839
rect 2729 1767 2735 1801
rect 2769 1767 2775 1801
rect 2729 1729 2775 1767
rect 2729 1695 2735 1729
rect 2769 1695 2775 1729
rect 2729 1657 2775 1695
rect 2729 1623 2735 1657
rect 2769 1623 2775 1657
rect 2729 1585 2775 1623
rect 2729 1551 2735 1585
rect 2769 1551 2775 1585
rect 2729 1513 2775 1551
rect 2729 1479 2735 1513
rect 2769 1479 2775 1513
rect 2729 1441 2775 1479
rect 2729 1407 2735 1441
rect 2769 1407 2775 1441
rect 2729 1369 2775 1407
rect 2729 1335 2735 1369
rect 2769 1335 2775 1369
rect 2729 1297 2775 1335
rect 2729 1263 2735 1297
rect 2769 1263 2775 1297
tri 2612 1232 2615 1235 sw
rect 2563 1226 2615 1232
rect 2563 1157 2615 1174
rect 2563 1088 2615 1105
rect 2563 1019 2615 1036
rect 2563 950 2615 967
rect 2563 892 2615 898
tri 2563 889 2566 892 ne
rect 2403 831 2409 865
rect 2443 831 2449 865
rect 2240 759 2246 793
rect 2280 759 2286 793
rect 2240 721 2286 759
rect 2240 687 2246 721
rect 2280 687 2286 721
rect 2240 649 2286 687
rect 2240 615 2246 649
rect 2280 615 2286 649
rect 2240 577 2286 615
rect 2240 543 2246 577
rect 2280 543 2286 577
rect 2240 505 2286 543
rect 2240 471 2246 505
rect 2280 471 2286 505
rect 2240 459 2286 471
tri 2400 809 2403 812 se
rect 2403 809 2449 831
rect 2566 865 2612 892
tri 2612 889 2615 892 nw
rect 2729 1225 2775 1263
rect 2892 1873 2938 1885
rect 2892 1839 2898 1873
rect 2932 1839 2938 1873
rect 2892 1801 2938 1839
rect 2892 1767 2898 1801
rect 2932 1767 2938 1801
rect 2892 1729 2938 1767
rect 2892 1695 2898 1729
rect 2932 1695 2938 1729
rect 2892 1657 2938 1695
rect 2892 1623 2898 1657
rect 2932 1623 2938 1657
rect 2892 1585 2938 1623
rect 2892 1551 2898 1585
rect 2932 1551 2938 1585
rect 2892 1513 2938 1551
rect 2892 1479 2898 1513
rect 2932 1479 2938 1513
rect 2892 1441 2938 1479
rect 2892 1407 2898 1441
rect 2932 1407 2938 1441
rect 2892 1369 2938 1407
rect 2892 1335 2898 1369
rect 2932 1335 2938 1369
rect 2892 1297 2938 1335
rect 2892 1263 2898 1297
rect 2932 1263 2938 1297
rect 2729 1191 2735 1225
rect 2769 1191 2775 1225
rect 2729 1153 2775 1191
rect 2729 1119 2735 1153
rect 2769 1119 2775 1153
rect 2729 1081 2775 1119
rect 2729 1047 2735 1081
rect 2769 1047 2775 1081
rect 2729 1009 2775 1047
rect 2729 975 2735 1009
rect 2769 975 2775 1009
rect 2729 937 2775 975
rect 2729 903 2735 937
rect 2769 903 2775 937
rect 2566 831 2572 865
rect 2606 831 2612 865
tri 2449 809 2452 812 sw
rect 2400 803 2452 809
rect 2400 735 2452 751
rect 2400 666 2452 683
rect 2400 597 2452 614
rect 2400 543 2409 545
rect 2443 543 2452 545
rect 2400 528 2452 543
rect 2400 471 2409 476
rect 2443 471 2452 476
rect 2400 470 2452 471
tri 2400 467 2403 470 ne
rect 2403 459 2449 470
tri 2449 467 2452 470 nw
rect 2566 793 2612 831
rect 2729 865 2775 903
tri 2889 1232 2892 1235 se
rect 2892 1232 2938 1263
rect 3055 1873 3101 1885
rect 3055 1839 3061 1873
rect 3095 1839 3101 1873
rect 3055 1801 3101 1839
rect 3055 1767 3061 1801
rect 3095 1767 3101 1801
rect 3055 1729 3101 1767
rect 3055 1695 3061 1729
rect 3095 1695 3101 1729
rect 3055 1657 3101 1695
rect 3055 1623 3061 1657
rect 3095 1623 3101 1657
rect 3055 1585 3101 1623
rect 3055 1551 3061 1585
rect 3095 1551 3101 1585
rect 3055 1513 3101 1551
rect 3055 1479 3061 1513
rect 3095 1479 3101 1513
rect 3055 1441 3101 1479
rect 3055 1407 3061 1441
rect 3095 1407 3101 1441
rect 3055 1369 3101 1407
rect 3055 1335 3061 1369
rect 3095 1335 3101 1369
rect 3055 1297 3101 1335
rect 3055 1263 3061 1297
rect 3095 1263 3101 1297
tri 2938 1232 2941 1235 sw
rect 2889 1226 2941 1232
rect 2889 1157 2941 1174
rect 2889 1088 2941 1105
rect 2889 1019 2941 1036
rect 2889 950 2941 967
rect 2889 892 2941 898
tri 2889 889 2892 892 ne
rect 2729 831 2735 865
rect 2769 831 2775 865
rect 2566 759 2572 793
rect 2606 759 2612 793
rect 2566 721 2612 759
rect 2566 687 2572 721
rect 2606 687 2612 721
rect 2566 649 2612 687
rect 2566 615 2572 649
rect 2606 615 2612 649
rect 2566 577 2612 615
rect 2566 543 2572 577
rect 2606 543 2612 577
rect 2566 505 2612 543
rect 2566 471 2572 505
rect 2606 471 2612 505
rect 2566 459 2612 471
tri 2726 809 2729 812 se
rect 2729 809 2775 831
rect 2892 865 2938 892
tri 2938 889 2941 892 nw
rect 3055 1225 3101 1263
rect 3055 1191 3061 1225
rect 3095 1191 3101 1225
rect 3055 1153 3101 1191
rect 3055 1119 3061 1153
rect 3095 1119 3101 1153
rect 3055 1081 3101 1119
rect 3055 1047 3061 1081
rect 3095 1047 3101 1081
rect 3055 1009 3101 1047
rect 3055 975 3061 1009
rect 3095 975 3101 1009
rect 3055 937 3101 975
rect 3055 903 3061 937
rect 3095 903 3101 937
rect 2892 831 2898 865
rect 2932 831 2938 865
tri 2775 809 2778 812 sw
rect 2726 803 2778 809
rect 2726 735 2778 751
rect 2726 666 2778 683
rect 2726 597 2778 614
rect 2726 543 2735 545
rect 2769 543 2778 545
rect 2726 528 2778 543
rect 2726 471 2735 476
rect 2769 471 2778 476
rect 2726 470 2778 471
tri 2726 467 2729 470 ne
rect 2729 459 2775 470
tri 2775 467 2778 470 nw
rect 2892 793 2938 831
rect 3055 865 3101 903
rect 3055 831 3061 865
rect 3095 831 3101 865
rect 2892 759 2898 793
rect 2932 759 2938 793
rect 2892 721 2938 759
rect 2892 687 2898 721
rect 2932 687 2938 721
rect 2892 649 2938 687
rect 2892 615 2898 649
rect 2932 615 2938 649
rect 2892 577 2938 615
rect 2892 543 2898 577
rect 2932 543 2938 577
rect 2892 505 2938 543
rect 2892 471 2898 505
rect 2932 471 2938 505
rect 2892 459 2938 471
tri 3052 809 3055 812 se
rect 3055 809 3101 831
rect 3186 1868 3211 1920
rect 3263 1868 3288 1920
rect 3186 1848 3220 1868
rect 3254 1848 3288 1868
rect 3186 1835 3288 1848
rect 3186 1783 3211 1835
rect 3263 1783 3288 1835
rect 3186 1775 3220 1783
rect 3254 1775 3288 1783
rect 3186 1736 3288 1775
rect 3186 1702 3220 1736
rect 3254 1702 3288 1736
rect 3186 1663 3288 1702
rect 3186 1629 3220 1663
rect 3254 1629 3288 1663
rect 3186 1590 3288 1629
rect 3186 1556 3220 1590
rect 3254 1556 3288 1590
rect 3186 1517 3288 1556
rect 3186 1483 3220 1517
rect 3254 1483 3288 1517
rect 3186 1444 3288 1483
rect 3186 1410 3220 1444
rect 3254 1410 3288 1444
rect 3186 1371 3288 1410
rect 3186 1337 3220 1371
rect 3254 1337 3288 1371
rect 3186 1298 3288 1337
rect 3186 1264 3220 1298
rect 3254 1264 3288 1298
rect 3186 1225 3288 1264
rect 3186 1191 3220 1225
rect 3254 1191 3288 1225
rect 3186 1151 3288 1191
rect 3186 1117 3220 1151
rect 3254 1117 3288 1151
rect 3186 1077 3288 1117
rect 3186 1043 3220 1077
rect 3254 1043 3288 1077
rect 3186 1003 3288 1043
rect 3186 969 3220 1003
rect 3254 969 3288 1003
rect 3186 929 3288 969
rect 3186 895 3220 929
rect 3254 895 3288 929
rect 3186 855 3288 895
rect 3186 821 3220 855
rect 3254 821 3288 855
tri 3101 809 3104 812 sw
rect 3052 803 3104 809
rect 3052 735 3104 751
rect 3052 666 3104 683
rect 3052 597 3104 614
rect 3052 543 3061 545
rect 3095 543 3104 545
rect 3052 528 3104 543
rect 3052 471 3061 476
rect 3095 471 3104 476
rect 3052 470 3104 471
tri 3052 467 3055 470 ne
rect 3055 459 3101 470
tri 3101 467 3104 470 nw
rect 3186 781 3288 821
rect 3186 747 3220 781
rect 3254 747 3288 781
rect 3186 707 3288 747
rect 3186 673 3220 707
rect 3254 673 3288 707
rect 3186 633 3288 673
rect 3186 599 3220 633
rect 3254 599 3288 633
rect 3186 559 3288 599
rect 3186 525 3220 559
rect 3254 525 3288 559
rect 3186 485 3288 525
rect 2058 441 2160 451
rect 3186 451 3220 485
rect 3254 451 3288 485
tri 3185 446 3186 447 se
rect 3186 446 3288 451
tri 2160 441 2165 446 sw
tri 3180 441 3185 446 se
rect 3185 441 3288 446
rect 2058 411 2165 441
tri 2165 411 2195 441 sw
tri 3150 411 3180 441 se
rect 3180 411 3288 441
rect 2058 401 2195 411
tri 2195 401 2205 411 sw
tri 3140 401 3150 411 se
rect 3150 401 3220 411
rect 2058 377 3220 401
rect 3254 377 3288 411
rect 2058 367 3288 377
rect 2058 333 2136 367
rect 2170 333 2230 367
rect 2264 333 2323 367
rect 2357 333 2416 367
rect 2450 333 2492 367
rect 2526 333 2568 367
rect 2602 333 2644 367
rect 2678 333 2720 367
rect 2754 333 2796 367
rect 2830 333 2872 367
rect 2906 333 2948 367
rect 2982 333 3023 367
rect 3057 333 3098 367
rect 3132 333 3288 367
rect 2058 299 3288 333
rect 3435 2102 3469 2136
rect 3503 2102 3537 2136
rect 3435 2062 3537 2102
rect 3435 2028 3469 2062
rect 3503 2028 3537 2062
rect 3435 1988 3537 2028
rect 3435 1954 3469 1988
rect 3503 1954 3537 1988
rect 3435 1914 3537 1954
rect 3435 1880 3469 1914
rect 3503 1880 3537 1914
rect 3435 1840 3537 1880
rect 3435 1806 3469 1840
rect 3503 1806 3537 1840
rect 3435 1766 3537 1806
rect 3435 1732 3469 1766
rect 3503 1732 3537 1766
rect 3435 1692 3537 1732
rect 3435 1658 3469 1692
rect 3503 1658 3537 1692
rect 3435 1618 3537 1658
rect 3435 1584 3469 1618
rect 3503 1584 3537 1618
rect 3435 1544 3537 1584
rect 3435 1510 3469 1544
rect 3503 1510 3537 1544
rect 3435 1470 3537 1510
rect 3435 1436 3469 1470
rect 3503 1436 3537 1470
rect 3435 1396 3537 1436
rect 3435 1362 3469 1396
rect 3503 1362 3537 1396
rect 3435 1322 3537 1362
rect 3435 1288 3469 1322
rect 3503 1288 3537 1322
rect 3435 1248 3537 1288
rect 3435 1214 3469 1248
rect 3503 1214 3537 1248
rect 3435 1174 3537 1214
rect 3435 1140 3469 1174
rect 3503 1140 3537 1174
rect 3435 1100 3537 1140
rect 3435 1066 3469 1100
rect 3503 1066 3537 1100
rect 3435 1026 3537 1066
rect 3435 992 3469 1026
rect 3503 992 3537 1026
rect 3435 952 3537 992
rect 3435 918 3469 952
rect 3503 918 3537 952
rect 3435 879 3537 918
rect 3435 845 3469 879
rect 3503 845 3537 879
rect 3435 806 3537 845
rect 3435 772 3469 806
rect 3503 772 3537 806
rect 3435 733 3537 772
rect 3435 699 3469 733
rect 3503 699 3537 733
rect 3435 660 3537 699
rect 3435 626 3469 660
rect 3503 626 3537 660
rect 3435 587 3537 626
rect 3435 553 3469 587
rect 3503 553 3537 587
rect 3435 514 3537 553
rect 3435 480 3469 514
rect 3503 480 3537 514
rect 3435 441 3537 480
rect 3435 407 3469 441
rect 3503 407 3537 441
rect 3435 368 3537 407
rect 3435 334 3469 368
rect 3503 334 3537 368
rect 1641 243 1648 277
rect 1682 243 1720 277
rect 1754 243 1792 277
rect 1826 243 1864 277
rect 1898 243 1905 277
rect 1641 222 1905 243
rect 3435 295 3537 334
rect 3435 261 3469 295
rect 3503 261 3537 295
tri 1905 222 1913 230 sw
rect 3435 222 3537 261
tri 1639 204 1641 206 se
rect 1641 204 1913 222
rect -24 170 78 188
tri 1607 172 1639 204 se
rect 1639 172 1648 204
tri 78 170 80 172 sw
tri 1605 170 1607 172 se
rect 1607 170 1648 172
rect 1682 170 1720 204
rect 1754 170 1792 204
rect 1826 170 1864 204
rect 1898 188 1913 204
tri 1913 188 1947 222 sw
rect 3435 188 3469 222
rect 3503 188 3537 222
rect 1898 180 1947 188
tri 1947 180 1955 188 sw
rect 1898 170 1955 180
rect -24 156 80 170
tri 80 156 94 170 sw
tri 1591 156 1605 170 se
rect 1605 156 1955 170
tri 1955 156 1979 180 sw
tri 3419 156 3435 172 se
rect 3435 156 3537 188
rect -24 148 94 156
rect -24 114 10 148
rect 44 138 94 148
tri 94 138 112 156 sw
tri 1573 138 1591 156 se
rect 1591 138 1979 156
tri 1979 138 1997 156 sw
tri 3409 146 3419 156 se
rect 3419 146 3537 156
tri 3401 138 3409 146 se
rect 3409 138 3537 146
rect 44 114 3537 138
rect -24 104 3537 114
rect -24 70 128 104
rect 162 70 201 104
rect 235 70 274 104
rect 308 70 347 104
rect 381 70 420 104
rect 454 70 493 104
rect 527 70 566 104
rect 600 70 639 104
rect 673 70 712 104
rect 746 70 785 104
rect 819 70 858 104
rect 892 70 931 104
rect 965 70 1004 104
rect 1038 70 1077 104
rect 1111 70 1150 104
rect 1184 70 1223 104
rect 1257 70 1296 104
rect 1330 70 1369 104
rect 1403 70 1442 104
rect 1476 70 1515 104
rect 1549 70 1588 104
rect 1622 70 1661 104
rect 1695 70 1734 104
rect 1768 70 1807 104
rect 1841 70 1880 104
rect 1914 70 1953 104
rect 1987 70 2026 104
rect 2060 70 2099 104
rect 2133 70 2172 104
rect 2206 70 2245 104
rect 2279 70 2318 104
rect 2352 70 2391 104
rect 2425 70 2464 104
rect 2498 70 2537 104
rect 2571 70 2611 104
rect 2645 70 2685 104
rect 2719 70 2759 104
rect 2793 70 2833 104
rect 2867 70 2907 104
rect 2941 70 2981 104
rect 3015 70 3055 104
rect 3089 70 3129 104
rect 3163 70 3203 104
rect 3237 70 3277 104
rect 3311 70 3351 104
rect 3385 70 3425 104
rect 3459 70 3537 104
rect -24 36 3537 70
rect 3750 2328 10257 2362
rect 3750 2294 3828 2328
rect 3862 2294 3922 2328
rect 3956 2294 4015 2328
rect 4049 2294 4108 2328
rect 4142 2294 4184 2328
rect 4218 2294 4258 2328
rect 4292 2294 4332 2328
rect 4366 2294 4406 2328
rect 4440 2294 4480 2328
rect 4514 2294 4554 2328
rect 4588 2294 4628 2328
rect 4662 2294 4702 2328
rect 4736 2294 4776 2328
rect 4810 2294 4850 2328
rect 4884 2294 4924 2328
rect 4958 2294 4998 2328
rect 5032 2294 5072 2328
rect 5106 2294 5146 2328
rect 5180 2294 5220 2328
rect 5254 2294 5294 2328
rect 5328 2294 5368 2328
rect 5402 2294 5442 2328
rect 5476 2294 5516 2328
rect 5550 2294 5590 2328
rect 5624 2294 5663 2328
rect 5697 2294 5736 2328
rect 5770 2294 5809 2328
rect 5843 2294 5882 2328
rect 5916 2294 5955 2328
rect 5989 2294 6028 2328
rect 6062 2294 6101 2328
rect 6135 2294 6174 2328
rect 6208 2294 6247 2328
rect 6281 2294 6320 2328
rect 6354 2294 6393 2328
rect 6427 2294 6466 2328
rect 6500 2294 6539 2328
rect 6573 2294 6612 2328
rect 6646 2294 6685 2328
rect 6719 2294 6758 2328
rect 6792 2294 6956 2328
rect 6990 2294 7028 2328
rect 7062 2294 7100 2328
rect 7134 2294 7172 2328
rect 7206 2294 7244 2328
rect 7278 2294 7316 2328
rect 7350 2294 7388 2328
rect 7422 2294 7460 2328
rect 7494 2294 7532 2328
rect 7566 2294 7604 2328
rect 7638 2294 7676 2328
rect 7710 2294 7748 2328
rect 7782 2294 7820 2328
rect 7854 2294 7892 2328
rect 7926 2294 7964 2328
rect 7998 2294 8036 2328
rect 8070 2294 8108 2328
rect 8142 2294 8181 2328
rect 8215 2294 8254 2328
rect 8288 2294 8327 2328
rect 8361 2294 8400 2328
rect 8434 2294 8473 2328
rect 8507 2294 8546 2328
rect 8580 2294 8619 2328
rect 8653 2294 8692 2328
rect 8726 2294 8765 2328
rect 8799 2294 8838 2328
rect 8872 2294 8911 2328
rect 8945 2294 8984 2328
rect 9018 2294 9057 2328
rect 9091 2294 9133 2328
rect 9167 2294 9205 2328
rect 9239 2294 9277 2328
rect 9311 2294 9349 2328
rect 9383 2294 9421 2328
rect 9455 2294 9493 2328
rect 9527 2294 9565 2328
rect 9599 2294 9637 2328
rect 9671 2294 9709 2328
rect 9743 2294 9781 2328
rect 9815 2294 9853 2328
rect 9887 2294 9926 2328
rect 9960 2294 9999 2328
rect 10033 2294 10072 2328
rect 10106 2294 10145 2328
rect 10179 2294 10257 2328
rect 3750 2284 10257 2294
rect 3750 2260 6876 2284
rect 3750 2250 3876 2260
tri 3876 2250 3886 2260 nw
tri 6808 2250 6818 2260 ne
rect 6818 2250 6876 2260
rect 6910 2260 10257 2284
rect 6910 2250 6958 2260
rect 3750 2210 3852 2250
tri 3852 2226 3876 2250 nw
tri 6818 2226 6842 2250 ne
rect 6842 2226 6958 2250
tri 6958 2226 6992 2260 nw
tri 10121 2226 10155 2260 ne
rect 3750 2176 3784 2210
rect 3818 2176 3852 2210
rect 3750 2137 3852 2176
rect 3750 2103 3784 2137
rect 3818 2103 3852 2137
rect 3750 2064 3852 2103
rect 6842 2210 6944 2226
tri 6944 2212 6958 2226 nw
rect 10155 2212 10257 2260
rect 6842 2176 6876 2210
rect 6910 2176 6944 2210
rect 6842 2136 6944 2176
rect 6842 2102 6876 2136
rect 6910 2102 6944 2136
rect 10155 2178 10189 2212
rect 10223 2178 10257 2212
rect 10155 2140 10257 2178
rect 3750 2030 3784 2064
rect 3818 2030 3852 2064
rect 3750 2005 3852 2030
rect 3750 1953 3775 2005
rect 3827 1953 3852 2005
rect 3750 1920 3852 1953
rect 3750 1868 3775 1920
rect 3827 1868 3852 1920
rect 3750 1845 3852 1868
rect 3750 1835 3784 1845
rect 3818 1835 3852 1845
rect 3750 1783 3775 1835
rect 3827 1783 3852 1835
rect 3750 1772 3852 1783
rect 3750 1738 3784 1772
rect 3818 1738 3852 1772
rect 3750 1699 3852 1738
rect 3750 1665 3784 1699
rect 3818 1665 3852 1699
rect 3750 1626 3852 1665
rect 3750 1592 3784 1626
rect 3818 1592 3852 1626
rect 3750 1553 3852 1592
rect 3750 1519 3784 1553
rect 3818 1519 3852 1553
rect 3750 1480 3852 1519
rect 3750 1446 3784 1480
rect 3818 1446 3852 1480
rect 3750 1407 3852 1446
rect 3750 1373 3784 1407
rect 3818 1373 3852 1407
rect 3750 1334 3852 1373
rect 3750 1300 3784 1334
rect 3818 1300 3852 1334
rect 3750 1261 3852 1300
rect 3750 1227 3784 1261
rect 3818 1227 3852 1261
rect 3750 1188 3852 1227
rect 3750 1154 3784 1188
rect 3818 1154 3852 1188
rect 3750 1115 3852 1154
rect 3750 1081 3784 1115
rect 3818 1081 3852 1115
rect 3750 1042 3852 1081
rect 3750 1008 3784 1042
rect 3818 1008 3852 1042
rect 3750 969 3852 1008
rect 3750 935 3784 969
rect 3818 935 3852 969
rect 3750 896 3852 935
rect 3750 862 3784 896
rect 3818 862 3852 896
rect 3750 822 3852 862
rect 3750 788 3784 822
rect 3818 788 3852 822
rect 3999 2073 6695 2079
rect 3999 2039 4099 2073
rect 4133 2039 4179 2073
rect 4213 2039 4252 2073
rect 4286 2039 4325 2073
rect 4359 2039 4398 2073
rect 4432 2039 4471 2073
rect 4505 2039 4544 2073
rect 4578 2039 4617 2073
rect 4651 2039 4690 2073
rect 4724 2039 4763 2073
rect 4797 2039 4836 2073
rect 4870 2039 4909 2073
rect 4943 2039 4982 2073
rect 5016 2039 5055 2073
rect 5089 2039 5128 2073
rect 5162 2039 5201 2073
rect 5235 2039 5274 2073
rect 5308 2039 5347 2073
rect 5381 2039 5420 2073
rect 5454 2039 5493 2073
rect 5527 2039 5566 2073
rect 5600 2039 5639 2073
rect 5673 2039 5712 2073
rect 5746 2039 5785 2073
rect 5819 2039 5858 2073
rect 5892 2039 5931 2073
rect 5965 2039 6004 2073
rect 6038 2039 6077 2073
rect 6111 2039 6150 2073
rect 6184 2039 6223 2073
rect 6257 2039 6295 2073
rect 6329 2039 6367 2073
rect 6401 2039 6439 2073
rect 6473 2039 6511 2073
rect 6545 2039 6583 2073
rect 6617 2039 6695 2073
rect 3999 2033 6695 2039
rect 3999 2028 4074 2033
tri 4074 2028 4079 2033 nw
rect 3999 2001 4047 2028
tri 4047 2001 4074 2028 nw
rect 6649 2001 6695 2033
rect 3999 1999 4045 2001
tri 4045 1999 4047 2001 nw
rect 3999 1965 4005 1999
rect 4039 1965 4045 1999
rect 6649 1967 6655 2001
rect 6689 1967 6695 2001
rect 3999 1925 4045 1965
rect 3999 1891 4005 1925
rect 4039 1891 4045 1925
rect 4164 1957 4612 1966
rect 4164 1923 4176 1957
rect 4210 1923 4250 1957
rect 4284 1923 4323 1957
rect 4357 1923 4396 1957
rect 4430 1923 4469 1957
rect 4503 1923 4542 1957
rect 4576 1923 4612 1957
rect 4164 1914 4612 1923
rect 4664 1914 4676 1966
rect 4728 1914 4734 1966
rect 5447 1957 5897 1966
rect 5447 1923 5459 1957
rect 5493 1923 5535 1957
rect 5569 1923 5611 1957
rect 5645 1923 5687 1957
rect 5721 1923 5763 1957
rect 5797 1923 5838 1957
rect 5872 1923 5897 1957
rect 5447 1914 5897 1923
rect 5949 1914 5976 1966
rect 6028 1914 6034 1966
rect 6649 1926 6695 1967
rect 3999 1851 4045 1891
rect 6649 1892 6655 1926
rect 6689 1892 6695 1926
rect 3999 1817 4005 1851
rect 4039 1817 4045 1851
rect 3999 1777 4045 1817
rect 3999 1743 4005 1777
rect 4039 1743 4045 1777
rect 3999 1703 4045 1743
rect 3999 1669 4005 1703
rect 4039 1669 4045 1703
rect 3999 1629 4045 1669
rect 3999 1595 4005 1629
rect 4039 1595 4045 1629
rect 3999 1555 4045 1595
rect 3999 1521 4005 1555
rect 4039 1521 4045 1555
rect 3999 1481 4045 1521
rect 3999 1447 4005 1481
rect 4039 1447 4045 1481
rect 3999 1407 4045 1447
rect 3999 1373 4005 1407
rect 4039 1373 4045 1407
rect 3999 1333 4045 1373
rect 3999 1299 4005 1333
rect 4039 1299 4045 1333
rect 3999 1259 4045 1299
rect 3999 1225 4005 1259
rect 4039 1225 4045 1259
rect 3999 1185 4045 1225
rect 3999 1151 4005 1185
rect 4039 1151 4045 1185
rect 3999 1111 4045 1151
rect 3999 1077 4005 1111
rect 4039 1077 4045 1111
rect 3999 1037 4045 1077
rect 3999 1003 4005 1037
rect 4039 1003 4045 1037
rect 3999 963 4045 1003
rect 3999 929 4005 963
rect 4039 929 4045 963
rect 3999 889 4045 929
rect 3999 855 4005 889
rect 4039 855 4045 889
rect 3999 814 4045 855
rect 3750 748 3852 788
rect 3750 714 3784 748
rect 3818 714 3852 748
rect 3750 674 3852 714
rect 3750 640 3784 674
rect 3818 640 3852 674
rect 3750 600 3852 640
rect 3750 566 3784 600
rect 3818 566 3852 600
rect 3750 526 3852 566
rect 3750 492 3784 526
rect 3818 492 3852 526
rect 3750 452 3852 492
tri 3996 809 3999 812 se
rect 3999 809 4005 814
rect 3996 803 4005 809
rect 4039 811 4045 814
rect 4125 1873 4171 1885
rect 4125 1839 4131 1873
rect 4165 1839 4171 1873
rect 4125 1801 4171 1839
rect 4125 1767 4131 1801
rect 4165 1767 4171 1801
rect 4125 1729 4171 1767
rect 4125 1695 4131 1729
rect 4165 1695 4171 1729
rect 4125 1657 4171 1695
rect 4125 1623 4131 1657
rect 4165 1623 4171 1657
rect 4125 1585 4171 1623
rect 4125 1551 4131 1585
rect 4165 1551 4171 1585
rect 4125 1513 4171 1551
rect 4125 1479 4131 1513
rect 4165 1479 4171 1513
rect 4125 1441 4171 1479
rect 4125 1407 4131 1441
rect 4165 1407 4171 1441
rect 4125 1369 4171 1407
rect 4125 1335 4131 1369
rect 4165 1335 4171 1369
rect 4125 1297 4171 1335
rect 4125 1263 4131 1297
rect 4165 1263 4171 1297
rect 4125 1225 4171 1263
rect 4288 1873 4334 1885
rect 4288 1839 4294 1873
rect 4328 1839 4334 1873
rect 4288 1801 4334 1839
rect 4288 1767 4294 1801
rect 4328 1767 4334 1801
rect 4288 1729 4334 1767
rect 4288 1695 4294 1729
rect 4328 1695 4334 1729
rect 4288 1657 4334 1695
rect 4288 1623 4294 1657
rect 4328 1623 4334 1657
rect 4288 1585 4334 1623
rect 4288 1551 4294 1585
rect 4328 1551 4334 1585
rect 4288 1513 4334 1551
rect 4288 1479 4294 1513
rect 4328 1479 4334 1513
rect 4288 1441 4334 1479
rect 4288 1407 4294 1441
rect 4328 1407 4334 1441
rect 4288 1369 4334 1407
rect 4288 1335 4294 1369
rect 4328 1335 4334 1369
rect 4288 1297 4334 1335
rect 4288 1263 4294 1297
rect 4328 1263 4334 1297
rect 4125 1191 4131 1225
rect 4165 1191 4171 1225
rect 4125 1153 4171 1191
rect 4125 1119 4131 1153
rect 4165 1119 4171 1153
rect 4125 1081 4171 1119
rect 4125 1047 4131 1081
rect 4165 1047 4171 1081
rect 4125 1009 4171 1047
rect 4125 975 4131 1009
rect 4165 975 4171 1009
rect 4125 937 4171 975
rect 4125 903 4131 937
rect 4165 903 4171 937
rect 4125 865 4171 903
tri 4285 1232 4288 1235 se
rect 4288 1232 4334 1263
rect 4451 1873 4497 1885
rect 4451 1839 4457 1873
rect 4491 1839 4497 1873
rect 4451 1801 4497 1839
rect 4451 1767 4457 1801
rect 4491 1767 4497 1801
rect 4451 1729 4497 1767
rect 4451 1695 4457 1729
rect 4491 1695 4497 1729
rect 4451 1657 4497 1695
rect 4451 1623 4457 1657
rect 4491 1623 4497 1657
rect 4451 1585 4497 1623
rect 4451 1551 4457 1585
rect 4491 1551 4497 1585
rect 4451 1513 4497 1551
rect 4451 1479 4457 1513
rect 4491 1479 4497 1513
rect 4451 1441 4497 1479
rect 4451 1407 4457 1441
rect 4491 1407 4497 1441
rect 4451 1369 4497 1407
rect 4451 1335 4457 1369
rect 4491 1335 4497 1369
rect 4451 1297 4497 1335
rect 4451 1263 4457 1297
rect 4491 1263 4497 1297
tri 4334 1232 4337 1235 sw
rect 4285 1226 4337 1232
rect 4285 1157 4337 1174
rect 4285 1088 4337 1105
rect 4285 1019 4337 1036
rect 4285 950 4337 967
rect 4285 892 4337 898
tri 4285 889 4288 892 ne
rect 4125 831 4131 865
rect 4165 831 4171 865
tri 4045 811 4046 812 sw
tri 4124 811 4125 812 se
rect 4125 811 4171 831
rect 4288 865 4334 892
tri 4334 889 4337 892 nw
rect 4451 1225 4497 1263
rect 4614 1873 4660 1885
rect 4614 1839 4620 1873
rect 4654 1839 4660 1873
rect 4614 1801 4660 1839
rect 4614 1767 4620 1801
rect 4654 1767 4660 1801
rect 4614 1729 4660 1767
rect 4614 1695 4620 1729
rect 4654 1695 4660 1729
rect 4614 1657 4660 1695
rect 4614 1623 4620 1657
rect 4654 1623 4660 1657
rect 4614 1585 4660 1623
rect 4614 1551 4620 1585
rect 4654 1551 4660 1585
rect 4614 1513 4660 1551
rect 4614 1479 4620 1513
rect 4654 1479 4660 1513
rect 4614 1441 4660 1479
rect 4614 1407 4620 1441
rect 4654 1407 4660 1441
rect 4614 1369 4660 1407
rect 4614 1335 4620 1369
rect 4654 1335 4660 1369
rect 4614 1297 4660 1335
rect 4614 1263 4620 1297
rect 4654 1263 4660 1297
rect 4451 1191 4457 1225
rect 4491 1191 4497 1225
rect 4451 1153 4497 1191
rect 4451 1119 4457 1153
rect 4491 1119 4497 1153
rect 4451 1081 4497 1119
rect 4451 1047 4457 1081
rect 4491 1047 4497 1081
rect 4451 1009 4497 1047
rect 4451 975 4457 1009
rect 4491 975 4497 1009
rect 4451 937 4497 975
rect 4451 903 4457 937
rect 4491 903 4497 937
rect 4288 831 4294 865
rect 4328 831 4334 865
tri 4171 811 4172 812 sw
rect 4039 809 4046 811
tri 4046 809 4048 811 sw
rect 4039 803 4048 809
rect 3996 739 4048 751
rect 3996 735 4005 739
rect 4039 735 4048 739
rect 3996 666 4048 683
rect 3996 597 4048 614
rect 3996 528 4048 545
rect 3996 470 4048 476
tri 3996 469 3997 470 ne
rect 3997 469 4047 470
tri 4047 469 4048 470 nw
tri 4122 809 4124 811 se
rect 4124 809 4172 811
tri 4172 809 4174 811 sw
rect 4122 803 4174 809
rect 4122 735 4174 751
rect 4122 666 4174 683
rect 4122 597 4174 614
rect 4122 543 4131 545
rect 4165 543 4174 545
rect 4122 528 4174 543
rect 4122 471 4131 476
rect 4165 471 4174 476
rect 4122 470 4174 471
tri 4122 469 4123 470 ne
rect 4123 469 4173 470
tri 4173 469 4174 470 nw
rect 4288 793 4334 831
rect 4451 865 4497 903
tri 4611 1232 4614 1235 se
rect 4614 1232 4660 1263
rect 4777 1873 4823 1885
rect 4777 1839 4783 1873
rect 4817 1839 4823 1873
rect 4777 1801 4823 1839
rect 4777 1767 4783 1801
rect 4817 1767 4823 1801
rect 4777 1729 4823 1767
rect 4777 1695 4783 1729
rect 4817 1695 4823 1729
rect 4777 1657 4823 1695
rect 4777 1623 4783 1657
rect 4817 1623 4823 1657
rect 4777 1585 4823 1623
rect 4777 1551 4783 1585
rect 4817 1551 4823 1585
rect 4777 1513 4823 1551
rect 4777 1479 4783 1513
rect 4817 1479 4823 1513
rect 4777 1441 4823 1479
rect 4777 1407 4783 1441
rect 4817 1407 4823 1441
rect 4777 1369 4823 1407
rect 4777 1335 4783 1369
rect 4817 1335 4823 1369
rect 4777 1297 4823 1335
rect 4777 1263 4783 1297
rect 4817 1263 4823 1297
tri 4660 1232 4663 1235 sw
rect 4611 1226 4663 1232
rect 4611 1157 4663 1174
rect 4611 1088 4663 1105
rect 4611 1019 4663 1036
rect 4611 950 4663 967
rect 4611 892 4663 898
tri 4611 889 4614 892 ne
rect 4451 831 4457 865
rect 4491 831 4497 865
tri 4450 811 4451 812 se
rect 4451 811 4497 831
rect 4614 865 4660 892
tri 4660 889 4663 892 nw
rect 4777 1225 4823 1263
rect 4940 1873 4986 1885
rect 4940 1839 4946 1873
rect 4980 1839 4986 1873
rect 4940 1801 4986 1839
rect 4940 1767 4946 1801
rect 4980 1767 4986 1801
rect 4940 1729 4986 1767
rect 4940 1695 4946 1729
rect 4980 1695 4986 1729
rect 4940 1657 4986 1695
rect 4940 1623 4946 1657
rect 4980 1623 4986 1657
rect 4940 1585 4986 1623
rect 4940 1551 4946 1585
rect 4980 1551 4986 1585
rect 4940 1513 4986 1551
rect 4940 1479 4946 1513
rect 4980 1479 4986 1513
rect 4940 1441 4986 1479
rect 4940 1407 4946 1441
rect 4980 1407 4986 1441
rect 4940 1369 4986 1407
rect 4940 1335 4946 1369
rect 4980 1335 4986 1369
rect 4940 1297 4986 1335
rect 4940 1263 4946 1297
rect 4980 1263 4986 1297
rect 4777 1191 4783 1225
rect 4817 1191 4823 1225
rect 4777 1153 4823 1191
rect 4777 1119 4783 1153
rect 4817 1119 4823 1153
rect 4777 1081 4823 1119
rect 4777 1047 4783 1081
rect 4817 1047 4823 1081
rect 4777 1009 4823 1047
rect 4777 975 4783 1009
rect 4817 975 4823 1009
rect 4777 937 4823 975
rect 4777 903 4783 937
rect 4817 903 4823 937
rect 4614 831 4620 865
rect 4654 831 4660 865
tri 4497 811 4498 812 sw
rect 4288 759 4294 793
rect 4328 759 4334 793
rect 4288 721 4334 759
rect 4288 687 4294 721
rect 4328 687 4334 721
rect 4288 649 4334 687
rect 4288 615 4294 649
rect 4328 615 4334 649
rect 4288 577 4334 615
rect 4288 543 4294 577
rect 4328 543 4334 577
rect 4288 505 4334 543
rect 4288 471 4294 505
rect 4328 471 4334 505
tri 3997 467 3999 469 ne
rect 3750 418 3784 452
rect 3818 418 3852 452
rect 3750 378 3852 418
rect 3750 344 3784 378
rect 3818 344 3852 378
rect 3750 304 3852 344
rect 3999 439 4045 469
tri 4045 467 4047 469 nw
tri 4123 467 4125 469 ne
rect 4125 459 4171 469
tri 4171 467 4173 469 nw
rect 4288 459 4334 471
tri 4448 809 4450 811 se
rect 4450 809 4498 811
tri 4498 809 4500 811 sw
rect 4448 803 4500 809
rect 4448 735 4500 751
rect 4448 666 4500 683
rect 4448 597 4500 614
rect 4448 543 4457 545
rect 4491 543 4500 545
rect 4448 528 4500 543
rect 4448 471 4457 476
rect 4491 471 4500 476
rect 4448 470 4500 471
tri 4448 469 4449 470 ne
rect 4449 469 4499 470
tri 4499 469 4500 470 nw
rect 4614 793 4660 831
rect 4777 865 4823 903
tri 4937 1232 4940 1235 se
rect 4940 1232 4986 1263
rect 5103 1873 5149 1885
rect 5103 1839 5109 1873
rect 5143 1839 5149 1873
rect 5103 1801 5149 1839
rect 5103 1767 5109 1801
rect 5143 1767 5149 1801
rect 5103 1729 5149 1767
rect 5103 1695 5109 1729
rect 5143 1695 5149 1729
rect 5103 1657 5149 1695
rect 5103 1623 5109 1657
rect 5143 1623 5149 1657
rect 5103 1585 5149 1623
rect 5103 1551 5109 1585
rect 5143 1551 5149 1585
rect 5103 1513 5149 1551
rect 5103 1479 5109 1513
rect 5143 1479 5149 1513
rect 5103 1441 5149 1479
rect 5103 1407 5109 1441
rect 5143 1407 5149 1441
rect 5103 1369 5149 1407
rect 5103 1335 5109 1369
rect 5143 1335 5149 1369
rect 5103 1297 5149 1335
rect 5103 1263 5109 1297
rect 5143 1263 5149 1297
tri 4986 1232 4989 1235 sw
rect 4937 1226 4989 1232
rect 4937 1157 4989 1174
rect 4937 1088 4989 1105
rect 4937 1019 4989 1036
rect 4937 950 4989 967
rect 4937 892 4989 898
tri 4937 889 4940 892 ne
rect 4777 831 4783 865
rect 4817 831 4823 865
tri 4776 811 4777 812 se
rect 4777 811 4823 831
rect 4940 865 4986 892
tri 4986 889 4989 892 nw
rect 5103 1225 5149 1263
rect 5266 1873 5312 1885
rect 5266 1839 5272 1873
rect 5306 1839 5312 1873
rect 5266 1801 5312 1839
rect 5266 1767 5272 1801
rect 5306 1767 5312 1801
rect 5266 1729 5312 1767
rect 5266 1695 5272 1729
rect 5306 1695 5312 1729
rect 5389 1873 5435 1885
rect 5389 1839 5395 1873
rect 5429 1839 5435 1873
rect 5389 1801 5435 1839
rect 5389 1767 5395 1801
rect 5429 1767 5435 1801
rect 5389 1729 5435 1767
rect 5266 1657 5312 1695
rect 5266 1623 5272 1657
rect 5306 1623 5312 1657
rect 5266 1585 5312 1623
rect 5266 1551 5272 1585
rect 5306 1551 5312 1585
rect 5266 1513 5312 1551
rect 5266 1479 5272 1513
rect 5306 1479 5312 1513
rect 5266 1441 5312 1479
rect 5266 1407 5272 1441
rect 5306 1407 5312 1441
rect 5266 1369 5312 1407
rect 5266 1335 5272 1369
rect 5306 1335 5312 1369
tri 5386 1723 5389 1726 se
rect 5389 1723 5395 1729
rect 5386 1717 5395 1723
rect 5429 1723 5435 1729
rect 5552 1873 5598 1885
rect 5552 1839 5558 1873
rect 5592 1839 5598 1873
rect 5552 1801 5598 1839
rect 5552 1767 5558 1801
rect 5592 1767 5598 1801
rect 5552 1729 5598 1767
tri 5435 1723 5438 1726 sw
rect 5429 1717 5438 1723
rect 5386 1657 5438 1665
rect 5386 1638 5395 1657
rect 5429 1638 5438 1657
rect 5386 1585 5438 1586
rect 5386 1559 5395 1585
rect 5429 1559 5438 1585
rect 5386 1480 5395 1507
rect 5429 1480 5438 1507
rect 5386 1407 5395 1428
rect 5429 1407 5438 1428
rect 5386 1401 5438 1407
rect 5386 1343 5395 1349
tri 5386 1340 5389 1343 ne
rect 5266 1297 5312 1335
rect 5266 1263 5272 1297
rect 5306 1263 5312 1297
rect 5103 1191 5109 1225
rect 5143 1191 5149 1225
rect 5103 1153 5149 1191
rect 5103 1119 5109 1153
rect 5143 1119 5149 1153
rect 5103 1081 5149 1119
rect 5103 1047 5109 1081
rect 5143 1047 5149 1081
rect 5103 1009 5149 1047
rect 5103 975 5109 1009
rect 5143 975 5149 1009
rect 5103 937 5149 975
rect 5103 903 5109 937
rect 5143 903 5149 937
rect 4940 831 4946 865
rect 4980 831 4986 865
tri 4823 811 4824 812 sw
rect 4614 759 4620 793
rect 4654 759 4660 793
rect 4614 721 4660 759
rect 4614 687 4620 721
rect 4654 687 4660 721
rect 4614 649 4660 687
rect 4614 615 4620 649
rect 4654 615 4660 649
rect 4614 577 4660 615
rect 4614 543 4620 577
rect 4654 543 4660 577
rect 4614 505 4660 543
rect 4614 471 4620 505
rect 4654 471 4660 505
tri 4449 467 4451 469 ne
rect 4451 459 4497 469
tri 4497 467 4499 469 nw
rect 4614 459 4660 471
tri 4774 809 4776 811 se
rect 4776 809 4824 811
tri 4824 809 4826 811 sw
rect 4774 803 4826 809
rect 4774 735 4826 751
rect 4774 666 4826 683
rect 4774 597 4826 614
rect 4774 543 4783 545
rect 4817 543 4826 545
rect 4774 528 4826 543
rect 4774 471 4783 476
rect 4817 471 4826 476
rect 4774 470 4826 471
tri 4774 469 4775 470 ne
rect 4775 469 4825 470
tri 4825 469 4826 470 nw
rect 4940 793 4986 831
rect 5103 865 5149 903
tri 5263 1232 5266 1235 se
rect 5266 1232 5312 1263
rect 5389 1335 5395 1343
rect 5429 1343 5438 1349
rect 5429 1335 5435 1343
tri 5435 1340 5438 1343 nw
rect 5552 1695 5558 1729
rect 5592 1695 5598 1729
rect 5715 1873 5761 1885
rect 5715 1839 5721 1873
rect 5755 1839 5761 1873
rect 5715 1801 5761 1839
rect 5715 1767 5721 1801
rect 5755 1767 5761 1801
rect 5715 1729 5761 1767
rect 5552 1657 5598 1695
rect 5552 1623 5558 1657
rect 5592 1623 5598 1657
rect 5552 1585 5598 1623
rect 5552 1551 5558 1585
rect 5592 1551 5598 1585
rect 5552 1513 5598 1551
rect 5552 1479 5558 1513
rect 5592 1479 5598 1513
rect 5552 1441 5598 1479
rect 5552 1407 5558 1441
rect 5592 1407 5598 1441
rect 5552 1369 5598 1407
rect 5389 1297 5435 1335
rect 5389 1263 5395 1297
rect 5429 1263 5435 1297
tri 5312 1232 5315 1235 sw
rect 5263 1226 5315 1232
rect 5263 1157 5315 1174
rect 5263 1088 5315 1105
rect 5263 1019 5315 1036
rect 5263 950 5315 967
rect 5263 892 5315 898
tri 5263 889 5266 892 ne
rect 5103 831 5109 865
rect 5143 831 5149 865
tri 5102 811 5103 812 se
rect 5103 811 5149 831
rect 5266 865 5312 892
tri 5312 889 5315 892 nw
rect 5389 1225 5435 1263
rect 5389 1191 5395 1225
rect 5429 1191 5435 1225
rect 5389 1153 5435 1191
rect 5389 1119 5395 1153
rect 5429 1119 5435 1153
rect 5389 1081 5435 1119
rect 5389 1047 5395 1081
rect 5429 1047 5435 1081
rect 5389 1009 5435 1047
rect 5389 975 5395 1009
rect 5429 975 5435 1009
rect 5389 937 5435 975
rect 5389 903 5395 937
rect 5429 903 5435 937
rect 5266 831 5272 865
rect 5306 831 5312 865
tri 5149 811 5150 812 sw
rect 4940 759 4946 793
rect 4980 759 4986 793
rect 4940 721 4986 759
rect 4940 687 4946 721
rect 4980 687 4986 721
rect 4940 649 4986 687
rect 4940 615 4946 649
rect 4980 615 4986 649
rect 4940 577 4986 615
rect 4940 543 4946 577
rect 4980 543 4986 577
rect 4940 505 4986 543
rect 4940 471 4946 505
rect 4980 471 4986 505
tri 4775 467 4777 469 ne
rect 4777 459 4823 469
tri 4823 467 4825 469 nw
rect 4940 459 4986 471
tri 5100 809 5102 811 se
rect 5102 809 5150 811
tri 5150 809 5152 811 sw
rect 5100 803 5152 809
rect 5100 735 5152 751
rect 5100 666 5152 683
rect 5100 597 5152 614
rect 5100 543 5109 545
rect 5143 543 5152 545
rect 5100 528 5152 543
rect 5100 471 5109 476
rect 5143 471 5152 476
rect 5100 470 5152 471
tri 5100 469 5101 470 ne
rect 5101 469 5151 470
tri 5151 469 5152 470 nw
rect 5266 793 5312 831
rect 5266 759 5272 793
rect 5306 759 5312 793
rect 5266 721 5312 759
rect 5266 687 5272 721
rect 5306 687 5312 721
rect 5266 649 5312 687
rect 5266 615 5272 649
rect 5306 615 5312 649
rect 5266 577 5312 615
rect 5266 543 5272 577
rect 5306 543 5312 577
rect 5266 505 5312 543
rect 5266 471 5272 505
rect 5306 471 5312 505
tri 5101 467 5103 469 ne
rect 5103 459 5149 469
tri 5149 467 5151 469 nw
rect 5266 459 5312 471
rect 5389 865 5435 903
rect 5389 831 5395 865
rect 5429 831 5435 865
rect 5389 793 5435 831
rect 5552 1335 5558 1369
rect 5592 1335 5598 1369
tri 5712 1723 5715 1726 se
rect 5715 1723 5721 1729
rect 5712 1717 5721 1723
rect 5755 1723 5761 1729
rect 5878 1873 5924 1885
rect 5878 1839 5884 1873
rect 5918 1839 5924 1873
rect 5878 1801 5924 1839
rect 5878 1767 5884 1801
rect 5918 1767 5924 1801
rect 5878 1729 5924 1767
tri 5761 1723 5764 1726 sw
rect 5755 1717 5764 1723
rect 5712 1657 5764 1665
rect 5712 1638 5721 1657
rect 5755 1638 5764 1657
rect 5712 1585 5764 1586
rect 5712 1559 5721 1585
rect 5755 1559 5764 1585
rect 5712 1480 5721 1507
rect 5755 1480 5764 1507
rect 5712 1407 5721 1428
rect 5755 1407 5764 1428
rect 5712 1401 5764 1407
rect 5712 1343 5721 1349
tri 5712 1340 5715 1343 ne
rect 5552 1297 5598 1335
rect 5552 1263 5558 1297
rect 5592 1263 5598 1297
rect 5552 1225 5598 1263
rect 5552 1191 5558 1225
rect 5592 1191 5598 1225
rect 5552 1153 5598 1191
rect 5552 1119 5558 1153
rect 5592 1119 5598 1153
rect 5552 1081 5598 1119
rect 5552 1047 5558 1081
rect 5592 1047 5598 1081
rect 5552 1009 5598 1047
rect 5552 975 5558 1009
rect 5592 975 5598 1009
rect 5552 937 5598 975
rect 5552 903 5558 937
rect 5592 903 5598 937
rect 5552 865 5598 903
rect 5552 831 5558 865
rect 5592 831 5598 865
tri 5551 811 5552 812 se
rect 5552 811 5598 831
rect 5715 1335 5721 1343
rect 5755 1343 5764 1349
rect 5755 1335 5761 1343
tri 5761 1340 5764 1343 nw
rect 5878 1695 5884 1729
rect 5918 1695 5924 1729
rect 6041 1873 6087 1885
rect 6041 1839 6047 1873
rect 6081 1839 6087 1873
rect 6041 1801 6087 1839
rect 6041 1767 6047 1801
rect 6081 1767 6087 1801
rect 6041 1729 6087 1767
rect 5878 1657 5924 1695
rect 5878 1623 5884 1657
rect 5918 1623 5924 1657
rect 5878 1585 5924 1623
rect 5878 1551 5884 1585
rect 5918 1551 5924 1585
rect 5878 1513 5924 1551
rect 5878 1479 5884 1513
rect 5918 1479 5924 1513
rect 5878 1441 5924 1479
rect 5878 1407 5884 1441
rect 5918 1407 5924 1441
rect 5878 1369 5924 1407
rect 5715 1297 5761 1335
rect 5715 1263 5721 1297
rect 5755 1263 5761 1297
rect 5715 1225 5761 1263
rect 5715 1191 5721 1225
rect 5755 1191 5761 1225
rect 5715 1153 5761 1191
rect 5715 1119 5721 1153
rect 5755 1119 5761 1153
rect 5715 1081 5761 1119
rect 5715 1047 5721 1081
rect 5755 1047 5761 1081
rect 5715 1009 5761 1047
rect 5715 975 5721 1009
rect 5755 975 5761 1009
rect 5715 937 5761 975
rect 5715 903 5721 937
rect 5755 903 5761 937
rect 5715 865 5761 903
rect 5715 831 5721 865
rect 5755 831 5761 865
tri 5598 811 5599 812 sw
rect 5389 759 5395 793
rect 5429 759 5435 793
rect 5389 721 5435 759
rect 5389 687 5395 721
rect 5429 687 5435 721
rect 5389 649 5435 687
rect 5389 615 5395 649
rect 5429 615 5435 649
rect 5389 577 5435 615
rect 5389 543 5395 577
rect 5429 543 5435 577
rect 5389 505 5435 543
rect 5389 471 5395 505
rect 5429 471 5435 505
rect 5389 459 5435 471
tri 5549 809 5551 811 se
rect 5551 809 5599 811
tri 5599 809 5601 811 sw
rect 5549 803 5601 809
rect 5549 735 5601 751
rect 5549 666 5601 683
rect 5549 597 5601 614
rect 5549 543 5558 545
rect 5592 543 5601 545
rect 5549 528 5601 543
rect 5549 471 5558 476
rect 5592 471 5601 476
rect 5549 470 5601 471
tri 5549 469 5550 470 ne
rect 5550 469 5600 470
tri 5600 469 5601 470 nw
rect 5715 793 5761 831
rect 5878 1335 5884 1369
rect 5918 1335 5924 1369
tri 6038 1723 6041 1726 se
rect 6041 1723 6047 1729
rect 6038 1717 6047 1723
rect 6081 1723 6087 1729
rect 6204 1873 6250 1885
rect 6204 1839 6210 1873
rect 6244 1839 6250 1873
rect 6204 1801 6250 1839
rect 6204 1767 6210 1801
rect 6244 1767 6250 1801
rect 6204 1729 6250 1767
tri 6087 1723 6090 1726 sw
rect 6081 1717 6090 1723
rect 6038 1657 6090 1665
rect 6038 1638 6047 1657
rect 6081 1638 6090 1657
rect 6038 1585 6090 1586
rect 6038 1559 6047 1585
rect 6081 1559 6090 1585
rect 6038 1480 6047 1507
rect 6081 1480 6090 1507
rect 6038 1407 6047 1428
rect 6081 1407 6090 1428
rect 6038 1401 6090 1407
rect 6038 1343 6047 1349
tri 6038 1340 6041 1343 ne
rect 5878 1297 5924 1335
rect 5878 1263 5884 1297
rect 5918 1263 5924 1297
rect 5878 1225 5924 1263
rect 5878 1191 5884 1225
rect 5918 1191 5924 1225
rect 5878 1153 5924 1191
rect 5878 1119 5884 1153
rect 5918 1119 5924 1153
rect 5878 1081 5924 1119
rect 5878 1047 5884 1081
rect 5918 1047 5924 1081
rect 5878 1009 5924 1047
rect 5878 975 5884 1009
rect 5918 975 5924 1009
rect 5878 937 5924 975
rect 5878 903 5884 937
rect 5918 903 5924 937
rect 5878 865 5924 903
rect 5878 831 5884 865
rect 5918 831 5924 865
tri 5877 811 5878 812 se
rect 5878 811 5924 831
rect 6041 1335 6047 1343
rect 6081 1343 6090 1349
rect 6081 1335 6087 1343
tri 6087 1340 6090 1343 nw
rect 6204 1695 6210 1729
rect 6244 1695 6250 1729
rect 6367 1873 6413 1885
rect 6367 1839 6373 1873
rect 6407 1839 6413 1873
rect 6367 1801 6413 1839
rect 6367 1767 6373 1801
rect 6407 1767 6413 1801
rect 6367 1729 6413 1767
rect 6204 1657 6250 1695
rect 6204 1623 6210 1657
rect 6244 1623 6250 1657
rect 6204 1585 6250 1623
rect 6204 1551 6210 1585
rect 6244 1551 6250 1585
rect 6204 1513 6250 1551
rect 6204 1479 6210 1513
rect 6244 1479 6250 1513
rect 6204 1441 6250 1479
rect 6204 1407 6210 1441
rect 6244 1407 6250 1441
rect 6204 1369 6250 1407
rect 6041 1297 6087 1335
rect 6041 1263 6047 1297
rect 6081 1263 6087 1297
rect 6041 1225 6087 1263
rect 6041 1191 6047 1225
rect 6081 1191 6087 1225
rect 6041 1153 6087 1191
rect 6041 1119 6047 1153
rect 6081 1119 6087 1153
rect 6041 1081 6087 1119
rect 6041 1047 6047 1081
rect 6081 1047 6087 1081
rect 6041 1009 6087 1047
rect 6041 975 6047 1009
rect 6081 975 6087 1009
rect 6041 937 6087 975
rect 6041 903 6047 937
rect 6081 903 6087 937
rect 6041 865 6087 903
rect 6041 831 6047 865
rect 6081 831 6087 865
tri 5924 811 5925 812 sw
rect 5715 759 5721 793
rect 5755 759 5761 793
rect 5715 721 5761 759
rect 5715 687 5721 721
rect 5755 687 5761 721
rect 5715 649 5761 687
rect 5715 615 5721 649
rect 5755 615 5761 649
rect 5715 577 5761 615
rect 5715 543 5721 577
rect 5755 543 5761 577
rect 5715 505 5761 543
rect 5715 471 5721 505
rect 5755 471 5761 505
tri 5550 467 5552 469 ne
rect 5552 459 5598 469
tri 5598 467 5600 469 nw
rect 5715 459 5761 471
tri 5875 809 5877 811 se
rect 5877 809 5925 811
tri 5925 809 5927 811 sw
rect 5875 803 5927 809
rect 5875 735 5927 751
rect 5875 666 5927 683
rect 5875 597 5927 614
rect 5875 543 5884 545
rect 5918 543 5927 545
rect 5875 528 5927 543
rect 5875 471 5884 476
rect 5918 471 5927 476
rect 5875 470 5927 471
tri 5875 469 5876 470 ne
rect 5876 469 5926 470
tri 5926 469 5927 470 nw
rect 6041 793 6087 831
rect 6204 1335 6210 1369
rect 6244 1335 6250 1369
tri 6364 1723 6367 1726 se
rect 6367 1723 6373 1729
rect 6364 1717 6373 1723
rect 6407 1723 6413 1729
rect 6530 1873 6576 1885
rect 6530 1839 6536 1873
rect 6570 1839 6576 1873
rect 6530 1801 6576 1839
rect 6530 1767 6536 1801
rect 6570 1767 6576 1801
rect 6530 1729 6576 1767
tri 6413 1723 6416 1726 sw
rect 6407 1717 6416 1723
rect 6364 1657 6416 1665
rect 6364 1638 6373 1657
rect 6407 1638 6416 1657
rect 6364 1585 6416 1586
rect 6364 1559 6373 1585
rect 6407 1559 6416 1585
rect 6364 1480 6373 1507
rect 6407 1480 6416 1507
rect 6364 1407 6373 1428
rect 6407 1407 6416 1428
rect 6364 1401 6416 1407
rect 6364 1343 6373 1349
tri 6364 1340 6367 1343 ne
rect 6204 1297 6250 1335
rect 6204 1263 6210 1297
rect 6244 1263 6250 1297
rect 6204 1225 6250 1263
rect 6204 1191 6210 1225
rect 6244 1191 6250 1225
rect 6204 1153 6250 1191
rect 6204 1119 6210 1153
rect 6244 1119 6250 1153
rect 6204 1081 6250 1119
rect 6204 1047 6210 1081
rect 6244 1047 6250 1081
rect 6204 1009 6250 1047
rect 6204 975 6210 1009
rect 6244 975 6250 1009
rect 6204 937 6250 975
rect 6204 903 6210 937
rect 6244 903 6250 937
rect 6204 865 6250 903
rect 6204 831 6210 865
rect 6244 831 6250 865
tri 6203 811 6204 812 se
rect 6204 811 6250 831
rect 6367 1335 6373 1343
rect 6407 1343 6416 1349
rect 6407 1335 6413 1343
tri 6413 1340 6416 1343 nw
rect 6530 1695 6536 1729
rect 6570 1695 6576 1729
rect 6530 1657 6576 1695
rect 6530 1623 6536 1657
rect 6570 1623 6576 1657
rect 6530 1585 6576 1623
rect 6530 1551 6536 1585
rect 6570 1551 6576 1585
rect 6530 1513 6576 1551
rect 6530 1479 6536 1513
rect 6570 1479 6576 1513
rect 6530 1441 6576 1479
rect 6530 1407 6536 1441
rect 6570 1407 6576 1441
rect 6530 1369 6576 1407
rect 6367 1297 6413 1335
rect 6367 1263 6373 1297
rect 6407 1263 6413 1297
rect 6367 1225 6413 1263
rect 6367 1191 6373 1225
rect 6407 1191 6413 1225
rect 6367 1153 6413 1191
rect 6367 1119 6373 1153
rect 6407 1119 6413 1153
rect 6367 1081 6413 1119
rect 6367 1047 6373 1081
rect 6407 1047 6413 1081
rect 6367 1009 6413 1047
rect 6367 975 6373 1009
rect 6407 975 6413 1009
rect 6367 937 6413 975
rect 6367 903 6373 937
rect 6407 903 6413 937
rect 6367 865 6413 903
rect 6367 831 6373 865
rect 6407 831 6413 865
tri 6250 811 6251 812 sw
rect 6041 759 6047 793
rect 6081 759 6087 793
rect 6041 721 6087 759
rect 6041 687 6047 721
rect 6081 687 6087 721
rect 6041 649 6087 687
rect 6041 615 6047 649
rect 6081 615 6087 649
rect 6041 577 6087 615
rect 6041 543 6047 577
rect 6081 543 6087 577
rect 6041 505 6087 543
rect 6041 471 6047 505
rect 6081 471 6087 505
tri 5876 467 5878 469 ne
rect 5878 459 5924 469
tri 5924 467 5926 469 nw
rect 6041 459 6087 471
tri 6201 809 6203 811 se
rect 6203 809 6251 811
tri 6251 809 6253 811 sw
rect 6201 803 6253 809
rect 6201 735 6253 751
rect 6201 666 6253 683
rect 6201 597 6253 614
rect 6201 543 6210 545
rect 6244 543 6253 545
rect 6201 528 6253 543
rect 6201 471 6210 476
rect 6244 471 6253 476
rect 6201 470 6253 471
tri 6201 469 6202 470 ne
rect 6202 469 6252 470
tri 6252 469 6253 470 nw
rect 6367 793 6413 831
rect 6530 1335 6536 1369
rect 6570 1335 6576 1369
rect 6530 1297 6576 1335
rect 6530 1263 6536 1297
rect 6570 1263 6576 1297
rect 6530 1225 6576 1263
rect 6530 1191 6536 1225
rect 6570 1191 6576 1225
rect 6530 1153 6576 1191
rect 6530 1119 6536 1153
rect 6570 1119 6576 1153
rect 6530 1081 6576 1119
rect 6530 1047 6536 1081
rect 6570 1047 6576 1081
rect 6530 1009 6576 1047
rect 6530 975 6536 1009
rect 6570 975 6576 1009
rect 6530 937 6576 975
rect 6530 903 6536 937
rect 6570 903 6576 937
rect 6530 865 6576 903
rect 6530 831 6536 865
rect 6570 831 6576 865
tri 6529 811 6530 812 se
rect 6530 811 6576 831
rect 6649 1851 6695 1892
rect 6649 1817 6655 1851
rect 6689 1817 6695 1851
rect 6649 1776 6695 1817
rect 6649 1742 6655 1776
rect 6689 1742 6695 1776
rect 6649 1701 6695 1742
rect 6649 1667 6655 1701
rect 6689 1667 6695 1701
rect 6649 1626 6695 1667
rect 6649 1592 6655 1626
rect 6689 1592 6695 1626
rect 6649 1551 6695 1592
rect 6649 1517 6655 1551
rect 6689 1517 6695 1551
rect 6649 1477 6695 1517
rect 6649 1443 6655 1477
rect 6689 1443 6695 1477
rect 6649 1403 6695 1443
rect 6649 1369 6655 1403
rect 6689 1369 6695 1403
rect 6649 1329 6695 1369
rect 6649 1295 6655 1329
rect 6689 1295 6695 1329
rect 6649 1255 6695 1295
rect 6649 1221 6655 1255
rect 6689 1221 6695 1255
rect 6649 1181 6695 1221
rect 6649 1147 6655 1181
rect 6689 1147 6695 1181
rect 6649 1107 6695 1147
rect 6649 1073 6655 1107
rect 6689 1073 6695 1107
rect 6649 1033 6695 1073
rect 6649 999 6655 1033
rect 6689 999 6695 1033
rect 6649 959 6695 999
rect 6649 925 6655 959
rect 6689 925 6695 959
rect 6649 885 6695 925
rect 6649 851 6655 885
rect 6689 851 6695 885
tri 6576 811 6577 812 sw
tri 6648 811 6649 812 se
rect 6649 811 6695 851
rect 6842 2062 6944 2102
rect 6842 2028 6876 2062
rect 6910 2028 6944 2062
rect 6842 1988 6944 2028
rect 6842 1954 6876 1988
rect 6910 1954 6944 1988
rect 6842 1914 6944 1954
rect 6842 1880 6876 1914
rect 6910 1880 6944 1914
rect 6842 1840 6944 1880
rect 6842 1806 6876 1840
rect 6910 1806 6944 1840
rect 6842 1766 6944 1806
rect 6842 1732 6876 1766
rect 6910 1732 6944 1766
rect 7091 2107 10003 2113
rect 7091 2073 7170 2107
rect 7204 2073 7243 2107
rect 7277 2073 7316 2107
rect 7350 2073 7389 2107
rect 7423 2073 7463 2107
rect 7497 2073 7537 2107
rect 7571 2073 7611 2107
rect 7645 2073 7685 2107
rect 7719 2073 7759 2107
rect 7793 2073 7833 2107
rect 7867 2073 7907 2107
rect 7941 2073 7981 2107
rect 8015 2073 8055 2107
rect 8089 2073 8129 2107
rect 8163 2073 8203 2107
rect 8237 2073 8277 2107
rect 8311 2073 8351 2107
rect 8385 2073 8425 2107
rect 8459 2073 8499 2107
rect 8533 2073 8573 2107
rect 8607 2073 8647 2107
rect 8681 2073 8721 2107
rect 8755 2073 8795 2107
rect 8829 2073 8869 2107
rect 8903 2073 8943 2107
rect 8977 2073 9017 2107
rect 9051 2073 9091 2107
rect 9125 2073 9165 2107
rect 9199 2073 9239 2107
rect 9273 2073 9313 2107
rect 9347 2073 9387 2107
rect 9421 2073 9461 2107
rect 9495 2073 9535 2107
rect 9569 2073 9645 2107
rect 9679 2073 9727 2107
rect 9761 2073 9809 2107
rect 9843 2073 9891 2107
rect 9925 2073 10003 2107
rect 7091 2067 10003 2073
rect 7091 2035 7138 2067
rect 7091 2001 7097 2035
rect 7131 2034 7138 2035
tri 7138 2034 7171 2067 nw
tri 9923 2034 9956 2067 ne
rect 9956 2034 10003 2067
rect 7131 2001 7137 2034
tri 7137 2033 7138 2034 nw
rect 7091 1960 7137 2001
rect 7261 2025 7286 2034
rect 7338 2025 7351 2034
rect 7261 1991 7273 2025
rect 7338 1991 7346 2025
rect 7261 1982 7286 1991
rect 7338 1982 7351 1991
rect 7403 1982 7416 2034
rect 7468 1982 7481 2034
rect 7533 1982 7546 2034
rect 7598 2025 7611 2034
rect 7663 2025 7676 2034
rect 7728 2025 8195 2034
rect 7599 1991 7611 2025
rect 7672 1991 7676 2025
rect 7745 1991 7784 2025
rect 7818 1991 7857 2025
rect 7891 1991 7930 2025
rect 7964 1991 8003 2025
rect 8037 1991 8075 2025
rect 8109 1991 8147 2025
rect 8181 1991 8195 2025
rect 7598 1982 7611 1991
rect 7663 1982 7676 1991
rect 7728 1982 8195 1991
rect 8242 1982 8248 2034
rect 8300 1982 8312 2034
rect 8364 2025 9778 2034
tri 9956 2033 9957 2034 ne
rect 9957 2033 10003 2034
rect 8364 1991 8544 2025
rect 8578 1991 8619 2025
rect 8653 1991 8694 2025
rect 8728 1991 8769 2025
rect 8803 1991 8844 2025
rect 8878 1991 8918 2025
rect 8952 1991 8992 2025
rect 9026 1991 9066 2025
rect 9100 1991 9140 2025
rect 9174 1991 9214 2025
rect 9248 1991 9288 2025
rect 9322 1991 9362 2025
rect 9396 1991 9436 2025
rect 9470 1991 9510 2025
rect 9544 1991 9584 2025
rect 9618 1991 9658 2025
rect 9692 1991 9732 2025
rect 9766 1991 9778 2025
rect 8364 1982 9778 1991
rect 9957 1999 9963 2033
rect 9997 1999 10003 2033
rect 7091 1926 7097 1960
rect 7131 1926 7137 1960
rect 9957 1959 10003 1999
rect 7091 1885 7137 1926
rect 7091 1851 7097 1885
rect 7131 1851 7137 1885
rect 7091 1810 7137 1851
rect 7091 1776 7097 1810
rect 7131 1776 7137 1810
rect 6842 1692 6944 1732
rect 6842 1658 6876 1692
rect 6910 1658 6944 1692
rect 6842 1618 6944 1658
rect 6842 1584 6876 1618
rect 6910 1584 6944 1618
rect 6842 1544 6944 1584
rect 6842 1510 6876 1544
rect 6910 1510 6944 1544
rect 6842 1471 6944 1510
rect 6842 1437 6876 1471
rect 6910 1437 6944 1471
rect 6842 1398 6944 1437
rect 6842 1364 6876 1398
rect 6910 1364 6944 1398
tri 7088 1738 7091 1741 se
rect 7091 1738 7137 1776
rect 7210 1941 7256 1953
rect 7210 1907 7216 1941
rect 7250 1907 7256 1941
rect 7210 1869 7256 1907
rect 7210 1835 7216 1869
rect 7250 1835 7256 1869
rect 7210 1797 7256 1835
rect 7210 1763 7216 1797
rect 7250 1763 7256 1797
tri 7137 1738 7140 1741 sw
rect 7088 1735 7140 1738
rect 7088 1732 7097 1735
rect 7131 1732 7140 1735
rect 7088 1661 7140 1680
rect 7088 1590 7140 1609
rect 7088 1518 7140 1538
rect 7088 1446 7140 1466
rect 7088 1388 7140 1394
tri 7088 1386 7090 1388 ne
rect 7090 1386 7138 1388
tri 7138 1386 7140 1388 nw
rect 7210 1725 7256 1763
rect 7373 1941 7419 1953
rect 7373 1907 7379 1941
rect 7413 1907 7419 1941
rect 7373 1869 7419 1907
rect 7373 1835 7379 1869
rect 7413 1835 7419 1869
rect 7373 1797 7419 1835
rect 7373 1763 7379 1797
rect 7413 1763 7419 1797
rect 7210 1691 7216 1725
rect 7250 1691 7256 1725
rect 7210 1653 7256 1691
rect 7210 1619 7216 1653
rect 7250 1619 7256 1653
rect 7210 1581 7256 1619
rect 7210 1547 7216 1581
rect 7250 1547 7256 1581
rect 7210 1509 7256 1547
rect 7210 1475 7216 1509
rect 7250 1475 7256 1509
rect 7210 1437 7256 1475
rect 7210 1403 7216 1437
rect 7250 1403 7256 1437
tri 7090 1385 7091 1386 ne
rect 6842 1325 6944 1364
rect 6842 1291 6876 1325
rect 6910 1291 6944 1325
rect 6842 1252 6944 1291
rect 6842 1218 6876 1252
rect 6910 1218 6944 1252
rect 6842 1179 6944 1218
rect 6842 1145 6876 1179
rect 6910 1145 6944 1179
rect 6842 1106 6944 1145
rect 6842 1072 6876 1106
rect 6910 1072 6944 1106
rect 6842 1033 6944 1072
rect 6842 999 6876 1033
rect 6910 999 6944 1033
rect 6842 960 6944 999
rect 6842 926 6876 960
rect 6910 926 6944 960
rect 6842 887 6944 926
rect 6842 853 6876 887
rect 6910 853 6944 887
rect 6842 814 6944 853
rect 6367 759 6373 793
rect 6407 759 6413 793
rect 6367 721 6413 759
rect 6367 687 6373 721
rect 6407 687 6413 721
rect 6367 649 6413 687
rect 6367 615 6373 649
rect 6407 615 6413 649
rect 6367 577 6413 615
rect 6367 543 6373 577
rect 6407 543 6413 577
rect 6367 505 6413 543
rect 6367 471 6373 505
rect 6407 471 6413 505
tri 6202 467 6204 469 ne
rect 6204 459 6250 469
tri 6250 467 6252 469 nw
rect 6367 459 6413 471
tri 6527 809 6529 811 se
rect 6529 809 6577 811
tri 6577 809 6579 811 sw
rect 6527 803 6579 809
rect 6527 735 6579 751
rect 6527 666 6579 683
rect 6527 597 6579 614
rect 6527 543 6536 545
rect 6570 543 6579 545
rect 6527 528 6579 543
rect 6527 471 6536 476
rect 6570 471 6579 476
rect 6527 470 6579 471
tri 6527 469 6528 470 ne
rect 6528 469 6578 470
tri 6578 469 6579 470 nw
tri 6646 809 6648 811 se
rect 6648 809 6655 811
rect 6646 803 6655 809
rect 6689 809 6695 811
tri 6695 809 6698 812 sw
rect 6689 803 6698 809
rect 6646 737 6698 751
rect 6646 735 6655 737
rect 6689 735 6698 737
rect 6646 666 6698 683
rect 6646 597 6698 614
rect 6646 528 6698 545
rect 6646 470 6698 476
tri 6646 469 6647 470 ne
rect 6647 469 6697 470
tri 6697 469 6698 470 nw
rect 6842 780 6876 814
rect 6910 780 6944 814
rect 6842 741 6944 780
rect 6842 707 6876 741
rect 6910 707 6944 741
rect 6842 668 6944 707
rect 6842 634 6876 668
rect 6910 634 6944 668
rect 6842 595 6944 634
rect 6842 561 6876 595
rect 6910 561 6944 595
rect 6842 522 6944 561
rect 6842 488 6876 522
rect 6910 488 6944 522
tri 6528 467 6530 469 ne
rect 6530 459 6576 469
tri 6576 467 6578 469 nw
tri 6647 467 6649 469 ne
rect 3999 405 4005 439
rect 4039 405 4045 439
rect 6649 441 6695 469
tri 6695 467 6697 469 nw
rect 6649 407 6655 441
rect 6689 407 6695 441
rect 3999 404 4045 405
tri 4045 404 4048 407 sw
tri 6646 404 6649 407 se
rect 6649 404 6695 407
rect 3999 376 4048 404
tri 4048 376 4076 404 sw
tri 6618 376 6646 404 se
rect 6646 376 6695 404
rect 3999 373 4076 376
tri 4076 373 4079 376 sw
tri 6615 373 6618 376 se
rect 6618 373 6695 376
rect 3999 367 6695 373
rect 3999 333 4078 367
rect 4112 333 4151 367
rect 4185 333 4224 367
rect 4258 333 4297 367
rect 4331 333 4370 367
rect 4404 333 4443 367
rect 4477 333 4516 367
rect 4550 333 4589 367
rect 4623 333 4662 367
rect 4696 333 4735 367
rect 4769 333 4808 367
rect 4842 333 4881 367
rect 4915 333 4955 367
rect 4989 333 5029 367
rect 5063 333 5103 367
rect 5137 333 5177 367
rect 5211 333 5251 367
rect 5285 333 5325 367
rect 5359 333 5399 367
rect 5433 333 5473 367
rect 5507 333 5547 367
rect 5581 333 5621 367
rect 5655 333 5695 367
rect 5729 333 5769 367
rect 5803 333 5843 367
rect 5877 333 5917 367
rect 5951 333 5991 367
rect 6025 333 6065 367
rect 6099 333 6139 367
rect 6173 333 6213 367
rect 6247 333 6287 367
rect 6321 333 6361 367
rect 6395 333 6435 367
rect 6469 333 6509 367
rect 6543 333 6583 367
rect 6617 333 6695 367
rect 3999 327 6695 333
rect 6842 449 6944 488
rect 6842 415 6876 449
rect 6910 415 6944 449
rect 7091 1360 7137 1386
tri 7137 1385 7138 1386 nw
rect 7091 1326 7097 1360
rect 7131 1326 7137 1360
rect 7091 1285 7137 1326
rect 7091 1251 7097 1285
rect 7131 1251 7137 1285
rect 7091 1210 7137 1251
rect 7210 1365 7256 1403
tri 7370 1738 7373 1741 se
rect 7373 1738 7419 1763
rect 7536 1941 7582 1953
rect 7536 1907 7542 1941
rect 7576 1907 7582 1941
rect 7536 1869 7582 1907
rect 7536 1835 7542 1869
rect 7576 1835 7582 1869
rect 7536 1797 7582 1835
rect 7536 1763 7542 1797
rect 7576 1763 7582 1797
tri 7419 1738 7422 1741 sw
rect 7370 1732 7422 1738
rect 7370 1661 7422 1680
rect 7370 1590 7422 1609
rect 7370 1518 7422 1538
rect 7370 1446 7422 1466
rect 7370 1388 7422 1394
tri 7370 1386 7372 1388 ne
rect 7372 1386 7420 1388
tri 7420 1386 7422 1388 nw
rect 7536 1725 7582 1763
rect 7699 1941 7745 1953
rect 7699 1907 7705 1941
rect 7739 1907 7745 1941
rect 7699 1869 7745 1907
rect 7699 1835 7705 1869
rect 7739 1835 7745 1869
rect 7699 1797 7745 1835
rect 7699 1763 7705 1797
rect 7739 1763 7745 1797
rect 7536 1691 7542 1725
rect 7576 1691 7582 1725
rect 7536 1653 7582 1691
rect 7536 1619 7542 1653
rect 7576 1619 7582 1653
rect 7536 1581 7582 1619
rect 7536 1547 7542 1581
rect 7576 1547 7582 1581
rect 7536 1509 7582 1547
rect 7536 1475 7542 1509
rect 7576 1475 7582 1509
rect 7536 1437 7582 1475
rect 7536 1403 7542 1437
rect 7576 1403 7582 1437
tri 7372 1385 7373 1386 ne
rect 7210 1331 7216 1365
rect 7250 1331 7256 1365
rect 7210 1293 7256 1331
rect 7210 1259 7216 1293
rect 7250 1259 7256 1293
rect 7091 1176 7097 1210
rect 7131 1176 7137 1210
rect 7091 1135 7137 1176
rect 7091 1101 7097 1135
rect 7131 1101 7137 1135
rect 7091 1061 7137 1101
rect 7091 1027 7097 1061
rect 7131 1027 7137 1061
rect 7091 987 7137 1027
rect 7091 953 7097 987
rect 7131 953 7137 987
rect 7091 913 7137 953
rect 7091 879 7097 913
rect 7131 879 7137 913
tri 7207 1232 7210 1235 se
rect 7210 1232 7256 1259
rect 7373 1365 7419 1386
tri 7419 1385 7420 1386 nw
rect 7373 1331 7379 1365
rect 7413 1331 7419 1365
rect 7373 1293 7419 1331
rect 7373 1259 7379 1293
rect 7413 1259 7419 1293
tri 7256 1232 7259 1235 sw
rect 7207 1226 7259 1232
rect 7207 1157 7259 1174
rect 7207 1088 7259 1105
rect 7207 1019 7259 1036
rect 7207 950 7259 967
rect 7207 892 7259 898
tri 7207 889 7210 892 ne
rect 7091 839 7137 879
rect 7091 805 7097 839
rect 7131 805 7137 839
rect 7091 765 7137 805
rect 7091 731 7097 765
rect 7131 731 7137 765
rect 7091 691 7137 731
rect 7091 657 7097 691
rect 7131 657 7137 691
rect 7091 617 7137 657
rect 7091 583 7097 617
rect 7131 583 7137 617
rect 7091 543 7137 583
rect 7091 509 7097 543
rect 7131 509 7137 543
rect 7210 861 7256 892
tri 7256 889 7259 892 nw
rect 7373 1221 7419 1259
rect 7536 1365 7582 1403
tri 7696 1738 7699 1741 se
rect 7699 1738 7745 1763
rect 7862 1941 7908 1953
rect 7862 1907 7868 1941
rect 7902 1907 7908 1941
rect 7862 1869 7908 1907
rect 7862 1835 7868 1869
rect 7902 1835 7908 1869
rect 7862 1797 7908 1835
rect 7862 1763 7868 1797
rect 7902 1763 7908 1797
tri 7745 1738 7748 1741 sw
rect 7696 1732 7748 1738
rect 7696 1661 7748 1680
rect 7696 1590 7748 1609
rect 7696 1518 7748 1538
rect 7696 1446 7748 1466
rect 7696 1388 7748 1394
tri 7696 1386 7698 1388 ne
rect 7698 1386 7746 1388
tri 7746 1386 7748 1388 nw
rect 7862 1725 7908 1763
rect 8025 1941 8071 1953
rect 8025 1907 8031 1941
rect 8065 1907 8071 1941
rect 8025 1869 8071 1907
rect 8025 1835 8031 1869
rect 8065 1835 8071 1869
rect 8025 1797 8071 1835
rect 8025 1763 8031 1797
rect 8065 1763 8071 1797
rect 7862 1691 7868 1725
rect 7902 1691 7908 1725
rect 7862 1653 7908 1691
rect 7862 1619 7868 1653
rect 7902 1619 7908 1653
rect 7862 1581 7908 1619
rect 7862 1547 7868 1581
rect 7902 1547 7908 1581
rect 7862 1509 7908 1547
rect 7862 1475 7868 1509
rect 7902 1475 7908 1509
rect 7862 1437 7908 1475
rect 7862 1403 7868 1437
rect 7902 1403 7908 1437
tri 7698 1385 7699 1386 ne
rect 7536 1331 7542 1365
rect 7576 1331 7582 1365
rect 7536 1293 7582 1331
rect 7536 1259 7542 1293
rect 7576 1259 7582 1293
rect 7373 1187 7379 1221
rect 7413 1187 7419 1221
rect 7373 1149 7419 1187
rect 7373 1115 7379 1149
rect 7413 1115 7419 1149
rect 7373 1077 7419 1115
rect 7373 1043 7379 1077
rect 7413 1043 7419 1077
rect 7373 1005 7419 1043
rect 7373 971 7379 1005
rect 7413 971 7419 1005
rect 7373 933 7419 971
rect 7373 899 7379 933
rect 7413 899 7419 933
rect 7210 827 7216 861
rect 7250 827 7256 861
rect 7210 789 7256 827
rect 7210 755 7216 789
rect 7250 755 7256 789
rect 7210 717 7256 755
rect 7210 683 7216 717
rect 7250 683 7256 717
rect 7210 645 7256 683
rect 7210 611 7216 645
rect 7250 611 7256 645
rect 7210 573 7256 611
rect 7210 539 7216 573
rect 7250 539 7256 573
rect 7210 527 7256 539
rect 7373 861 7419 899
tri 7533 1232 7536 1235 se
rect 7536 1232 7582 1259
rect 7699 1365 7745 1386
tri 7745 1385 7746 1386 nw
rect 7699 1331 7705 1365
rect 7739 1331 7745 1365
rect 7699 1293 7745 1331
rect 7699 1259 7705 1293
rect 7739 1259 7745 1293
tri 7582 1232 7585 1235 sw
rect 7533 1226 7585 1232
rect 7533 1157 7585 1174
rect 7533 1088 7585 1105
rect 7533 1019 7585 1036
rect 7533 950 7585 967
rect 7533 892 7585 898
tri 7533 889 7536 892 ne
rect 7373 827 7379 861
rect 7413 827 7419 861
rect 7373 789 7419 827
rect 7373 755 7379 789
rect 7413 755 7419 789
rect 7373 717 7419 755
rect 7373 683 7379 717
rect 7413 683 7419 717
rect 7373 645 7419 683
rect 7373 611 7379 645
rect 7413 611 7419 645
rect 7373 573 7419 611
rect 7373 539 7379 573
rect 7413 539 7419 573
rect 7373 527 7419 539
rect 7536 861 7582 892
tri 7582 889 7585 892 nw
rect 7699 1221 7745 1259
rect 7862 1365 7908 1403
tri 8022 1738 8025 1741 se
rect 8025 1738 8071 1763
rect 8188 1941 8234 1953
rect 8188 1907 8194 1941
rect 8228 1907 8234 1941
rect 8188 1869 8234 1907
rect 8188 1835 8194 1869
rect 8228 1835 8234 1869
rect 8188 1797 8234 1835
rect 8188 1763 8194 1797
rect 8228 1763 8234 1797
tri 8071 1738 8074 1741 sw
rect 8022 1732 8074 1738
rect 8022 1661 8074 1680
rect 8022 1590 8074 1609
rect 8022 1518 8074 1538
rect 8022 1446 8074 1466
rect 8022 1388 8074 1394
tri 8022 1386 8024 1388 ne
rect 8024 1386 8072 1388
tri 8072 1386 8074 1388 nw
rect 8188 1725 8234 1763
rect 8188 1691 8194 1725
rect 8228 1691 8234 1725
rect 8188 1653 8234 1691
rect 8188 1619 8194 1653
rect 8228 1619 8234 1653
rect 8188 1581 8234 1619
rect 8188 1547 8194 1581
rect 8228 1547 8234 1581
rect 8188 1509 8234 1547
rect 8188 1475 8194 1509
rect 8228 1475 8234 1509
rect 8188 1437 8234 1475
rect 8188 1403 8194 1437
rect 8228 1403 8234 1437
tri 8024 1385 8025 1386 ne
rect 7862 1331 7868 1365
rect 7902 1331 7908 1365
rect 7862 1293 7908 1331
rect 7862 1259 7868 1293
rect 7902 1259 7908 1293
rect 7699 1187 7705 1221
rect 7739 1187 7745 1221
rect 7699 1149 7745 1187
rect 7699 1115 7705 1149
rect 7739 1115 7745 1149
rect 7699 1077 7745 1115
rect 7699 1043 7705 1077
rect 7739 1043 7745 1077
rect 7699 1005 7745 1043
rect 7699 971 7705 1005
rect 7739 971 7745 1005
rect 7699 933 7745 971
rect 7699 899 7705 933
rect 7739 899 7745 933
rect 7536 827 7542 861
rect 7576 827 7582 861
rect 7536 789 7582 827
rect 7536 755 7542 789
rect 7576 755 7582 789
rect 7536 717 7582 755
rect 7536 683 7542 717
rect 7576 683 7582 717
rect 7536 645 7582 683
rect 7536 611 7542 645
rect 7576 611 7582 645
rect 7536 573 7582 611
rect 7536 539 7542 573
rect 7576 539 7582 573
rect 7536 527 7582 539
rect 7699 861 7745 899
tri 7859 1232 7862 1235 se
rect 7862 1232 7908 1259
rect 8025 1365 8071 1386
tri 8071 1385 8072 1386 nw
rect 8025 1331 8031 1365
rect 8065 1331 8071 1365
rect 8025 1293 8071 1331
rect 8025 1259 8031 1293
rect 8065 1259 8071 1293
tri 7908 1232 7911 1235 sw
rect 7859 1226 7911 1232
rect 7859 1157 7911 1174
rect 7859 1088 7911 1105
rect 7859 1019 7911 1036
rect 7859 950 7911 967
rect 7859 892 7911 898
tri 7859 889 7862 892 ne
rect 7699 827 7705 861
rect 7739 827 7745 861
rect 7699 789 7745 827
rect 7699 755 7705 789
rect 7739 755 7745 789
rect 7699 717 7745 755
rect 7699 683 7705 717
rect 7739 683 7745 717
rect 7699 645 7745 683
rect 7699 611 7705 645
rect 7739 611 7745 645
rect 7699 573 7745 611
rect 7699 539 7705 573
rect 7739 539 7745 573
rect 7699 527 7745 539
rect 7862 861 7908 892
tri 7908 889 7911 892 nw
rect 8025 1221 8071 1259
rect 8188 1365 8234 1403
rect 8188 1331 8194 1365
rect 8228 1331 8234 1365
rect 8188 1293 8234 1331
rect 8188 1259 8194 1293
rect 8228 1259 8234 1293
rect 8025 1187 8031 1221
rect 8065 1187 8071 1221
rect 8025 1149 8071 1187
rect 8025 1115 8031 1149
rect 8065 1115 8071 1149
rect 8025 1077 8071 1115
rect 8025 1043 8031 1077
rect 8065 1043 8071 1077
rect 8025 1005 8071 1043
rect 8025 971 8031 1005
rect 8065 971 8071 1005
rect 8025 933 8071 971
rect 8025 899 8031 933
rect 8065 899 8071 933
rect 7862 827 7868 861
rect 7902 827 7908 861
rect 7862 789 7908 827
rect 7862 755 7868 789
rect 7902 755 7908 789
rect 7862 717 7908 755
rect 7862 683 7868 717
rect 7902 683 7908 717
rect 7862 645 7908 683
rect 7862 611 7868 645
rect 7902 611 7908 645
rect 7862 573 7908 611
rect 7862 539 7868 573
rect 7902 539 7908 573
rect 7862 527 7908 539
rect 8025 861 8071 899
tri 8185 1232 8188 1235 se
rect 8188 1232 8234 1259
rect 8351 1941 8520 1953
rect 8351 1907 8357 1941
rect 8391 1907 8520 1941
rect 9957 1925 9963 1959
rect 9997 1925 10003 1959
rect 8351 1899 8520 1907
rect 8351 1869 8480 1899
rect 8351 1835 8357 1869
rect 8391 1865 8480 1869
rect 8514 1865 8520 1899
rect 8391 1835 8520 1865
rect 8351 1824 8520 1835
rect 8351 1797 8480 1824
rect 8351 1763 8357 1797
rect 8391 1790 8480 1797
rect 8514 1790 8520 1824
rect 8391 1763 8520 1790
rect 8351 1749 8520 1763
rect 8351 1725 8480 1749
rect 8351 1691 8357 1725
rect 8391 1715 8480 1725
rect 8514 1715 8520 1749
rect 8391 1691 8520 1715
rect 8351 1674 8520 1691
rect 8351 1653 8480 1674
rect 8351 1619 8357 1653
rect 8391 1640 8480 1653
rect 8514 1640 8520 1674
rect 8391 1619 8520 1640
rect 8351 1599 8520 1619
rect 8351 1581 8480 1599
rect 8351 1547 8357 1581
rect 8391 1565 8480 1581
rect 8514 1565 8520 1599
rect 8391 1547 8520 1565
rect 8351 1524 8520 1547
rect 8351 1509 8480 1524
rect 8351 1475 8357 1509
rect 8391 1490 8480 1509
rect 8514 1490 8520 1524
rect 8391 1475 8520 1490
rect 8351 1449 8520 1475
rect 8351 1437 8480 1449
rect 8351 1403 8357 1437
rect 8391 1415 8480 1437
rect 8514 1415 8520 1449
rect 8391 1403 8520 1415
rect 8351 1374 8520 1403
rect 8351 1365 8480 1374
rect 8351 1331 8357 1365
rect 8391 1340 8480 1365
rect 8514 1340 8520 1374
rect 8391 1331 8520 1340
rect 8637 1897 9009 1909
rect 8637 1863 8643 1897
rect 8677 1863 8969 1897
rect 9003 1863 9009 1897
rect 8637 1824 9009 1863
rect 8637 1790 8643 1824
rect 8677 1790 8969 1824
rect 9003 1790 9009 1824
rect 8637 1751 9009 1790
rect 8637 1717 8643 1751
rect 8677 1717 8969 1751
rect 9003 1717 9009 1751
rect 8637 1678 9009 1717
rect 8637 1644 8643 1678
rect 8677 1644 8969 1678
rect 9003 1644 9009 1678
rect 8637 1605 9009 1644
rect 8637 1571 8643 1605
rect 8677 1571 8969 1605
rect 9003 1571 9009 1605
rect 8637 1531 9009 1571
rect 8637 1497 8643 1531
rect 8677 1497 8969 1531
rect 9003 1497 9009 1531
rect 8637 1457 9009 1497
rect 8637 1423 8643 1457
rect 8677 1423 8969 1457
rect 9003 1423 9009 1457
rect 8637 1383 9009 1423
rect 8637 1349 8643 1383
rect 8677 1349 8969 1383
rect 9003 1349 9009 1383
rect 8637 1337 9009 1349
rect 9289 1897 9661 1909
rect 9289 1863 9295 1897
rect 9329 1863 9621 1897
rect 9655 1863 9661 1897
rect 9289 1824 9661 1863
rect 9289 1790 9295 1824
rect 9329 1790 9621 1824
rect 9655 1790 9661 1824
rect 9289 1751 9661 1790
rect 9289 1717 9295 1751
rect 9329 1717 9621 1751
rect 9655 1717 9661 1751
rect 9289 1678 9661 1717
rect 9289 1644 9295 1678
rect 9329 1644 9621 1678
rect 9655 1644 9661 1678
rect 9289 1605 9661 1644
rect 9289 1571 9295 1605
rect 9329 1571 9621 1605
rect 9655 1571 9661 1605
rect 9289 1531 9661 1571
rect 9289 1497 9295 1531
rect 9329 1497 9621 1531
rect 9655 1497 9661 1531
rect 9289 1457 9661 1497
rect 9289 1423 9295 1457
rect 9329 1423 9621 1457
rect 9655 1423 9661 1457
rect 9289 1383 9661 1423
rect 9289 1349 9295 1383
rect 9329 1349 9621 1383
rect 9655 1349 9661 1383
rect 9289 1337 9661 1349
rect 9957 1885 10003 1925
rect 9957 1851 9963 1885
rect 9997 1851 10003 1885
rect 9957 1811 10003 1851
rect 9957 1777 9963 1811
rect 9997 1777 10003 1811
rect 9957 1737 10003 1777
rect 9957 1703 9963 1737
rect 9997 1703 10003 1737
rect 9957 1663 10003 1703
rect 9957 1629 9963 1663
rect 9997 1629 10003 1663
rect 9957 1589 10003 1629
rect 9957 1555 9963 1589
rect 9997 1555 10003 1589
rect 9957 1515 10003 1555
rect 9957 1481 9963 1515
rect 9997 1481 10003 1515
rect 9957 1441 10003 1481
rect 9957 1407 9963 1441
rect 9997 1407 10003 1441
rect 9957 1366 10003 1407
rect 8351 1299 8520 1331
rect 8351 1293 8480 1299
rect 8351 1259 8357 1293
rect 8391 1265 8480 1293
rect 8514 1265 8520 1299
rect 8391 1259 8520 1265
tri 8234 1232 8237 1235 sw
rect 8185 1226 8237 1232
rect 8185 1157 8237 1174
rect 8185 1088 8237 1105
rect 8185 1019 8237 1036
rect 8185 950 8237 967
rect 8185 892 8237 898
tri 8185 889 8188 892 ne
rect 8025 827 8031 861
rect 8065 827 8071 861
rect 8025 789 8071 827
rect 8025 755 8031 789
rect 8065 755 8071 789
rect 8025 717 8071 755
rect 8025 683 8031 717
rect 8065 683 8071 717
rect 8025 645 8071 683
rect 8025 611 8031 645
rect 8065 611 8071 645
rect 8025 573 8071 611
rect 8025 539 8031 573
rect 8065 539 8071 573
rect 8025 527 8071 539
rect 8188 861 8234 892
tri 8234 889 8237 892 nw
rect 8351 1224 8520 1259
rect 8351 1221 8480 1224
rect 8351 1187 8357 1221
rect 8391 1190 8480 1221
rect 8514 1190 8520 1224
rect 9957 1332 9963 1366
rect 9997 1332 10003 1366
rect 9957 1291 10003 1332
rect 9957 1257 9963 1291
rect 9997 1257 10003 1291
rect 9957 1216 10003 1257
rect 8391 1187 8520 1190
rect 8351 1182 8520 1187
tri 8520 1182 8533 1195 sw
rect 9957 1182 9963 1216
rect 9997 1182 10003 1216
rect 8351 1170 8533 1182
tri 8533 1170 8545 1182 sw
rect 8351 1149 8545 1170
rect 8351 1115 8357 1149
rect 8391 1115 8480 1149
rect 8514 1141 8545 1149
tri 8545 1141 8574 1170 sw
rect 9957 1141 10003 1182
rect 8514 1115 8574 1141
rect 8351 1107 8574 1115
tri 8574 1107 8608 1141 sw
tri 9931 1107 9957 1133 se
rect 9957 1107 9963 1141
rect 9997 1107 10003 1141
rect 8351 1099 8608 1107
tri 8608 1099 8616 1107 sw
tri 9923 1099 9931 1107 se
rect 9931 1099 10003 1107
rect 8351 1093 10003 1099
rect 8351 1077 8494 1093
rect 8351 1043 8357 1077
rect 8391 1073 8494 1077
rect 8391 1043 8480 1073
rect 8351 1039 8480 1043
rect 8546 1041 8568 1093
rect 8620 1041 8642 1093
rect 8694 1041 8716 1093
rect 8768 1041 8790 1093
rect 8842 1087 10003 1093
rect 8842 1053 9132 1087
rect 9166 1053 9458 1087
rect 9492 1053 9784 1087
rect 9818 1066 10003 1087
rect 9818 1053 9963 1066
rect 8842 1041 9963 1053
rect 8514 1039 9963 1041
rect 8351 1032 9963 1039
rect 9997 1032 10003 1066
rect 8351 1023 10003 1032
rect 8351 1005 8494 1023
rect 8351 971 8357 1005
rect 8391 997 8494 1005
rect 8391 971 8480 997
rect 8546 971 8568 1023
rect 8620 971 8642 1023
rect 8694 971 8716 1023
rect 8768 971 8790 1023
rect 8842 1009 10003 1023
rect 8842 975 9132 1009
rect 9166 975 9458 1009
rect 9492 975 9784 1009
rect 9818 991 10003 1009
rect 9818 975 9963 991
rect 8842 971 9963 975
rect 8351 963 8480 971
rect 8514 963 9963 971
rect 8351 957 9963 963
rect 9997 957 10003 991
rect 8351 953 10003 957
rect 8351 933 8494 953
rect 8351 899 8357 933
rect 8391 921 8494 933
rect 8391 899 8480 921
rect 8546 901 8568 953
rect 8620 901 8642 953
rect 8694 901 8716 953
rect 8768 901 8790 953
rect 8842 931 10003 953
rect 8842 901 9132 931
rect 8188 827 8194 861
rect 8228 827 8234 861
rect 8188 789 8234 827
rect 8188 755 8194 789
rect 8228 755 8234 789
rect 8188 717 8234 755
rect 8188 683 8194 717
rect 8228 683 8234 717
rect 8188 645 8234 683
rect 8188 611 8194 645
rect 8228 611 8234 645
rect 8188 573 8234 611
rect 8188 539 8194 573
rect 8228 539 8234 573
rect 8188 527 8234 539
rect 8351 887 8480 899
rect 8514 897 8806 901
rect 8840 897 9132 901
rect 9166 897 9458 931
rect 9492 897 9784 931
rect 9818 916 10003 931
rect 9818 897 9963 916
rect 8514 887 9963 897
rect 8351 883 9963 887
rect 8351 861 8494 883
rect 8351 827 8357 861
rect 8391 845 8494 861
rect 8391 827 8480 845
rect 8546 831 8568 883
rect 8620 831 8642 883
rect 8694 831 8716 883
rect 8768 831 8790 883
rect 8842 882 9963 883
rect 9997 882 10003 916
rect 8842 853 10003 882
rect 8842 831 9132 853
rect 8351 811 8480 827
rect 8514 819 8806 831
rect 8840 819 9132 831
rect 9166 819 9458 853
rect 9492 819 9784 853
rect 9818 841 10003 853
rect 9818 819 9963 841
rect 8514 813 9963 819
rect 8351 789 8494 811
rect 8351 755 8357 789
rect 8391 769 8494 789
rect 8391 755 8480 769
rect 8546 761 8568 813
rect 8620 761 8642 813
rect 8694 761 8716 813
rect 8768 761 8790 813
rect 8842 807 9963 813
rect 9997 807 10003 841
rect 8842 775 10003 807
rect 8842 761 9132 775
rect 8351 735 8480 755
rect 8514 743 8806 761
rect 8840 743 9132 761
rect 8351 717 8494 735
rect 8351 683 8357 717
rect 8391 693 8494 717
rect 8391 683 8480 693
rect 8546 691 8568 743
rect 8620 691 8642 743
rect 8694 691 8716 743
rect 8768 691 8790 743
rect 8842 741 9132 743
rect 9166 741 9458 775
rect 9492 741 9784 775
rect 9818 766 10003 775
rect 9818 741 9963 766
rect 8842 732 9963 741
rect 9997 732 10003 766
rect 8842 697 10003 732
rect 8842 691 9132 697
rect 8351 659 8480 683
rect 8514 672 8806 691
rect 8840 672 9132 691
rect 8351 645 8494 659
rect 8351 611 8357 645
rect 8391 620 8494 645
rect 8546 620 8568 672
rect 8620 620 8642 672
rect 8694 620 8716 672
rect 8768 620 8790 672
rect 8842 663 9132 672
rect 9166 663 9458 697
rect 9492 663 9784 697
rect 9818 691 10003 697
rect 9818 663 9963 691
rect 8842 657 9963 663
rect 9997 657 10003 691
rect 8842 620 10003 657
rect 8391 619 10003 620
rect 8391 617 8806 619
rect 8391 611 8480 617
rect 8351 583 8480 611
rect 8514 585 8806 617
rect 8840 585 9132 619
rect 9166 585 9458 619
rect 9492 585 9784 619
rect 9818 616 10003 619
rect 9818 585 9963 616
rect 8514 583 9963 585
rect 8351 582 9963 583
rect 9997 582 10003 616
rect 8351 573 10003 582
rect 8351 539 8357 573
rect 8391 541 10003 573
rect 8391 539 8480 541
tri 8348 527 8351 530 se
rect 8351 527 8480 539
tri 8330 509 8348 527 se
rect 8348 509 8480 527
rect 7091 507 7137 509
tri 7137 507 7139 509 sw
tri 8328 507 8330 509 se
rect 8330 507 8480 509
rect 8514 507 8806 541
rect 8840 507 9132 541
rect 9166 507 9458 541
rect 9492 507 9784 541
rect 9818 507 9963 541
rect 9997 507 10003 541
rect 7091 477 7139 507
tri 7139 477 7169 507 sw
tri 8298 477 8328 507 se
rect 8328 477 10003 507
rect 7091 475 7169 477
tri 7169 475 7171 477 sw
tri 8296 475 8298 477 se
rect 8298 475 10003 477
rect 7091 469 10003 475
rect 7091 435 7169 469
rect 7203 435 7243 469
rect 7277 435 7317 469
rect 7351 435 7391 469
rect 7425 435 7465 469
rect 7499 435 7539 469
rect 7573 435 7613 469
rect 7647 435 7687 469
rect 7721 435 7761 469
rect 7795 435 7835 469
rect 7869 435 7909 469
rect 7943 435 7983 469
rect 8017 435 8057 469
rect 8091 435 8131 469
rect 8165 435 8205 469
rect 8239 435 8279 469
rect 8313 435 8353 469
rect 8387 435 8427 469
rect 8461 435 8501 469
rect 8535 435 8575 469
rect 8609 435 8649 469
rect 8683 435 8722 469
rect 8756 435 8795 469
rect 8829 435 8868 469
rect 8902 435 8941 469
rect 8975 435 9014 469
rect 9048 435 9087 469
rect 9121 435 9160 469
rect 9194 435 9233 469
rect 9267 435 9306 469
rect 9340 435 9379 469
rect 9413 435 9452 469
rect 9486 435 9525 469
rect 9559 435 9598 469
rect 9632 435 9671 469
rect 9705 435 9744 469
rect 9778 435 9817 469
rect 9851 435 9890 469
rect 9924 435 10003 469
rect 7091 429 10003 435
rect 10155 2106 10189 2140
rect 10223 2106 10257 2140
rect 10155 2068 10257 2106
rect 10155 2034 10189 2068
rect 10223 2034 10257 2068
rect 10155 1996 10257 2034
rect 10155 1962 10189 1996
rect 10223 1962 10257 1996
rect 10155 1924 10257 1962
rect 10155 1890 10189 1924
rect 10223 1890 10257 1924
rect 10155 1852 10257 1890
rect 10155 1818 10189 1852
rect 10223 1818 10257 1852
rect 10155 1780 10257 1818
rect 10155 1746 10189 1780
rect 10223 1746 10257 1780
rect 10155 1708 10257 1746
rect 10155 1674 10189 1708
rect 10223 1674 10257 1708
rect 10155 1636 10257 1674
rect 10155 1602 10189 1636
rect 10223 1602 10257 1636
rect 10155 1564 10257 1602
rect 10155 1530 10189 1564
rect 10223 1530 10257 1564
rect 10155 1492 10257 1530
rect 10155 1458 10189 1492
rect 10223 1458 10257 1492
rect 10155 1420 10257 1458
rect 10155 1386 10189 1420
rect 10223 1386 10257 1420
rect 10155 1348 10257 1386
rect 10155 1314 10189 1348
rect 10223 1314 10257 1348
rect 10155 1276 10257 1314
rect 10155 1242 10189 1276
rect 10223 1242 10257 1276
rect 10155 1204 10257 1242
rect 10155 1170 10189 1204
rect 10223 1170 10257 1204
rect 10155 1132 10257 1170
rect 10155 1098 10189 1132
rect 10223 1098 10257 1132
rect 10155 1060 10257 1098
rect 10155 1026 10189 1060
rect 10223 1026 10257 1060
rect 10155 988 10257 1026
rect 10155 954 10189 988
rect 10223 954 10257 988
rect 10155 915 10257 954
rect 10155 881 10189 915
rect 10223 881 10257 915
rect 10155 842 10257 881
rect 10155 808 10189 842
rect 10223 808 10257 842
rect 10155 769 10257 808
rect 10155 735 10189 769
rect 10223 735 10257 769
rect 10155 696 10257 735
rect 10155 662 10189 696
rect 10223 662 10257 696
rect 10155 623 10257 662
rect 10155 589 10189 623
rect 10223 589 10257 623
rect 10155 550 10257 589
rect 10155 516 10189 550
rect 10223 516 10257 550
rect 10155 477 10257 516
rect 10155 443 10189 477
rect 10223 443 10257 477
rect 6842 376 6944 415
rect 6842 342 6876 376
rect 6910 342 6944 376
rect 3750 270 3784 304
rect 3818 270 3852 304
rect 3750 230 3852 270
rect 3750 196 3784 230
rect 3818 196 3852 230
rect 3750 156 3852 196
rect 6842 303 6944 342
rect 6842 269 6876 303
rect 6910 269 6944 303
rect 10155 404 10257 443
rect 10155 370 10189 404
rect 10223 370 10257 404
rect 10155 331 10257 370
rect 10155 297 10189 331
rect 10223 297 10257 331
rect 6842 258 6944 269
tri 6944 258 6968 282 sw
tri 10131 258 10155 282 se
rect 10155 258 10257 297
rect 6842 248 6968 258
tri 6968 248 6978 258 sw
tri 10121 248 10131 258 se
rect 10131 248 10189 258
rect 6842 230 10189 248
rect 6842 196 6876 230
rect 6910 224 10189 230
rect 10223 224 10257 258
rect 6910 214 10257 224
rect 6910 196 6956 214
rect 6842 180 6956 196
rect 6990 180 7029 214
rect 7063 180 7102 214
rect 7136 180 7175 214
rect 7209 180 7248 214
rect 7282 180 7321 214
rect 7355 180 7394 214
rect 7428 180 7467 214
rect 7501 180 7540 214
rect 7574 180 7613 214
rect 7647 180 7686 214
rect 7720 180 7759 214
rect 7793 180 7832 214
rect 7866 180 7905 214
rect 7939 180 7978 214
rect 8012 180 8051 214
rect 8085 180 8124 214
rect 8158 180 8197 214
rect 8231 180 8270 214
rect 8304 180 8343 214
rect 8377 180 8416 214
rect 8450 180 8489 214
rect 8523 180 8561 214
rect 8595 180 8633 214
rect 8667 180 8705 214
rect 8739 180 8777 214
rect 8811 180 8849 214
rect 8883 180 8921 214
rect 8955 180 8993 214
rect 9027 180 9065 214
rect 9099 180 9137 214
rect 9171 180 9209 214
rect 9243 180 9281 214
rect 9315 180 9353 214
rect 9387 180 9425 214
rect 9459 180 9497 214
rect 9531 180 9569 214
rect 9603 180 9641 214
rect 9675 180 9713 214
rect 9747 180 9785 214
rect 9819 180 9857 214
rect 9891 180 9929 214
rect 9963 180 10001 214
rect 10035 180 10073 214
rect 10107 180 10257 214
rect 3750 122 3784 156
rect 3818 146 3852 156
tri 3852 146 3886 180 sw
tri 6808 146 6842 180 se
rect 6842 146 10257 180
rect 3818 138 6970 146
tri 6970 138 6978 146 nw
rect 3818 122 6944 138
rect 3750 112 6944 122
tri 6944 112 6970 138 nw
rect 3750 78 3902 112
rect 3936 78 3975 112
rect 4009 78 4048 112
rect 4082 78 4121 112
rect 4155 78 4194 112
rect 4228 78 4267 112
rect 4301 78 4340 112
rect 4374 78 4413 112
rect 4447 78 4486 112
rect 4520 78 4559 112
rect 4593 78 4632 112
rect 4666 78 4705 112
rect 4739 78 4778 112
rect 4812 78 4851 112
rect 4885 78 4924 112
rect 4958 78 4997 112
rect 5031 78 5070 112
rect 5104 78 5143 112
rect 5177 78 5216 112
rect 5250 78 5289 112
rect 5323 78 5362 112
rect 5396 78 5435 112
rect 5469 78 5508 112
rect 5542 78 5581 112
rect 5615 78 5654 112
rect 5688 78 5727 112
rect 5761 78 5800 112
rect 5834 78 5873 112
rect 5907 78 5946 112
rect 5980 78 6019 112
rect 6053 78 6092 112
rect 6126 78 6166 112
rect 6200 78 6240 112
rect 6274 78 6314 112
rect 6348 78 6388 112
rect 6422 78 6462 112
rect 6496 78 6536 112
rect 6570 78 6610 112
rect 6644 78 6684 112
rect 6718 78 6758 112
rect 6792 78 6832 112
rect 6866 78 6944 112
rect 3750 44 6944 78
<< via1 >>
rect 421 1957 473 1966
rect 421 1923 427 1957
rect 427 1923 461 1957
rect 461 1923 473 1957
rect 421 1914 473 1923
rect 485 1957 537 1966
rect 485 1923 506 1957
rect 506 1923 537 1957
rect 485 1914 537 1923
rect 353 1839 362 1873
rect 362 1839 396 1873
rect 396 1839 405 1873
rect 353 1821 405 1839
rect 353 1767 362 1800
rect 362 1767 396 1800
rect 396 1767 405 1800
rect 353 1748 405 1767
rect 353 1695 362 1726
rect 362 1695 396 1726
rect 396 1695 405 1726
rect 353 1674 405 1695
rect 353 1623 362 1652
rect 362 1623 396 1652
rect 396 1623 405 1652
rect 353 1600 405 1623
rect 353 1551 362 1578
rect 362 1551 396 1578
rect 396 1551 405 1578
rect 353 1526 405 1551
rect 353 1479 362 1504
rect 362 1479 396 1504
rect 396 1479 405 1504
rect 353 1452 405 1479
rect 353 1407 362 1430
rect 362 1407 396 1430
rect 396 1407 405 1430
rect 353 1378 405 1407
rect 679 1839 688 1873
rect 688 1839 722 1873
rect 722 1839 731 1873
rect 679 1821 731 1839
rect 679 1767 688 1800
rect 688 1767 722 1800
rect 722 1767 731 1800
rect 679 1748 731 1767
rect 679 1695 688 1726
rect 688 1695 722 1726
rect 722 1695 731 1726
rect 679 1674 731 1695
rect 679 1623 688 1652
rect 688 1623 722 1652
rect 722 1623 731 1652
rect 679 1600 731 1623
rect 679 1551 688 1578
rect 688 1551 722 1578
rect 722 1551 731 1578
rect 679 1526 731 1551
rect 679 1479 688 1504
rect 688 1479 722 1504
rect 722 1479 731 1504
rect 679 1452 731 1479
rect 679 1407 688 1430
rect 688 1407 722 1430
rect 722 1407 731 1430
rect 679 1378 731 1407
rect 1005 1839 1014 1853
rect 1014 1839 1048 1853
rect 1048 1839 1057 1853
rect 1005 1801 1057 1839
rect 1005 1767 1014 1775
rect 1014 1767 1048 1775
rect 1048 1767 1057 1775
rect 1005 1729 1057 1767
rect 1005 1723 1014 1729
rect 1014 1723 1048 1729
rect 1048 1723 1057 1729
rect 1005 1695 1014 1696
rect 1014 1695 1048 1696
rect 1048 1695 1057 1696
rect 1005 1657 1057 1695
rect 1005 1644 1014 1657
rect 1014 1644 1048 1657
rect 1048 1644 1057 1657
rect 1005 1585 1057 1617
rect 1005 1565 1014 1585
rect 1014 1565 1048 1585
rect 1048 1565 1057 1585
rect 1005 1513 1057 1538
rect 1005 1486 1014 1513
rect 1014 1486 1048 1513
rect 1048 1486 1057 1513
rect 1331 1839 1340 1853
rect 1340 1839 1374 1853
rect 1374 1839 1383 1853
rect 1331 1801 1383 1839
rect 1331 1767 1340 1775
rect 1340 1767 1374 1775
rect 1374 1767 1383 1775
rect 1331 1729 1383 1767
rect 1331 1723 1340 1729
rect 1340 1723 1374 1729
rect 1374 1723 1383 1729
rect 1331 1695 1340 1696
rect 1340 1695 1374 1696
rect 1374 1695 1383 1696
rect 1331 1657 1383 1695
rect 1331 1644 1340 1657
rect 1340 1644 1374 1657
rect 1374 1644 1383 1657
rect 1331 1585 1383 1617
rect 1331 1565 1340 1585
rect 1340 1565 1374 1585
rect 1374 1565 1383 1585
rect 1331 1513 1383 1538
rect 1331 1486 1340 1513
rect 1340 1486 1374 1513
rect 1374 1486 1383 1513
rect 516 793 568 803
rect 516 759 525 793
rect 525 759 559 793
rect 559 759 568 793
rect 516 751 568 759
rect 516 721 568 735
rect 516 687 525 721
rect 525 687 559 721
rect 559 687 568 721
rect 516 683 568 687
rect 516 649 568 666
rect 516 615 525 649
rect 525 615 559 649
rect 559 615 568 649
rect 516 614 568 615
rect 516 577 568 597
rect 516 545 525 577
rect 525 545 559 577
rect 559 545 568 577
rect 516 505 568 528
rect 516 476 525 505
rect 525 476 559 505
rect 559 476 568 505
rect 842 793 894 803
rect 842 759 851 793
rect 851 759 885 793
rect 885 759 894 793
rect 842 751 894 759
rect 842 721 894 735
rect 842 687 851 721
rect 851 687 885 721
rect 885 687 894 721
rect 842 683 894 687
rect 842 649 894 666
rect 842 615 851 649
rect 851 615 885 649
rect 885 615 894 649
rect 842 614 894 615
rect 842 577 894 597
rect 842 545 851 577
rect 851 545 885 577
rect 885 545 894 577
rect 842 505 894 528
rect 842 476 851 505
rect 851 476 885 505
rect 885 476 894 505
rect 1168 793 1220 803
rect 1168 759 1177 793
rect 1177 759 1211 793
rect 1211 759 1220 793
rect 1168 751 1220 759
rect 1168 721 1220 735
rect 1168 687 1177 721
rect 1177 687 1211 721
rect 1211 687 1220 721
rect 1168 683 1220 687
rect 1168 649 1220 666
rect 1168 615 1177 649
rect 1177 615 1211 649
rect 1211 615 1220 649
rect 1168 614 1220 615
rect 1168 577 1220 597
rect 1168 545 1177 577
rect 1177 545 1211 577
rect 1211 545 1220 577
rect 1168 505 1220 528
rect 1168 476 1177 505
rect 1177 476 1211 505
rect 1211 476 1220 505
rect 2297 1957 2349 1966
rect 2297 1923 2303 1957
rect 2303 1923 2337 1957
rect 2337 1923 2349 1957
rect 2297 1914 2349 1923
rect 2361 1957 2413 1966
rect 2361 1923 2382 1957
rect 2382 1923 2413 1957
rect 2361 1914 2413 1923
rect 3211 1955 3263 2005
rect 3211 1953 3220 1955
rect 3220 1953 3254 1955
rect 3254 1953 3263 1955
rect 2237 1225 2289 1226
rect 2237 1191 2246 1225
rect 2246 1191 2280 1225
rect 2280 1191 2289 1225
rect 2237 1174 2289 1191
rect 2237 1153 2289 1157
rect 2237 1119 2246 1153
rect 2246 1119 2280 1153
rect 2280 1119 2289 1153
rect 2237 1105 2289 1119
rect 2237 1081 2289 1088
rect 2237 1047 2246 1081
rect 2246 1047 2280 1081
rect 2280 1047 2289 1081
rect 2237 1036 2289 1047
rect 2237 1009 2289 1019
rect 2237 975 2246 1009
rect 2246 975 2280 1009
rect 2280 975 2289 1009
rect 2237 967 2289 975
rect 2237 937 2289 950
rect 2237 903 2246 937
rect 2246 903 2280 937
rect 2280 903 2289 937
rect 2237 898 2289 903
rect 2563 1225 2615 1226
rect 2563 1191 2572 1225
rect 2572 1191 2606 1225
rect 2606 1191 2615 1225
rect 2563 1174 2615 1191
rect 2563 1153 2615 1157
rect 2563 1119 2572 1153
rect 2572 1119 2606 1153
rect 2606 1119 2615 1153
rect 2563 1105 2615 1119
rect 2563 1081 2615 1088
rect 2563 1047 2572 1081
rect 2572 1047 2606 1081
rect 2606 1047 2615 1081
rect 2563 1036 2615 1047
rect 2563 1009 2615 1019
rect 2563 975 2572 1009
rect 2572 975 2606 1009
rect 2606 975 2615 1009
rect 2563 967 2615 975
rect 2563 937 2615 950
rect 2563 903 2572 937
rect 2572 903 2606 937
rect 2606 903 2615 937
rect 2563 898 2615 903
rect 2400 793 2452 803
rect 2400 759 2409 793
rect 2409 759 2443 793
rect 2443 759 2452 793
rect 2400 751 2452 759
rect 2400 721 2452 735
rect 2400 687 2409 721
rect 2409 687 2443 721
rect 2443 687 2452 721
rect 2400 683 2452 687
rect 2400 649 2452 666
rect 2400 615 2409 649
rect 2409 615 2443 649
rect 2443 615 2452 649
rect 2400 614 2452 615
rect 2400 577 2452 597
rect 2400 545 2409 577
rect 2409 545 2443 577
rect 2443 545 2452 577
rect 2400 505 2452 528
rect 2400 476 2409 505
rect 2409 476 2443 505
rect 2443 476 2452 505
rect 2889 1225 2941 1226
rect 2889 1191 2898 1225
rect 2898 1191 2932 1225
rect 2932 1191 2941 1225
rect 2889 1174 2941 1191
rect 2889 1153 2941 1157
rect 2889 1119 2898 1153
rect 2898 1119 2932 1153
rect 2932 1119 2941 1153
rect 2889 1105 2941 1119
rect 2889 1081 2941 1088
rect 2889 1047 2898 1081
rect 2898 1047 2932 1081
rect 2932 1047 2941 1081
rect 2889 1036 2941 1047
rect 2889 1009 2941 1019
rect 2889 975 2898 1009
rect 2898 975 2932 1009
rect 2932 975 2941 1009
rect 2889 967 2941 975
rect 2889 937 2941 950
rect 2889 903 2898 937
rect 2898 903 2932 937
rect 2932 903 2941 937
rect 2889 898 2941 903
rect 2726 793 2778 803
rect 2726 759 2735 793
rect 2735 759 2769 793
rect 2769 759 2778 793
rect 2726 751 2778 759
rect 2726 721 2778 735
rect 2726 687 2735 721
rect 2735 687 2769 721
rect 2769 687 2778 721
rect 2726 683 2778 687
rect 2726 649 2778 666
rect 2726 615 2735 649
rect 2735 615 2769 649
rect 2769 615 2778 649
rect 2726 614 2778 615
rect 2726 577 2778 597
rect 2726 545 2735 577
rect 2735 545 2769 577
rect 2769 545 2778 577
rect 2726 505 2778 528
rect 2726 476 2735 505
rect 2735 476 2769 505
rect 2769 476 2778 505
rect 3211 1882 3263 1920
rect 3211 1868 3220 1882
rect 3220 1868 3254 1882
rect 3254 1868 3263 1882
rect 3211 1809 3263 1835
rect 3211 1783 3220 1809
rect 3220 1783 3254 1809
rect 3254 1783 3263 1809
rect 3052 793 3104 803
rect 3052 759 3061 793
rect 3061 759 3095 793
rect 3095 759 3104 793
rect 3052 751 3104 759
rect 3052 721 3104 735
rect 3052 687 3061 721
rect 3061 687 3095 721
rect 3095 687 3104 721
rect 3052 683 3104 687
rect 3052 649 3104 666
rect 3052 615 3061 649
rect 3061 615 3095 649
rect 3095 615 3104 649
rect 3052 614 3104 615
rect 3052 577 3104 597
rect 3052 545 3061 577
rect 3061 545 3095 577
rect 3095 545 3104 577
rect 3052 505 3104 528
rect 3052 476 3061 505
rect 3061 476 3095 505
rect 3095 476 3104 505
rect 3775 1991 3827 2005
rect 3775 1957 3784 1991
rect 3784 1957 3818 1991
rect 3818 1957 3827 1991
rect 3775 1953 3827 1957
rect 3775 1918 3827 1920
rect 3775 1884 3784 1918
rect 3784 1884 3818 1918
rect 3818 1884 3827 1918
rect 3775 1868 3827 1884
rect 3775 1811 3784 1835
rect 3784 1811 3818 1835
rect 3818 1811 3827 1835
rect 3775 1783 3827 1811
rect 4612 1957 4664 1966
rect 4612 1923 4615 1957
rect 4615 1923 4649 1957
rect 4649 1923 4664 1957
rect 4612 1914 4664 1923
rect 4676 1957 4728 1966
rect 4676 1923 4688 1957
rect 4688 1923 4722 1957
rect 4722 1923 4728 1957
rect 4676 1914 4728 1923
rect 5897 1957 5949 1966
rect 5897 1923 5913 1957
rect 5913 1923 5947 1957
rect 5947 1923 5949 1957
rect 5897 1914 5949 1923
rect 5976 1957 6028 1966
rect 5976 1923 5988 1957
rect 5988 1923 6022 1957
rect 6022 1923 6028 1957
rect 5976 1914 6028 1923
rect 4285 1225 4337 1226
rect 4285 1191 4294 1225
rect 4294 1191 4328 1225
rect 4328 1191 4337 1225
rect 4285 1174 4337 1191
rect 4285 1153 4337 1157
rect 4285 1119 4294 1153
rect 4294 1119 4328 1153
rect 4328 1119 4337 1153
rect 4285 1105 4337 1119
rect 4285 1081 4337 1088
rect 4285 1047 4294 1081
rect 4294 1047 4328 1081
rect 4328 1047 4337 1081
rect 4285 1036 4337 1047
rect 4285 1009 4337 1019
rect 4285 975 4294 1009
rect 4294 975 4328 1009
rect 4328 975 4337 1009
rect 4285 967 4337 975
rect 4285 937 4337 950
rect 4285 903 4294 937
rect 4294 903 4328 937
rect 4328 903 4337 937
rect 4285 898 4337 903
rect 3996 780 4005 803
rect 4005 780 4039 803
rect 4039 780 4048 803
rect 3996 751 4048 780
rect 3996 705 4005 735
rect 4005 705 4039 735
rect 4039 705 4048 735
rect 3996 683 4048 705
rect 3996 664 4048 666
rect 3996 630 4005 664
rect 4005 630 4039 664
rect 4039 630 4048 664
rect 3996 614 4048 630
rect 3996 589 4048 597
rect 3996 555 4005 589
rect 4005 555 4039 589
rect 4039 555 4048 589
rect 3996 545 4048 555
rect 3996 514 4048 528
rect 3996 480 4005 514
rect 4005 480 4039 514
rect 4039 480 4048 514
rect 3996 476 4048 480
rect 4122 793 4174 803
rect 4122 759 4131 793
rect 4131 759 4165 793
rect 4165 759 4174 793
rect 4122 751 4174 759
rect 4122 721 4174 735
rect 4122 687 4131 721
rect 4131 687 4165 721
rect 4165 687 4174 721
rect 4122 683 4174 687
rect 4122 649 4174 666
rect 4122 615 4131 649
rect 4131 615 4165 649
rect 4165 615 4174 649
rect 4122 614 4174 615
rect 4122 577 4174 597
rect 4122 545 4131 577
rect 4131 545 4165 577
rect 4165 545 4174 577
rect 4122 505 4174 528
rect 4122 476 4131 505
rect 4131 476 4165 505
rect 4165 476 4174 505
rect 4611 1225 4663 1226
rect 4611 1191 4620 1225
rect 4620 1191 4654 1225
rect 4654 1191 4663 1225
rect 4611 1174 4663 1191
rect 4611 1153 4663 1157
rect 4611 1119 4620 1153
rect 4620 1119 4654 1153
rect 4654 1119 4663 1153
rect 4611 1105 4663 1119
rect 4611 1081 4663 1088
rect 4611 1047 4620 1081
rect 4620 1047 4654 1081
rect 4654 1047 4663 1081
rect 4611 1036 4663 1047
rect 4611 1009 4663 1019
rect 4611 975 4620 1009
rect 4620 975 4654 1009
rect 4654 975 4663 1009
rect 4611 967 4663 975
rect 4611 937 4663 950
rect 4611 903 4620 937
rect 4620 903 4654 937
rect 4654 903 4663 937
rect 4611 898 4663 903
rect 4448 793 4500 803
rect 4448 759 4457 793
rect 4457 759 4491 793
rect 4491 759 4500 793
rect 4448 751 4500 759
rect 4448 721 4500 735
rect 4448 687 4457 721
rect 4457 687 4491 721
rect 4491 687 4500 721
rect 4448 683 4500 687
rect 4448 649 4500 666
rect 4448 615 4457 649
rect 4457 615 4491 649
rect 4491 615 4500 649
rect 4448 614 4500 615
rect 4448 577 4500 597
rect 4448 545 4457 577
rect 4457 545 4491 577
rect 4491 545 4500 577
rect 4448 505 4500 528
rect 4448 476 4457 505
rect 4457 476 4491 505
rect 4491 476 4500 505
rect 4937 1225 4989 1226
rect 4937 1191 4946 1225
rect 4946 1191 4980 1225
rect 4980 1191 4989 1225
rect 4937 1174 4989 1191
rect 4937 1153 4989 1157
rect 4937 1119 4946 1153
rect 4946 1119 4980 1153
rect 4980 1119 4989 1153
rect 4937 1105 4989 1119
rect 4937 1081 4989 1088
rect 4937 1047 4946 1081
rect 4946 1047 4980 1081
rect 4980 1047 4989 1081
rect 4937 1036 4989 1047
rect 4937 1009 4989 1019
rect 4937 975 4946 1009
rect 4946 975 4980 1009
rect 4980 975 4989 1009
rect 4937 967 4989 975
rect 4937 937 4989 950
rect 4937 903 4946 937
rect 4946 903 4980 937
rect 4980 903 4989 937
rect 4937 898 4989 903
rect 5386 1695 5395 1717
rect 5395 1695 5429 1717
rect 5429 1695 5438 1717
rect 5386 1665 5438 1695
rect 5386 1623 5395 1638
rect 5395 1623 5429 1638
rect 5429 1623 5438 1638
rect 5386 1586 5438 1623
rect 5386 1551 5395 1559
rect 5395 1551 5429 1559
rect 5429 1551 5438 1559
rect 5386 1513 5438 1551
rect 5386 1507 5395 1513
rect 5395 1507 5429 1513
rect 5429 1507 5438 1513
rect 5386 1479 5395 1480
rect 5395 1479 5429 1480
rect 5429 1479 5438 1480
rect 5386 1441 5438 1479
rect 5386 1428 5395 1441
rect 5395 1428 5429 1441
rect 5429 1428 5438 1441
rect 5386 1369 5438 1401
rect 5386 1349 5395 1369
rect 5395 1349 5429 1369
rect 5429 1349 5438 1369
rect 4774 793 4826 803
rect 4774 759 4783 793
rect 4783 759 4817 793
rect 4817 759 4826 793
rect 4774 751 4826 759
rect 4774 721 4826 735
rect 4774 687 4783 721
rect 4783 687 4817 721
rect 4817 687 4826 721
rect 4774 683 4826 687
rect 4774 649 4826 666
rect 4774 615 4783 649
rect 4783 615 4817 649
rect 4817 615 4826 649
rect 4774 614 4826 615
rect 4774 577 4826 597
rect 4774 545 4783 577
rect 4783 545 4817 577
rect 4817 545 4826 577
rect 4774 505 4826 528
rect 4774 476 4783 505
rect 4783 476 4817 505
rect 4817 476 4826 505
rect 5263 1225 5315 1226
rect 5263 1191 5272 1225
rect 5272 1191 5306 1225
rect 5306 1191 5315 1225
rect 5263 1174 5315 1191
rect 5263 1153 5315 1157
rect 5263 1119 5272 1153
rect 5272 1119 5306 1153
rect 5306 1119 5315 1153
rect 5263 1105 5315 1119
rect 5263 1081 5315 1088
rect 5263 1047 5272 1081
rect 5272 1047 5306 1081
rect 5306 1047 5315 1081
rect 5263 1036 5315 1047
rect 5263 1009 5315 1019
rect 5263 975 5272 1009
rect 5272 975 5306 1009
rect 5306 975 5315 1009
rect 5263 967 5315 975
rect 5263 937 5315 950
rect 5263 903 5272 937
rect 5272 903 5306 937
rect 5306 903 5315 937
rect 5263 898 5315 903
rect 5100 793 5152 803
rect 5100 759 5109 793
rect 5109 759 5143 793
rect 5143 759 5152 793
rect 5100 751 5152 759
rect 5100 721 5152 735
rect 5100 687 5109 721
rect 5109 687 5143 721
rect 5143 687 5152 721
rect 5100 683 5152 687
rect 5100 649 5152 666
rect 5100 615 5109 649
rect 5109 615 5143 649
rect 5143 615 5152 649
rect 5100 614 5152 615
rect 5100 577 5152 597
rect 5100 545 5109 577
rect 5109 545 5143 577
rect 5143 545 5152 577
rect 5100 505 5152 528
rect 5100 476 5109 505
rect 5109 476 5143 505
rect 5143 476 5152 505
rect 5712 1695 5721 1717
rect 5721 1695 5755 1717
rect 5755 1695 5764 1717
rect 5712 1665 5764 1695
rect 5712 1623 5721 1638
rect 5721 1623 5755 1638
rect 5755 1623 5764 1638
rect 5712 1586 5764 1623
rect 5712 1551 5721 1559
rect 5721 1551 5755 1559
rect 5755 1551 5764 1559
rect 5712 1513 5764 1551
rect 5712 1507 5721 1513
rect 5721 1507 5755 1513
rect 5755 1507 5764 1513
rect 5712 1479 5721 1480
rect 5721 1479 5755 1480
rect 5755 1479 5764 1480
rect 5712 1441 5764 1479
rect 5712 1428 5721 1441
rect 5721 1428 5755 1441
rect 5755 1428 5764 1441
rect 5712 1369 5764 1401
rect 5712 1349 5721 1369
rect 5721 1349 5755 1369
rect 5755 1349 5764 1369
rect 5549 793 5601 803
rect 5549 759 5558 793
rect 5558 759 5592 793
rect 5592 759 5601 793
rect 5549 751 5601 759
rect 5549 721 5601 735
rect 5549 687 5558 721
rect 5558 687 5592 721
rect 5592 687 5601 721
rect 5549 683 5601 687
rect 5549 649 5601 666
rect 5549 615 5558 649
rect 5558 615 5592 649
rect 5592 615 5601 649
rect 5549 614 5601 615
rect 5549 577 5601 597
rect 5549 545 5558 577
rect 5558 545 5592 577
rect 5592 545 5601 577
rect 5549 505 5601 528
rect 5549 476 5558 505
rect 5558 476 5592 505
rect 5592 476 5601 505
rect 6038 1695 6047 1717
rect 6047 1695 6081 1717
rect 6081 1695 6090 1717
rect 6038 1665 6090 1695
rect 6038 1623 6047 1638
rect 6047 1623 6081 1638
rect 6081 1623 6090 1638
rect 6038 1586 6090 1623
rect 6038 1551 6047 1559
rect 6047 1551 6081 1559
rect 6081 1551 6090 1559
rect 6038 1513 6090 1551
rect 6038 1507 6047 1513
rect 6047 1507 6081 1513
rect 6081 1507 6090 1513
rect 6038 1479 6047 1480
rect 6047 1479 6081 1480
rect 6081 1479 6090 1480
rect 6038 1441 6090 1479
rect 6038 1428 6047 1441
rect 6047 1428 6081 1441
rect 6081 1428 6090 1441
rect 6038 1369 6090 1401
rect 6038 1349 6047 1369
rect 6047 1349 6081 1369
rect 6081 1349 6090 1369
rect 5875 793 5927 803
rect 5875 759 5884 793
rect 5884 759 5918 793
rect 5918 759 5927 793
rect 5875 751 5927 759
rect 5875 721 5927 735
rect 5875 687 5884 721
rect 5884 687 5918 721
rect 5918 687 5927 721
rect 5875 683 5927 687
rect 5875 649 5927 666
rect 5875 615 5884 649
rect 5884 615 5918 649
rect 5918 615 5927 649
rect 5875 614 5927 615
rect 5875 577 5927 597
rect 5875 545 5884 577
rect 5884 545 5918 577
rect 5918 545 5927 577
rect 5875 505 5927 528
rect 5875 476 5884 505
rect 5884 476 5918 505
rect 5918 476 5927 505
rect 6364 1695 6373 1717
rect 6373 1695 6407 1717
rect 6407 1695 6416 1717
rect 6364 1665 6416 1695
rect 6364 1623 6373 1638
rect 6373 1623 6407 1638
rect 6407 1623 6416 1638
rect 6364 1586 6416 1623
rect 6364 1551 6373 1559
rect 6373 1551 6407 1559
rect 6407 1551 6416 1559
rect 6364 1513 6416 1551
rect 6364 1507 6373 1513
rect 6373 1507 6407 1513
rect 6407 1507 6416 1513
rect 6364 1479 6373 1480
rect 6373 1479 6407 1480
rect 6407 1479 6416 1480
rect 6364 1441 6416 1479
rect 6364 1428 6373 1441
rect 6373 1428 6407 1441
rect 6407 1428 6416 1441
rect 6364 1369 6416 1401
rect 6364 1349 6373 1369
rect 6373 1349 6407 1369
rect 6407 1349 6416 1369
rect 6201 793 6253 803
rect 6201 759 6210 793
rect 6210 759 6244 793
rect 6244 759 6253 793
rect 6201 751 6253 759
rect 6201 721 6253 735
rect 6201 687 6210 721
rect 6210 687 6244 721
rect 6244 687 6253 721
rect 6201 683 6253 687
rect 6201 649 6253 666
rect 6201 615 6210 649
rect 6210 615 6244 649
rect 6244 615 6253 649
rect 6201 614 6253 615
rect 6201 577 6253 597
rect 6201 545 6210 577
rect 6210 545 6244 577
rect 6244 545 6253 577
rect 6201 505 6253 528
rect 6201 476 6210 505
rect 6210 476 6244 505
rect 6244 476 6253 505
rect 7286 2025 7338 2034
rect 7351 2025 7403 2034
rect 7286 1991 7307 2025
rect 7307 1991 7338 2025
rect 7351 1991 7380 2025
rect 7380 1991 7403 2025
rect 7286 1982 7338 1991
rect 7351 1982 7403 1991
rect 7416 2025 7468 2034
rect 7416 1991 7419 2025
rect 7419 1991 7453 2025
rect 7453 1991 7468 2025
rect 7416 1982 7468 1991
rect 7481 2025 7533 2034
rect 7481 1991 7492 2025
rect 7492 1991 7526 2025
rect 7526 1991 7533 2025
rect 7481 1982 7533 1991
rect 7546 2025 7598 2034
rect 7611 2025 7663 2034
rect 7676 2025 7728 2034
rect 7546 1991 7565 2025
rect 7565 1991 7598 2025
rect 7611 1991 7638 2025
rect 7638 1991 7663 2025
rect 7676 1991 7711 2025
rect 7711 1991 7728 2025
rect 7546 1982 7598 1991
rect 7611 1982 7663 1991
rect 7676 1982 7728 1991
rect 8248 1982 8300 2034
rect 8312 1982 8364 2034
rect 7088 1701 7097 1732
rect 7097 1701 7131 1732
rect 7131 1701 7140 1732
rect 7088 1680 7140 1701
rect 7088 1660 7140 1661
rect 7088 1626 7097 1660
rect 7097 1626 7131 1660
rect 7131 1626 7140 1660
rect 7088 1609 7140 1626
rect 7088 1585 7140 1590
rect 7088 1551 7097 1585
rect 7097 1551 7131 1585
rect 7131 1551 7140 1585
rect 7088 1538 7140 1551
rect 7088 1510 7140 1518
rect 7088 1476 7097 1510
rect 7097 1476 7131 1510
rect 7131 1476 7140 1510
rect 7088 1466 7140 1476
rect 7088 1435 7140 1446
rect 7088 1401 7097 1435
rect 7097 1401 7131 1435
rect 7131 1401 7140 1435
rect 7088 1394 7140 1401
rect 6527 793 6579 803
rect 6527 759 6536 793
rect 6536 759 6570 793
rect 6570 759 6579 793
rect 6527 751 6579 759
rect 6527 721 6579 735
rect 6527 687 6536 721
rect 6536 687 6570 721
rect 6570 687 6579 721
rect 6527 683 6579 687
rect 6527 649 6579 666
rect 6527 615 6536 649
rect 6536 615 6570 649
rect 6570 615 6579 649
rect 6527 614 6579 615
rect 6527 577 6579 597
rect 6527 545 6536 577
rect 6536 545 6570 577
rect 6570 545 6579 577
rect 6527 505 6579 528
rect 6527 476 6536 505
rect 6536 476 6570 505
rect 6570 476 6579 505
rect 6646 777 6655 803
rect 6655 777 6689 803
rect 6689 777 6698 803
rect 6646 751 6698 777
rect 6646 703 6655 735
rect 6655 703 6689 735
rect 6689 703 6698 735
rect 6646 683 6698 703
rect 6646 663 6698 666
rect 6646 629 6655 663
rect 6655 629 6689 663
rect 6689 629 6698 663
rect 6646 614 6698 629
rect 6646 589 6698 597
rect 6646 555 6655 589
rect 6655 555 6689 589
rect 6689 555 6698 589
rect 6646 545 6698 555
rect 6646 515 6698 528
rect 6646 481 6655 515
rect 6655 481 6689 515
rect 6689 481 6698 515
rect 6646 476 6698 481
rect 7370 1725 7422 1732
rect 7370 1691 7379 1725
rect 7379 1691 7413 1725
rect 7413 1691 7422 1725
rect 7370 1680 7422 1691
rect 7370 1653 7422 1661
rect 7370 1619 7379 1653
rect 7379 1619 7413 1653
rect 7413 1619 7422 1653
rect 7370 1609 7422 1619
rect 7370 1581 7422 1590
rect 7370 1547 7379 1581
rect 7379 1547 7413 1581
rect 7413 1547 7422 1581
rect 7370 1538 7422 1547
rect 7370 1509 7422 1518
rect 7370 1475 7379 1509
rect 7379 1475 7413 1509
rect 7413 1475 7422 1509
rect 7370 1466 7422 1475
rect 7370 1437 7422 1446
rect 7370 1403 7379 1437
rect 7379 1403 7413 1437
rect 7413 1403 7422 1437
rect 7370 1394 7422 1403
rect 7207 1221 7259 1226
rect 7207 1187 7216 1221
rect 7216 1187 7250 1221
rect 7250 1187 7259 1221
rect 7207 1174 7259 1187
rect 7207 1149 7259 1157
rect 7207 1115 7216 1149
rect 7216 1115 7250 1149
rect 7250 1115 7259 1149
rect 7207 1105 7259 1115
rect 7207 1077 7259 1088
rect 7207 1043 7216 1077
rect 7216 1043 7250 1077
rect 7250 1043 7259 1077
rect 7207 1036 7259 1043
rect 7207 1005 7259 1019
rect 7207 971 7216 1005
rect 7216 971 7250 1005
rect 7250 971 7259 1005
rect 7207 967 7259 971
rect 7207 933 7259 950
rect 7207 899 7216 933
rect 7216 899 7250 933
rect 7250 899 7259 933
rect 7207 898 7259 899
rect 7696 1725 7748 1732
rect 7696 1691 7705 1725
rect 7705 1691 7739 1725
rect 7739 1691 7748 1725
rect 7696 1680 7748 1691
rect 7696 1653 7748 1661
rect 7696 1619 7705 1653
rect 7705 1619 7739 1653
rect 7739 1619 7748 1653
rect 7696 1609 7748 1619
rect 7696 1581 7748 1590
rect 7696 1547 7705 1581
rect 7705 1547 7739 1581
rect 7739 1547 7748 1581
rect 7696 1538 7748 1547
rect 7696 1509 7748 1518
rect 7696 1475 7705 1509
rect 7705 1475 7739 1509
rect 7739 1475 7748 1509
rect 7696 1466 7748 1475
rect 7696 1437 7748 1446
rect 7696 1403 7705 1437
rect 7705 1403 7739 1437
rect 7739 1403 7748 1437
rect 7696 1394 7748 1403
rect 7533 1221 7585 1226
rect 7533 1187 7542 1221
rect 7542 1187 7576 1221
rect 7576 1187 7585 1221
rect 7533 1174 7585 1187
rect 7533 1149 7585 1157
rect 7533 1115 7542 1149
rect 7542 1115 7576 1149
rect 7576 1115 7585 1149
rect 7533 1105 7585 1115
rect 7533 1077 7585 1088
rect 7533 1043 7542 1077
rect 7542 1043 7576 1077
rect 7576 1043 7585 1077
rect 7533 1036 7585 1043
rect 7533 1005 7585 1019
rect 7533 971 7542 1005
rect 7542 971 7576 1005
rect 7576 971 7585 1005
rect 7533 967 7585 971
rect 7533 933 7585 950
rect 7533 899 7542 933
rect 7542 899 7576 933
rect 7576 899 7585 933
rect 7533 898 7585 899
rect 8022 1725 8074 1732
rect 8022 1691 8031 1725
rect 8031 1691 8065 1725
rect 8065 1691 8074 1725
rect 8022 1680 8074 1691
rect 8022 1653 8074 1661
rect 8022 1619 8031 1653
rect 8031 1619 8065 1653
rect 8065 1619 8074 1653
rect 8022 1609 8074 1619
rect 8022 1581 8074 1590
rect 8022 1547 8031 1581
rect 8031 1547 8065 1581
rect 8065 1547 8074 1581
rect 8022 1538 8074 1547
rect 8022 1509 8074 1518
rect 8022 1475 8031 1509
rect 8031 1475 8065 1509
rect 8065 1475 8074 1509
rect 8022 1466 8074 1475
rect 8022 1437 8074 1446
rect 8022 1403 8031 1437
rect 8031 1403 8065 1437
rect 8065 1403 8074 1437
rect 8022 1394 8074 1403
rect 7859 1221 7911 1226
rect 7859 1187 7868 1221
rect 7868 1187 7902 1221
rect 7902 1187 7911 1221
rect 7859 1174 7911 1187
rect 7859 1149 7911 1157
rect 7859 1115 7868 1149
rect 7868 1115 7902 1149
rect 7902 1115 7911 1149
rect 7859 1105 7911 1115
rect 7859 1077 7911 1088
rect 7859 1043 7868 1077
rect 7868 1043 7902 1077
rect 7902 1043 7911 1077
rect 7859 1036 7911 1043
rect 7859 1005 7911 1019
rect 7859 971 7868 1005
rect 7868 971 7902 1005
rect 7902 971 7911 1005
rect 7859 967 7911 971
rect 7859 933 7911 950
rect 7859 899 7868 933
rect 7868 899 7902 933
rect 7902 899 7911 933
rect 7859 898 7911 899
rect 8185 1221 8237 1226
rect 8185 1187 8194 1221
rect 8194 1187 8228 1221
rect 8228 1187 8237 1221
rect 8185 1174 8237 1187
rect 8185 1149 8237 1157
rect 8185 1115 8194 1149
rect 8194 1115 8228 1149
rect 8228 1115 8237 1149
rect 8185 1105 8237 1115
rect 8185 1077 8237 1088
rect 8185 1043 8194 1077
rect 8194 1043 8228 1077
rect 8228 1043 8237 1077
rect 8185 1036 8237 1043
rect 8185 1005 8237 1019
rect 8185 971 8194 1005
rect 8194 971 8228 1005
rect 8228 971 8237 1005
rect 8185 967 8237 971
rect 8185 933 8237 950
rect 8185 899 8194 933
rect 8194 899 8228 933
rect 8228 899 8237 933
rect 8185 898 8237 899
rect 8494 1073 8546 1093
rect 8494 1041 8514 1073
rect 8514 1041 8546 1073
rect 8568 1041 8620 1093
rect 8642 1041 8694 1093
rect 8716 1041 8768 1093
rect 8790 1087 8842 1093
rect 8790 1053 8806 1087
rect 8806 1053 8840 1087
rect 8840 1053 8842 1087
rect 8790 1041 8842 1053
rect 8494 997 8546 1023
rect 8494 971 8514 997
rect 8514 971 8546 997
rect 8568 971 8620 1023
rect 8642 971 8694 1023
rect 8716 971 8768 1023
rect 8790 1009 8842 1023
rect 8790 975 8806 1009
rect 8806 975 8840 1009
rect 8840 975 8842 1009
rect 8790 971 8842 975
rect 8494 921 8546 953
rect 8494 901 8514 921
rect 8514 901 8546 921
rect 8568 901 8620 953
rect 8642 901 8694 953
rect 8716 901 8768 953
rect 8790 931 8842 953
rect 8790 901 8806 931
rect 8806 901 8840 931
rect 8840 901 8842 931
rect 8494 845 8546 883
rect 8494 831 8514 845
rect 8514 831 8546 845
rect 8568 831 8620 883
rect 8642 831 8694 883
rect 8716 831 8768 883
rect 8790 853 8842 883
rect 8790 831 8806 853
rect 8806 831 8840 853
rect 8840 831 8842 853
rect 8494 811 8514 813
rect 8514 811 8546 813
rect 8494 769 8546 811
rect 8494 761 8514 769
rect 8514 761 8546 769
rect 8568 761 8620 813
rect 8642 761 8694 813
rect 8716 761 8768 813
rect 8790 775 8842 813
rect 8790 761 8806 775
rect 8806 761 8840 775
rect 8840 761 8842 775
rect 8494 735 8514 743
rect 8514 735 8546 743
rect 8494 693 8546 735
rect 8494 691 8514 693
rect 8514 691 8546 693
rect 8568 691 8620 743
rect 8642 691 8694 743
rect 8716 691 8768 743
rect 8790 741 8806 743
rect 8806 741 8840 743
rect 8840 741 8842 743
rect 8790 697 8842 741
rect 8790 691 8806 697
rect 8806 691 8840 697
rect 8840 691 8842 697
rect 8494 659 8514 672
rect 8514 659 8546 672
rect 8494 620 8546 659
rect 8568 620 8620 672
rect 8642 620 8694 672
rect 8716 620 8768 672
rect 8790 663 8806 672
rect 8806 663 8840 672
rect 8840 663 8842 672
rect 8790 620 8842 663
<< metal2 >>
rect -24 2188 3941 2213
tri 3941 2188 3966 2213 sw
rect -24 2161 3966 2188
tri 3919 2128 3952 2161 ne
rect 3952 2128 3966 2161
tri 3966 2128 4026 2188 sw
rect -24 2115 3906 2128
tri 3906 2115 3919 2128 sw
tri 3952 2115 3965 2128 ne
rect 3965 2115 4026 2128
rect -24 2114 3919 2115
tri 3919 2114 3920 2115 sw
tri 3965 2114 3966 2115 ne
rect 3966 2114 4026 2115
tri 4026 2114 4040 2128 sw
rect -24 2092 3920 2114
tri 3920 2092 3942 2114 sw
tri 3966 2092 3988 2114 ne
rect 3988 2092 4040 2114
tri 4040 2092 4062 2114 sw
rect -24 2076 3942 2092
tri 3884 2048 3912 2076 ne
rect 3912 2074 3942 2076
tri 3942 2074 3960 2092 sw
tri 3988 2074 4006 2092 ne
rect 4006 2074 4062 2092
tri 4062 2074 4080 2092 sw
rect 3912 2068 3960 2074
tri 3960 2068 3966 2074 sw
tri 4006 2068 4012 2074 ne
rect 4012 2068 4080 2074
rect 3912 2048 3966 2068
rect -24 2040 2174 2048
tri 2174 2040 2182 2048 sw
tri 3912 2040 3920 2048 ne
rect 3920 2040 3966 2048
tri 3966 2040 3994 2068 sw
tri 4012 2040 4040 2068 ne
rect 4040 2040 4080 2068
tri 4080 2040 4114 2074 sw
tri 5643 2040 5677 2074 se
rect 5677 2040 7225 2074
rect -24 2034 2182 2040
tri 2182 2034 2188 2040 sw
tri 3920 2034 3926 2040 ne
rect 3926 2034 3994 2040
tri 3994 2034 4000 2040 sw
tri 4040 2034 4046 2040 ne
rect 4046 2034 4114 2040
tri 4114 2034 4120 2040 sw
tri 5637 2034 5643 2040 se
rect 5643 2034 7225 2040
tri 7225 2034 7265 2074 sw
rect -24 2018 2188 2034
tri 2188 2018 2204 2034 sw
tri 3926 2018 3942 2034 ne
rect 3942 2022 4000 2034
tri 4000 2022 4012 2034 sw
tri 4046 2022 4058 2034 ne
rect 4058 2022 4120 2034
tri 4120 2022 4132 2034 sw
tri 5625 2022 5637 2034 se
rect 5637 2022 7286 2034
rect 3942 2018 4012 2022
tri 4012 2018 4016 2022 sw
tri 4058 2018 4062 2022 ne
rect 4062 2018 4132 2022
tri 4132 2018 4136 2022 sw
tri 5621 2018 5625 2022 se
rect 5625 2018 5697 2022
rect -24 2011 2204 2018
tri 2204 2011 2211 2018 sw
tri 3942 2011 3949 2018 ne
rect 3949 2011 4016 2018
tri 4016 2011 4023 2018 sw
tri 4062 2011 4069 2018 ne
rect 4069 2011 4136 2018
tri 4136 2011 4143 2018 sw
tri 5614 2011 5621 2018 se
rect 5621 2011 5697 2018
tri 5697 2011 5708 2022 nw
tri 7183 2011 7194 2022 ne
rect 7194 2011 7286 2022
rect -24 2005 2211 2011
tri 2211 2005 2217 2011 sw
rect 3186 2005 3852 2011
rect -24 1996 2217 2005
tri 2152 1968 2180 1996 ne
rect 2180 1968 2217 1996
rect -24 1966 581 1968
tri 2180 1966 2182 1968 ne
rect 2182 1966 2217 1968
tri 2217 1966 2256 2005 sw
rect -24 1914 421 1966
rect 473 1914 485 1966
rect 537 1914 581 1966
tri 2182 1914 2234 1966 ne
rect 2234 1914 2297 1966
rect 2349 1914 2361 1966
rect 2413 1914 2419 1966
rect 3186 1953 3211 2005
rect 3263 1953 3775 2005
rect 3827 1953 3852 2005
tri 3949 1982 3978 2011 ne
rect 3978 1994 4023 2011
tri 4023 1994 4040 2011 sw
tri 4069 1994 4086 2011 ne
rect 4086 1994 4143 2011
rect 3978 1982 4040 1994
tri 4040 1982 4052 1994 sw
tri 4086 1982 4098 1994 ne
rect 4098 1982 4143 1994
tri 4143 1982 4172 2011 sw
tri 5585 1982 5614 2011 se
rect 5614 1982 5668 2011
tri 5668 1982 5697 2011 nw
tri 7194 1982 7223 2011 ne
rect 7223 1982 7286 2011
rect 7338 1982 7351 2034
rect 7403 1982 7416 2034
rect 7468 1982 7481 2034
rect 7533 1982 7546 2034
rect 7598 1982 7611 2034
rect 7663 1982 7676 2034
rect 7728 1982 7734 2034
tri 8198 1982 8242 2026 se
rect 8242 1982 8248 2034
rect 8300 1982 8312 2034
rect 8364 1982 8370 2034
tri 3978 1966 3994 1982 ne
rect 3994 1966 4052 1982
tri 4052 1966 4068 1982 sw
tri 4098 1966 4114 1982 ne
rect 4114 1966 4172 1982
tri 4172 1966 4188 1982 sw
tri 5569 1966 5585 1982 se
rect 5585 1966 5652 1982
tri 5652 1966 5668 1982 nw
tri 8182 1966 8198 1982 se
rect 8198 1966 8244 1982
rect 3186 1920 3852 1953
tri 3994 1944 4016 1966 ne
rect 4016 1944 4068 1966
tri 4068 1944 4090 1966 sw
tri 4114 1944 4136 1966 ne
rect 4136 1944 4612 1966
rect -24 1910 581 1914
rect 353 1873 731 1879
rect 405 1821 679 1873
rect 3186 1868 3211 1920
rect 3263 1868 3775 1920
rect 3827 1868 3852 1920
tri 4016 1914 4046 1944 ne
rect 4046 1920 4090 1944
tri 4090 1920 4114 1944 sw
tri 4136 1920 4160 1944 ne
rect 4160 1920 4612 1944
rect 4046 1914 4114 1920
tri 4114 1914 4120 1920 sw
tri 4160 1914 4166 1920 ne
rect 4166 1914 4612 1920
rect 4664 1914 4676 1966
rect 4728 1939 5625 1966
tri 5625 1939 5652 1966 nw
tri 5814 1939 5841 1966 se
rect 5841 1939 5897 1966
rect 4728 1914 5600 1939
tri 5600 1914 5625 1939 nw
tri 5789 1914 5814 1939 se
rect 5814 1914 5897 1939
rect 5949 1914 5976 1966
rect 6028 1954 6662 1966
tri 6662 1954 6674 1966 sw
tri 8170 1954 8182 1966 se
rect 8182 1954 8244 1966
tri 8244 1954 8272 1982 nw
rect 6028 1948 6674 1954
tri 6674 1948 6680 1954 sw
tri 8164 1948 8170 1954 se
rect 6028 1914 6680 1948
tri 6680 1914 6714 1948 sw
tri 8130 1914 8164 1948 se
rect 8164 1914 8170 1948
tri 4046 1870 4090 1914 ne
rect 4090 1892 4120 1914
tri 4120 1892 4142 1914 sw
tri 5767 1892 5789 1914 se
rect 5789 1892 5841 1914
tri 5841 1892 5863 1914 nw
tri 6640 1892 6662 1914 ne
rect 6662 1892 6714 1914
tri 6714 1892 6736 1914 sw
tri 8108 1892 8130 1914 se
rect 8130 1892 8170 1914
rect 4090 1870 4142 1892
tri 4142 1870 4164 1892 sw
tri 5745 1870 5767 1892 se
rect 5767 1870 5819 1892
tri 5819 1870 5841 1892 nw
tri 6662 1874 6680 1892 ne
rect 6680 1880 6736 1892
tri 6736 1880 6748 1892 sw
tri 8096 1880 8108 1892 se
rect 8108 1880 8170 1892
tri 8170 1880 8244 1954 nw
rect 6680 1874 6748 1880
tri 6748 1874 6754 1880 sw
tri 8090 1874 8096 1880 se
rect 8096 1874 8164 1880
tri 8164 1874 8170 1880 nw
tri 6680 1870 6684 1874 ne
rect 6684 1870 8112 1874
rect 1057 1859 1383 1860
rect 353 1800 731 1821
rect 405 1748 679 1800
rect 353 1726 731 1748
rect 405 1674 679 1726
rect 353 1652 731 1674
rect 405 1600 679 1652
rect 353 1578 731 1600
rect 405 1526 679 1578
rect 353 1504 731 1526
rect 405 1452 679 1504
rect 1005 1853 1383 1859
rect 1057 1801 1331 1853
rect 1005 1775 1383 1801
rect 3186 1835 3852 1868
rect 3186 1783 3211 1835
rect 3263 1783 3775 1835
rect 3827 1783 3852 1835
tri 4090 1818 4142 1870 ne
rect 4142 1818 5767 1870
tri 5767 1818 5819 1870 nw
tri 6684 1822 6732 1870 ne
rect 6732 1822 8112 1870
tri 8112 1822 8164 1874 nw
rect 3186 1777 3852 1783
rect 1057 1723 1331 1775
rect 7088 1732 8259 1738
rect 1005 1696 1383 1723
rect 1057 1644 1331 1696
rect 1005 1617 1383 1644
rect 1057 1565 1331 1617
rect 1005 1538 1383 1565
rect 1057 1486 1331 1538
rect 1005 1480 1383 1486
rect 5386 1717 5764 1723
rect 5438 1665 5712 1717
rect 5386 1638 5764 1665
rect 5438 1586 5712 1638
rect 5386 1559 5764 1586
rect 5438 1507 5712 1559
rect 5386 1480 5764 1507
rect 353 1430 731 1452
rect 405 1378 679 1430
rect 353 1372 731 1378
rect 5438 1428 5712 1480
rect 5386 1401 5764 1428
rect 5438 1349 5712 1401
rect 5386 1343 5764 1349
rect 6038 1717 6416 1723
rect 6090 1665 6364 1717
rect 6038 1638 6416 1665
rect 6090 1586 6364 1638
rect 6038 1559 6416 1586
rect 6090 1507 6364 1559
rect 6038 1480 6416 1507
rect 6090 1428 6364 1480
rect 6038 1401 6416 1428
rect 6090 1349 6364 1401
rect 7140 1680 7370 1732
rect 7422 1680 7696 1732
rect 7748 1680 8022 1732
rect 8074 1723 8259 1732
tri 8259 1723 8274 1738 sw
rect 8074 1680 8274 1723
rect 7088 1661 8274 1680
rect 7140 1609 7370 1661
rect 7422 1609 7696 1661
rect 7748 1609 8022 1661
rect 8074 1609 8274 1661
rect 7088 1590 8274 1609
rect 7140 1538 7370 1590
rect 7422 1538 7696 1590
rect 7748 1538 8022 1590
rect 8074 1538 8274 1590
rect 7088 1518 8274 1538
rect 7140 1466 7370 1518
rect 7422 1466 7696 1518
rect 7748 1466 8022 1518
rect 8074 1504 8274 1518
tri 8274 1504 8493 1723 sw
rect 8074 1466 8493 1504
rect 7088 1446 8493 1466
rect 7140 1394 7370 1446
rect 7422 1394 7696 1446
rect 7748 1394 8022 1446
rect 8074 1394 8493 1446
rect 7088 1388 8493 1394
tri 8493 1388 8609 1504 sw
rect 6038 1343 6416 1349
tri 8234 1343 8279 1388 ne
rect 8279 1343 8609 1388
tri 8279 1232 8390 1343 ne
rect 8390 1232 8609 1343
rect 2230 1226 8237 1232
rect 2230 1174 2237 1226
rect 2289 1174 2563 1226
rect 2615 1174 2889 1226
rect 2941 1174 4285 1226
rect 4337 1174 4611 1226
rect 4663 1174 4937 1226
rect 4989 1174 5263 1226
rect 5315 1174 7207 1226
rect 7259 1174 7533 1226
rect 7585 1174 7859 1226
rect 7911 1174 8185 1226
rect 2230 1157 8237 1174
rect 2230 1105 2237 1157
rect 2289 1105 2563 1157
rect 2615 1105 2889 1157
rect 2941 1105 4285 1157
rect 4337 1105 4611 1157
rect 4663 1105 4937 1157
rect 4989 1105 5263 1157
rect 5315 1105 7207 1157
rect 7259 1105 7533 1157
rect 7585 1105 7859 1157
rect 7911 1105 8185 1157
tri 8390 1129 8493 1232 ne
rect 8493 1154 8609 1232
tri 8609 1154 8843 1388 sw
rect 2230 1088 8237 1105
rect 2230 1036 2237 1088
rect 2289 1036 2563 1088
rect 2615 1036 2889 1088
rect 2941 1036 4285 1088
rect 4337 1036 4611 1088
rect 4663 1036 4937 1088
rect 4989 1036 5263 1088
rect 5315 1036 7207 1088
rect 7259 1036 7533 1088
rect 7585 1036 7859 1088
rect 7911 1036 8185 1088
rect 2230 1019 8237 1036
rect 2230 967 2237 1019
rect 2289 967 2563 1019
rect 2615 967 2889 1019
rect 2941 967 4285 1019
rect 4337 967 4611 1019
rect 4663 967 4937 1019
rect 4989 967 5263 1019
rect 5315 967 7207 1019
rect 7259 967 7533 1019
rect 7585 967 7859 1019
rect 7911 967 8185 1019
rect 2230 950 8237 967
rect 2230 898 2237 950
rect 2289 898 2563 950
rect 2615 898 2889 950
rect 2941 898 4285 950
rect 4337 898 4611 950
rect 4663 898 4937 950
rect 4989 898 5263 950
rect 5315 898 7207 950
rect 7259 898 7533 950
rect 7585 898 7859 950
rect 7911 898 8185 950
rect 2230 892 8237 898
rect 8493 1093 8843 1154
rect 8493 1041 8494 1093
rect 8546 1041 8568 1093
rect 8620 1041 8642 1093
rect 8694 1041 8716 1093
rect 8768 1041 8790 1093
rect 8842 1041 8843 1093
rect 8493 1023 8843 1041
rect 8493 971 8494 1023
rect 8546 971 8568 1023
rect 8620 971 8642 1023
rect 8694 971 8716 1023
rect 8768 971 8790 1023
rect 8842 971 8843 1023
rect 8493 953 8843 971
rect 8493 901 8494 953
rect 8546 901 8568 953
rect 8620 901 8642 953
rect 8694 901 8716 953
rect 8768 901 8790 953
rect 8842 901 8843 953
rect 8493 883 8843 901
rect 8493 831 8494 883
rect 8546 831 8568 883
rect 8620 831 8642 883
rect 8694 831 8716 883
rect 8768 831 8790 883
rect 8842 831 8843 883
rect 8493 813 8843 831
rect 353 803 6698 809
rect 353 751 516 803
rect 568 751 842 803
rect 894 751 1168 803
rect 1220 751 2400 803
rect 2452 751 2726 803
rect 2778 751 3052 803
rect 3104 751 3996 803
rect 4048 751 4122 803
rect 4174 751 4448 803
rect 4500 751 4774 803
rect 4826 751 5100 803
rect 5152 751 5549 803
rect 5601 751 5875 803
rect 5927 751 6201 803
rect 6253 751 6527 803
rect 6579 751 6646 803
rect 353 735 6698 751
rect 353 683 516 735
rect 568 683 842 735
rect 894 683 1168 735
rect 1220 683 2400 735
rect 2452 683 2726 735
rect 2778 683 3052 735
rect 3104 683 3996 735
rect 4048 683 4122 735
rect 4174 683 4448 735
rect 4500 683 4774 735
rect 4826 683 5100 735
rect 5152 683 5549 735
rect 5601 683 5875 735
rect 5927 683 6201 735
rect 6253 683 6527 735
rect 6579 683 6646 735
rect 353 666 6698 683
rect 353 614 516 666
rect 568 614 842 666
rect 894 614 1168 666
rect 1220 614 2400 666
rect 2452 614 2726 666
rect 2778 614 3052 666
rect 3104 614 3996 666
rect 4048 614 4122 666
rect 4174 614 4448 666
rect 4500 614 4774 666
rect 4826 614 5100 666
rect 5152 614 5549 666
rect 5601 614 5875 666
rect 5927 614 6201 666
rect 6253 614 6527 666
rect 6579 614 6646 666
rect 8493 761 8494 813
rect 8546 761 8568 813
rect 8620 761 8642 813
rect 8694 761 8716 813
rect 8768 761 8790 813
rect 8842 761 8843 813
rect 8493 743 8843 761
rect 8493 691 8494 743
rect 8546 691 8568 743
rect 8620 691 8642 743
rect 8694 691 8716 743
rect 8768 691 8790 743
rect 8842 691 8843 743
rect 8493 672 8843 691
rect 8493 620 8494 672
rect 8546 620 8568 672
rect 8620 620 8642 672
rect 8694 620 8716 672
rect 8768 620 8790 672
rect 8842 620 8843 672
rect 8493 614 8843 620
rect 353 597 6698 614
rect 353 545 516 597
rect 568 545 842 597
rect 894 545 1168 597
rect 1220 545 2400 597
rect 2452 545 2726 597
rect 2778 545 3052 597
rect 3104 545 3996 597
rect 4048 545 4122 597
rect 4174 545 4448 597
rect 4500 545 4774 597
rect 4826 545 5100 597
rect 5152 545 5549 597
rect 5601 545 5875 597
rect 5927 545 6201 597
rect 6253 545 6527 597
rect 6579 545 6646 597
rect 353 528 6698 545
rect 353 476 516 528
rect 568 476 842 528
rect 894 476 1168 528
rect 1220 476 2400 528
rect 2452 476 2726 528
rect 2778 476 3052 528
rect 3104 476 3996 528
rect 4048 476 4122 528
rect 4174 476 4448 528
rect 4500 476 4774 528
rect 4826 476 5100 528
rect 5152 476 5549 528
rect 5601 476 5875 528
rect 5927 476 6201 528
rect 6253 476 6527 528
rect 6579 476 6646 528
rect 353 470 6698 476
use sky130_fd_pr__pfet_01v8__example_55959141808564  sky130_fd_pr__pfet_01v8__example_55959141808564_0
timestamp 1624884095
transform -1 0 3043 0 1 475
box -35 0 780 697
use sky130_fd_pr__pfet_01v8__example_55959141808562  sky130_fd_pr__pfet_01v8__example_55959141808562_0
timestamp 1624884095
transform -1 0 1322 0 1 475
box -35 0 943 697
use sky130_fd_pr__nfet_01v8__example_55959141808560  sky130_fd_pr__nfet_01v8__example_55959141808560_0
timestamp 1624884095
transform -1 0 8339 0 1 543
box -35 0 1106 697
use sky130_fd_pr__nfet_01v8__example_55959141808560  sky130_fd_pr__nfet_01v8__example_55959141808560_1
timestamp 1624884095
transform 1 0 5447 0 1 475
box -35 0 1106 697
use sky130_fd_pr__nfet_01v8__example_55959141808560  sky130_fd_pr__nfet_01v8__example_55959141808560_2
timestamp 1624884095
transform -1 0 5254 0 1 475
box -35 0 1106 697
use sky130_fd_pr__nfet_01v8__example_55959141808558  sky130_fd_pr__nfet_01v8__example_55959141808558_0
timestamp 1624884095
transform -1 0 9766 0 1 543
box -35 0 1269 675
<< labels >>
flabel metal2 s 4567 965 5916 1232 3 FreeSans 520 0 0 0 AMUXBUS_HV
port 1 nsew
flabel metal2 s 518 1516 560 1698 3 FreeSans 520 0 0 0 PAD_HV_P0
port 2 nsew
flabel metal2 s -24 2002 97 2040 3 FreeSans 520 0 0 0 PG_AMX_VDDA_H_N
port 3 nsew
flabel metal2 s -24 2168 62 2209 3 FreeSans 520 0 0 0 NG_AMX_VPMP_H
port 4 nsew
flabel metal2 s -24 2081 105 2123 3 FreeSans 520 0 0 0 NG_PAD_VPMP_H
port 5 nsew
flabel metal2 s 1142 1669 1180 1718 3 FreeSans 520 0 0 0 PAD_HV_P1
port 6 nsew
flabel metal2 s -24 1921 117 1960 3 FreeSans 520 0 0 0 PG_PAD_VDDIOQ_H_N
port 7 nsew
flabel metal2 s 5499 1436 5697 1701 3 FreeSans 520 0 0 0 PAD_HV_N0
port 8 nsew
flabel metal2 s 6060 1618 6089 1682 3 FreeSans 520 0 0 0 PAD_HV_N1
port 9 nsew
flabel metal1 s 3168 2300 3222 2333 3 FreeSans 520 0 0 0 VSSD
port 10 nsew
flabel metal1 s 3891 2274 4015 2351 3 FreeSans 520 0 0 0 VDDA
port 11 nsew
flabel metal1 s 8781 1514 8899 1707 3 FreeSans 520 0 0 0 PAD_HV_N2
port 12 nsew
flabel metal1 s 218 1569 254 1648 3 FreeSans 520 0 0 0 VDDIO
port 13 nsew
flabel metal1 s 9421 1760 9451 1800 3 FreeSans 520 0 0 0 PAD_HV_N3
port 14 nsew
flabel comment s 8177 2165 8177 2165 0 FreeSans 440 0 0 0 CONDIODE
flabel comment s 5143 2155 5143 2155 0 FreeSans 440 0 0 0 CONDIODE
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 13625376
string GDS_START 13410064
<< end >>
