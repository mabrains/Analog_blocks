magic
tech sky130A
magscale 1 2
timestamp 1624883981
<< checkpaint >>
rect -1260 -1260 1960 2454
<< pwell >>
rect 0 66 700 1128
<< nmoslvt >>
rect 194 92 230 1102
rect 286 92 322 1102
rect 378 92 414 1102
rect 470 92 506 1102
<< ndiff >>
rect 138 1090 194 1102
rect 138 1056 149 1090
rect 183 1056 194 1090
rect 138 1022 194 1056
rect 138 988 149 1022
rect 183 988 194 1022
rect 138 954 194 988
rect 138 920 149 954
rect 183 920 194 954
rect 138 886 194 920
rect 138 852 149 886
rect 183 852 194 886
rect 138 818 194 852
rect 138 784 149 818
rect 183 784 194 818
rect 138 750 194 784
rect 138 716 149 750
rect 183 716 194 750
rect 138 682 194 716
rect 138 648 149 682
rect 183 648 194 682
rect 138 614 194 648
rect 138 580 149 614
rect 183 580 194 614
rect 138 546 194 580
rect 138 512 149 546
rect 183 512 194 546
rect 138 478 194 512
rect 138 444 149 478
rect 183 444 194 478
rect 138 410 194 444
rect 138 376 149 410
rect 183 376 194 410
rect 138 342 194 376
rect 138 308 149 342
rect 183 308 194 342
rect 138 274 194 308
rect 138 240 149 274
rect 183 240 194 274
rect 138 206 194 240
rect 138 172 149 206
rect 183 172 194 206
rect 138 138 194 172
rect 138 104 149 138
rect 183 104 194 138
rect 138 92 194 104
rect 230 1090 286 1102
rect 230 1056 241 1090
rect 275 1056 286 1090
rect 230 1022 286 1056
rect 230 988 241 1022
rect 275 988 286 1022
rect 230 954 286 988
rect 230 920 241 954
rect 275 920 286 954
rect 230 886 286 920
rect 230 852 241 886
rect 275 852 286 886
rect 230 818 286 852
rect 230 784 241 818
rect 275 784 286 818
rect 230 750 286 784
rect 230 716 241 750
rect 275 716 286 750
rect 230 682 286 716
rect 230 648 241 682
rect 275 648 286 682
rect 230 614 286 648
rect 230 580 241 614
rect 275 580 286 614
rect 230 546 286 580
rect 230 512 241 546
rect 275 512 286 546
rect 230 478 286 512
rect 230 444 241 478
rect 275 444 286 478
rect 230 410 286 444
rect 230 376 241 410
rect 275 376 286 410
rect 230 342 286 376
rect 230 308 241 342
rect 275 308 286 342
rect 230 274 286 308
rect 230 240 241 274
rect 275 240 286 274
rect 230 206 286 240
rect 230 172 241 206
rect 275 172 286 206
rect 230 138 286 172
rect 230 104 241 138
rect 275 104 286 138
rect 230 92 286 104
rect 322 1090 378 1102
rect 322 1056 333 1090
rect 367 1056 378 1090
rect 322 1022 378 1056
rect 322 988 333 1022
rect 367 988 378 1022
rect 322 954 378 988
rect 322 920 333 954
rect 367 920 378 954
rect 322 886 378 920
rect 322 852 333 886
rect 367 852 378 886
rect 322 818 378 852
rect 322 784 333 818
rect 367 784 378 818
rect 322 750 378 784
rect 322 716 333 750
rect 367 716 378 750
rect 322 682 378 716
rect 322 648 333 682
rect 367 648 378 682
rect 322 614 378 648
rect 322 580 333 614
rect 367 580 378 614
rect 322 546 378 580
rect 322 512 333 546
rect 367 512 378 546
rect 322 478 378 512
rect 322 444 333 478
rect 367 444 378 478
rect 322 410 378 444
rect 322 376 333 410
rect 367 376 378 410
rect 322 342 378 376
rect 322 308 333 342
rect 367 308 378 342
rect 322 274 378 308
rect 322 240 333 274
rect 367 240 378 274
rect 322 206 378 240
rect 322 172 333 206
rect 367 172 378 206
rect 322 138 378 172
rect 322 104 333 138
rect 367 104 378 138
rect 322 92 378 104
rect 414 1090 470 1102
rect 414 1056 425 1090
rect 459 1056 470 1090
rect 414 1022 470 1056
rect 414 988 425 1022
rect 459 988 470 1022
rect 414 954 470 988
rect 414 920 425 954
rect 459 920 470 954
rect 414 886 470 920
rect 414 852 425 886
rect 459 852 470 886
rect 414 818 470 852
rect 414 784 425 818
rect 459 784 470 818
rect 414 750 470 784
rect 414 716 425 750
rect 459 716 470 750
rect 414 682 470 716
rect 414 648 425 682
rect 459 648 470 682
rect 414 614 470 648
rect 414 580 425 614
rect 459 580 470 614
rect 414 546 470 580
rect 414 512 425 546
rect 459 512 470 546
rect 414 478 470 512
rect 414 444 425 478
rect 459 444 470 478
rect 414 410 470 444
rect 414 376 425 410
rect 459 376 470 410
rect 414 342 470 376
rect 414 308 425 342
rect 459 308 470 342
rect 414 274 470 308
rect 414 240 425 274
rect 459 240 470 274
rect 414 206 470 240
rect 414 172 425 206
rect 459 172 470 206
rect 414 138 470 172
rect 414 104 425 138
rect 459 104 470 138
rect 414 92 470 104
rect 506 1090 562 1102
rect 506 1056 517 1090
rect 551 1056 562 1090
rect 506 1022 562 1056
rect 506 988 517 1022
rect 551 988 562 1022
rect 506 954 562 988
rect 506 920 517 954
rect 551 920 562 954
rect 506 886 562 920
rect 506 852 517 886
rect 551 852 562 886
rect 506 818 562 852
rect 506 784 517 818
rect 551 784 562 818
rect 506 750 562 784
rect 506 716 517 750
rect 551 716 562 750
rect 506 682 562 716
rect 506 648 517 682
rect 551 648 562 682
rect 506 614 562 648
rect 506 580 517 614
rect 551 580 562 614
rect 506 546 562 580
rect 506 512 517 546
rect 551 512 562 546
rect 506 478 562 512
rect 506 444 517 478
rect 551 444 562 478
rect 506 410 562 444
rect 506 376 517 410
rect 551 376 562 410
rect 506 342 562 376
rect 506 308 517 342
rect 551 308 562 342
rect 506 274 562 308
rect 506 240 517 274
rect 551 240 562 274
rect 506 206 562 240
rect 506 172 517 206
rect 551 172 562 206
rect 506 138 562 172
rect 506 104 517 138
rect 551 104 562 138
rect 506 92 562 104
<< ndiffc >>
rect 149 1056 183 1090
rect 149 988 183 1022
rect 149 920 183 954
rect 149 852 183 886
rect 149 784 183 818
rect 149 716 183 750
rect 149 648 183 682
rect 149 580 183 614
rect 149 512 183 546
rect 149 444 183 478
rect 149 376 183 410
rect 149 308 183 342
rect 149 240 183 274
rect 149 172 183 206
rect 149 104 183 138
rect 241 1056 275 1090
rect 241 988 275 1022
rect 241 920 275 954
rect 241 852 275 886
rect 241 784 275 818
rect 241 716 275 750
rect 241 648 275 682
rect 241 580 275 614
rect 241 512 275 546
rect 241 444 275 478
rect 241 376 275 410
rect 241 308 275 342
rect 241 240 275 274
rect 241 172 275 206
rect 241 104 275 138
rect 333 1056 367 1090
rect 333 988 367 1022
rect 333 920 367 954
rect 333 852 367 886
rect 333 784 367 818
rect 333 716 367 750
rect 333 648 367 682
rect 333 580 367 614
rect 333 512 367 546
rect 333 444 367 478
rect 333 376 367 410
rect 333 308 367 342
rect 333 240 367 274
rect 333 172 367 206
rect 333 104 367 138
rect 425 1056 459 1090
rect 425 988 459 1022
rect 425 920 459 954
rect 425 852 459 886
rect 425 784 459 818
rect 425 716 459 750
rect 425 648 459 682
rect 425 580 459 614
rect 425 512 459 546
rect 425 444 459 478
rect 425 376 459 410
rect 425 308 459 342
rect 425 240 459 274
rect 425 172 459 206
rect 425 104 459 138
rect 517 1056 551 1090
rect 517 988 551 1022
rect 517 920 551 954
rect 517 852 551 886
rect 517 784 551 818
rect 517 716 551 750
rect 517 648 551 682
rect 517 580 551 614
rect 517 512 551 546
rect 517 444 551 478
rect 517 376 551 410
rect 517 308 551 342
rect 517 240 551 274
rect 517 172 551 206
rect 517 104 551 138
<< psubdiff >>
rect 26 1056 84 1102
rect 26 1022 38 1056
rect 72 1022 84 1056
rect 26 988 84 1022
rect 26 954 38 988
rect 72 954 84 988
rect 26 920 84 954
rect 26 886 38 920
rect 72 886 84 920
rect 26 852 84 886
rect 26 818 38 852
rect 72 818 84 852
rect 26 784 84 818
rect 26 750 38 784
rect 72 750 84 784
rect 26 716 84 750
rect 26 682 38 716
rect 72 682 84 716
rect 26 648 84 682
rect 26 614 38 648
rect 72 614 84 648
rect 26 580 84 614
rect 26 546 38 580
rect 72 546 84 580
rect 26 512 84 546
rect 26 478 38 512
rect 72 478 84 512
rect 26 444 84 478
rect 26 410 38 444
rect 72 410 84 444
rect 26 376 84 410
rect 26 342 38 376
rect 72 342 84 376
rect 26 308 84 342
rect 26 274 38 308
rect 72 274 84 308
rect 26 240 84 274
rect 26 206 38 240
rect 72 206 84 240
rect 26 172 84 206
rect 26 138 38 172
rect 72 138 84 172
rect 26 92 84 138
rect 616 1056 674 1102
rect 616 1022 628 1056
rect 662 1022 674 1056
rect 616 988 674 1022
rect 616 954 628 988
rect 662 954 674 988
rect 616 920 674 954
rect 616 886 628 920
rect 662 886 674 920
rect 616 852 674 886
rect 616 818 628 852
rect 662 818 674 852
rect 616 784 674 818
rect 616 750 628 784
rect 662 750 674 784
rect 616 716 674 750
rect 616 682 628 716
rect 662 682 674 716
rect 616 648 674 682
rect 616 614 628 648
rect 662 614 674 648
rect 616 580 674 614
rect 616 546 628 580
rect 662 546 674 580
rect 616 512 674 546
rect 616 478 628 512
rect 662 478 674 512
rect 616 444 674 478
rect 616 410 628 444
rect 662 410 674 444
rect 616 376 674 410
rect 616 342 628 376
rect 662 342 674 376
rect 616 308 674 342
rect 616 274 628 308
rect 662 274 674 308
rect 616 240 674 274
rect 616 206 628 240
rect 662 206 674 240
rect 616 172 674 206
rect 616 138 628 172
rect 662 138 674 172
rect 616 92 674 138
<< psubdiffcont >>
rect 38 1022 72 1056
rect 38 954 72 988
rect 38 886 72 920
rect 38 818 72 852
rect 38 750 72 784
rect 38 682 72 716
rect 38 614 72 648
rect 38 546 72 580
rect 38 478 72 512
rect 38 410 72 444
rect 38 342 72 376
rect 38 274 72 308
rect 38 206 72 240
rect 38 138 72 172
rect 628 1022 662 1056
rect 628 954 662 988
rect 628 886 662 920
rect 628 818 662 852
rect 628 750 662 784
rect 628 682 662 716
rect 628 614 662 648
rect 628 546 662 580
rect 628 478 662 512
rect 628 410 662 444
rect 628 342 662 376
rect 628 274 662 308
rect 628 206 662 240
rect 628 138 662 172
<< poly >>
rect 181 1174 519 1194
rect 181 1140 197 1174
rect 231 1140 265 1174
rect 299 1140 333 1174
rect 367 1140 401 1174
rect 435 1140 469 1174
rect 503 1140 519 1174
rect 181 1124 519 1140
rect 194 1102 230 1124
rect 286 1102 322 1124
rect 378 1102 414 1124
rect 470 1102 506 1124
rect 194 70 230 92
rect 286 70 322 92
rect 378 70 414 92
rect 470 70 506 92
rect 181 54 519 70
rect 181 20 197 54
rect 231 20 265 54
rect 299 20 333 54
rect 367 20 401 54
rect 435 20 469 54
rect 503 20 519 54
rect 181 0 519 20
<< polycont >>
rect 197 1140 231 1174
rect 265 1140 299 1174
rect 333 1140 367 1174
rect 401 1140 435 1174
rect 469 1140 503 1174
rect 197 20 231 54
rect 265 20 299 54
rect 333 20 367 54
rect 401 20 435 54
rect 469 20 503 54
<< locali >>
rect 181 1140 189 1174
rect 231 1140 261 1174
rect 299 1140 333 1174
rect 367 1140 401 1174
rect 439 1140 469 1174
rect 511 1140 519 1174
rect 149 1090 183 1106
rect 38 1010 72 1022
rect 38 938 72 954
rect 38 866 72 886
rect 38 794 72 818
rect 38 722 72 750
rect 38 650 72 682
rect 38 580 72 614
rect 38 512 72 544
rect 38 444 72 472
rect 38 376 72 400
rect 38 308 72 328
rect 38 240 72 256
rect 38 172 72 184
rect 149 1022 183 1048
rect 149 954 183 976
rect 149 886 183 904
rect 149 818 183 832
rect 149 750 183 760
rect 149 682 183 688
rect 149 614 183 616
rect 149 578 183 580
rect 149 506 183 512
rect 149 434 183 444
rect 149 362 183 376
rect 149 290 183 308
rect 149 218 183 240
rect 149 146 183 172
rect 149 88 183 104
rect 241 1090 275 1106
rect 241 1022 275 1048
rect 241 954 275 976
rect 241 886 275 904
rect 241 818 275 832
rect 241 750 275 760
rect 241 682 275 688
rect 241 614 275 616
rect 241 578 275 580
rect 241 506 275 512
rect 241 434 275 444
rect 241 362 275 376
rect 241 290 275 308
rect 241 218 275 240
rect 241 146 275 172
rect 241 88 275 104
rect 333 1090 367 1106
rect 333 1022 367 1048
rect 333 954 367 976
rect 333 886 367 904
rect 333 818 367 832
rect 333 750 367 760
rect 333 682 367 688
rect 333 614 367 616
rect 333 578 367 580
rect 333 506 367 512
rect 333 434 367 444
rect 333 362 367 376
rect 333 290 367 308
rect 333 218 367 240
rect 333 146 367 172
rect 333 88 367 104
rect 425 1090 459 1106
rect 425 1022 459 1048
rect 425 954 459 976
rect 425 886 459 904
rect 425 818 459 832
rect 425 750 459 760
rect 425 682 459 688
rect 425 614 459 616
rect 425 578 459 580
rect 425 506 459 512
rect 425 434 459 444
rect 425 362 459 376
rect 425 290 459 308
rect 425 218 459 240
rect 425 146 459 172
rect 425 88 459 104
rect 517 1090 551 1106
rect 517 1022 551 1048
rect 517 954 551 976
rect 517 886 551 904
rect 517 818 551 832
rect 517 750 551 760
rect 517 682 551 688
rect 517 614 551 616
rect 517 578 551 580
rect 517 506 551 512
rect 517 434 551 444
rect 517 362 551 376
rect 517 290 551 308
rect 517 218 551 240
rect 517 146 551 172
rect 628 1010 662 1022
rect 628 938 662 954
rect 628 866 662 886
rect 628 794 662 818
rect 628 722 662 750
rect 628 650 662 682
rect 628 580 662 614
rect 628 512 662 544
rect 628 444 662 472
rect 628 376 662 400
rect 628 308 662 328
rect 628 240 662 256
rect 628 172 662 184
rect 517 88 551 104
rect 181 20 189 54
rect 231 20 261 54
rect 299 20 333 54
rect 367 20 401 54
rect 439 20 469 54
rect 511 20 519 54
<< viali >>
rect 189 1140 197 1174
rect 197 1140 223 1174
rect 261 1140 265 1174
rect 265 1140 295 1174
rect 333 1140 367 1174
rect 405 1140 435 1174
rect 435 1140 439 1174
rect 477 1140 503 1174
rect 503 1140 511 1174
rect 38 1056 72 1082
rect 38 1048 72 1056
rect 38 988 72 1010
rect 38 976 72 988
rect 38 920 72 938
rect 38 904 72 920
rect 38 852 72 866
rect 38 832 72 852
rect 38 784 72 794
rect 38 760 72 784
rect 38 716 72 722
rect 38 688 72 716
rect 38 648 72 650
rect 38 616 72 648
rect 38 546 72 578
rect 38 544 72 546
rect 38 478 72 506
rect 38 472 72 478
rect 38 410 72 434
rect 38 400 72 410
rect 38 342 72 362
rect 38 328 72 342
rect 38 274 72 290
rect 38 256 72 274
rect 38 206 72 218
rect 38 184 72 206
rect 38 138 72 146
rect 38 112 72 138
rect 149 1056 183 1082
rect 149 1048 183 1056
rect 149 988 183 1010
rect 149 976 183 988
rect 149 920 183 938
rect 149 904 183 920
rect 149 852 183 866
rect 149 832 183 852
rect 149 784 183 794
rect 149 760 183 784
rect 149 716 183 722
rect 149 688 183 716
rect 149 648 183 650
rect 149 616 183 648
rect 149 546 183 578
rect 149 544 183 546
rect 149 478 183 506
rect 149 472 183 478
rect 149 410 183 434
rect 149 400 183 410
rect 149 342 183 362
rect 149 328 183 342
rect 149 274 183 290
rect 149 256 183 274
rect 149 206 183 218
rect 149 184 183 206
rect 149 138 183 146
rect 149 112 183 138
rect 241 1056 275 1082
rect 241 1048 275 1056
rect 241 988 275 1010
rect 241 976 275 988
rect 241 920 275 938
rect 241 904 275 920
rect 241 852 275 866
rect 241 832 275 852
rect 241 784 275 794
rect 241 760 275 784
rect 241 716 275 722
rect 241 688 275 716
rect 241 648 275 650
rect 241 616 275 648
rect 241 546 275 578
rect 241 544 275 546
rect 241 478 275 506
rect 241 472 275 478
rect 241 410 275 434
rect 241 400 275 410
rect 241 342 275 362
rect 241 328 275 342
rect 241 274 275 290
rect 241 256 275 274
rect 241 206 275 218
rect 241 184 275 206
rect 241 138 275 146
rect 241 112 275 138
rect 333 1056 367 1082
rect 333 1048 367 1056
rect 333 988 367 1010
rect 333 976 367 988
rect 333 920 367 938
rect 333 904 367 920
rect 333 852 367 866
rect 333 832 367 852
rect 333 784 367 794
rect 333 760 367 784
rect 333 716 367 722
rect 333 688 367 716
rect 333 648 367 650
rect 333 616 367 648
rect 333 546 367 578
rect 333 544 367 546
rect 333 478 367 506
rect 333 472 367 478
rect 333 410 367 434
rect 333 400 367 410
rect 333 342 367 362
rect 333 328 367 342
rect 333 274 367 290
rect 333 256 367 274
rect 333 206 367 218
rect 333 184 367 206
rect 333 138 367 146
rect 333 112 367 138
rect 425 1056 459 1082
rect 425 1048 459 1056
rect 425 988 459 1010
rect 425 976 459 988
rect 425 920 459 938
rect 425 904 459 920
rect 425 852 459 866
rect 425 832 459 852
rect 425 784 459 794
rect 425 760 459 784
rect 425 716 459 722
rect 425 688 459 716
rect 425 648 459 650
rect 425 616 459 648
rect 425 546 459 578
rect 425 544 459 546
rect 425 478 459 506
rect 425 472 459 478
rect 425 410 459 434
rect 425 400 459 410
rect 425 342 459 362
rect 425 328 459 342
rect 425 274 459 290
rect 425 256 459 274
rect 425 206 459 218
rect 425 184 459 206
rect 425 138 459 146
rect 425 112 459 138
rect 517 1056 551 1082
rect 517 1048 551 1056
rect 517 988 551 1010
rect 517 976 551 988
rect 517 920 551 938
rect 517 904 551 920
rect 517 852 551 866
rect 517 832 551 852
rect 517 784 551 794
rect 517 760 551 784
rect 517 716 551 722
rect 517 688 551 716
rect 517 648 551 650
rect 517 616 551 648
rect 517 546 551 578
rect 517 544 551 546
rect 517 478 551 506
rect 517 472 551 478
rect 517 410 551 434
rect 517 400 551 410
rect 517 342 551 362
rect 517 328 551 342
rect 517 274 551 290
rect 517 256 551 274
rect 517 206 551 218
rect 517 184 551 206
rect 517 138 551 146
rect 517 112 551 138
rect 628 1056 662 1082
rect 628 1048 662 1056
rect 628 988 662 1010
rect 628 976 662 988
rect 628 920 662 938
rect 628 904 662 920
rect 628 852 662 866
rect 628 832 662 852
rect 628 784 662 794
rect 628 760 662 784
rect 628 716 662 722
rect 628 688 662 716
rect 628 648 662 650
rect 628 616 662 648
rect 628 546 662 578
rect 628 544 662 546
rect 628 478 662 506
rect 628 472 662 478
rect 628 410 662 434
rect 628 400 662 410
rect 628 342 662 362
rect 628 328 662 342
rect 628 274 662 290
rect 628 256 662 274
rect 628 206 662 218
rect 628 184 662 206
rect 628 138 662 146
rect 628 112 662 138
rect 189 20 197 54
rect 197 20 223 54
rect 261 20 265 54
rect 265 20 295 54
rect 333 20 367 54
rect 405 20 435 54
rect 435 20 439 54
rect 477 20 503 54
rect 503 20 511 54
<< metal1 >>
rect 177 1174 523 1194
rect 177 1140 189 1174
rect 223 1140 261 1174
rect 295 1140 333 1174
rect 367 1140 405 1174
rect 439 1140 477 1174
rect 511 1140 523 1174
rect 177 1128 523 1140
rect 26 1082 84 1094
rect 26 1048 38 1082
rect 72 1048 84 1082
rect 26 1010 84 1048
rect 26 976 38 1010
rect 72 976 84 1010
rect 26 938 84 976
rect 26 904 38 938
rect 72 904 84 938
rect 26 866 84 904
rect 26 832 38 866
rect 72 832 84 866
rect 26 794 84 832
rect 26 760 38 794
rect 72 760 84 794
rect 26 722 84 760
rect 26 688 38 722
rect 72 688 84 722
rect 26 650 84 688
rect 26 616 38 650
rect 72 616 84 650
rect 26 578 84 616
rect 26 544 38 578
rect 72 544 84 578
rect 26 506 84 544
rect 26 472 38 506
rect 72 472 84 506
rect 26 434 84 472
rect 26 400 38 434
rect 72 400 84 434
rect 26 362 84 400
rect 26 328 38 362
rect 72 328 84 362
rect 26 290 84 328
rect 26 256 38 290
rect 72 256 84 290
rect 26 218 84 256
rect 26 184 38 218
rect 72 184 84 218
rect 26 146 84 184
rect 26 112 38 146
rect 72 112 84 146
rect 26 100 84 112
rect 140 1082 192 1094
rect 140 1048 149 1082
rect 183 1048 192 1082
rect 140 1010 192 1048
rect 140 976 149 1010
rect 183 976 192 1010
rect 140 938 192 976
rect 140 904 149 938
rect 183 904 192 938
rect 140 866 192 904
rect 140 832 149 866
rect 183 832 192 866
rect 140 794 192 832
rect 140 760 149 794
rect 183 760 192 794
rect 140 722 192 760
rect 140 688 149 722
rect 183 688 192 722
rect 140 650 192 688
rect 140 616 149 650
rect 183 616 192 650
rect 140 578 192 616
rect 140 544 149 578
rect 183 544 192 578
rect 140 542 192 544
rect 140 478 149 490
rect 183 478 192 490
rect 140 414 149 426
rect 183 414 192 426
rect 140 350 149 362
rect 183 350 192 362
rect 140 290 192 298
rect 140 286 149 290
rect 183 286 192 290
rect 140 222 192 234
rect 140 158 192 170
rect 140 100 192 106
rect 232 1088 284 1094
rect 232 1024 284 1036
rect 232 960 284 972
rect 232 904 241 908
rect 275 904 284 908
rect 232 896 284 904
rect 232 832 241 844
rect 275 832 284 844
rect 232 768 241 780
rect 275 768 284 780
rect 232 704 241 716
rect 275 704 284 716
rect 232 650 284 652
rect 232 616 241 650
rect 275 616 284 650
rect 232 578 284 616
rect 232 544 241 578
rect 275 544 284 578
rect 232 506 284 544
rect 232 472 241 506
rect 275 472 284 506
rect 232 434 284 472
rect 232 400 241 434
rect 275 400 284 434
rect 232 362 284 400
rect 232 328 241 362
rect 275 328 284 362
rect 232 290 284 328
rect 232 256 241 290
rect 275 256 284 290
rect 232 218 284 256
rect 232 184 241 218
rect 275 184 284 218
rect 232 146 284 184
rect 232 112 241 146
rect 275 112 284 146
rect 232 100 284 112
rect 324 1082 376 1094
rect 324 1048 333 1082
rect 367 1048 376 1082
rect 324 1010 376 1048
rect 324 976 333 1010
rect 367 976 376 1010
rect 324 938 376 976
rect 324 904 333 938
rect 367 904 376 938
rect 324 866 376 904
rect 324 832 333 866
rect 367 832 376 866
rect 324 794 376 832
rect 324 760 333 794
rect 367 760 376 794
rect 324 722 376 760
rect 324 688 333 722
rect 367 688 376 722
rect 324 650 376 688
rect 324 616 333 650
rect 367 616 376 650
rect 324 578 376 616
rect 324 544 333 578
rect 367 544 376 578
rect 324 542 376 544
rect 324 478 333 490
rect 367 478 376 490
rect 324 414 333 426
rect 367 414 376 426
rect 324 350 333 362
rect 367 350 376 362
rect 324 290 376 298
rect 324 286 333 290
rect 367 286 376 290
rect 324 222 376 234
rect 324 158 376 170
rect 324 100 376 106
rect 416 1088 468 1094
rect 416 1024 468 1036
rect 416 960 468 972
rect 416 904 425 908
rect 459 904 468 908
rect 416 896 468 904
rect 416 832 425 844
rect 459 832 468 844
rect 416 768 425 780
rect 459 768 468 780
rect 416 704 425 716
rect 459 704 468 716
rect 416 650 468 652
rect 416 616 425 650
rect 459 616 468 650
rect 416 578 468 616
rect 416 544 425 578
rect 459 544 468 578
rect 416 506 468 544
rect 416 472 425 506
rect 459 472 468 506
rect 416 434 468 472
rect 416 400 425 434
rect 459 400 468 434
rect 416 362 468 400
rect 416 328 425 362
rect 459 328 468 362
rect 416 290 468 328
rect 416 256 425 290
rect 459 256 468 290
rect 416 218 468 256
rect 416 184 425 218
rect 459 184 468 218
rect 416 146 468 184
rect 416 112 425 146
rect 459 112 468 146
rect 416 100 468 112
rect 508 1082 560 1094
rect 508 1048 517 1082
rect 551 1048 560 1082
rect 508 1010 560 1048
rect 508 976 517 1010
rect 551 976 560 1010
rect 508 938 560 976
rect 508 904 517 938
rect 551 904 560 938
rect 508 866 560 904
rect 508 832 517 866
rect 551 832 560 866
rect 508 794 560 832
rect 508 760 517 794
rect 551 760 560 794
rect 508 722 560 760
rect 508 688 517 722
rect 551 688 560 722
rect 508 650 560 688
rect 508 616 517 650
rect 551 616 560 650
rect 508 578 560 616
rect 508 544 517 578
rect 551 544 560 578
rect 508 542 560 544
rect 508 478 517 490
rect 551 478 560 490
rect 508 414 517 426
rect 551 414 560 426
rect 508 350 517 362
rect 551 350 560 362
rect 508 290 560 298
rect 508 286 517 290
rect 551 286 560 290
rect 508 222 560 234
rect 508 158 560 170
rect 508 100 560 106
rect 616 1082 674 1094
rect 616 1048 628 1082
rect 662 1048 674 1082
rect 616 1010 674 1048
rect 616 976 628 1010
rect 662 976 674 1010
rect 616 938 674 976
rect 616 904 628 938
rect 662 904 674 938
rect 616 866 674 904
rect 616 832 628 866
rect 662 832 674 866
rect 616 794 674 832
rect 616 760 628 794
rect 662 760 674 794
rect 616 722 674 760
rect 616 688 628 722
rect 662 688 674 722
rect 616 650 674 688
rect 616 616 628 650
rect 662 616 674 650
rect 616 578 674 616
rect 616 544 628 578
rect 662 544 674 578
rect 616 506 674 544
rect 616 472 628 506
rect 662 472 674 506
rect 616 434 674 472
rect 616 400 628 434
rect 662 400 674 434
rect 616 362 674 400
rect 616 328 628 362
rect 662 328 674 362
rect 616 290 674 328
rect 616 256 628 290
rect 662 256 674 290
rect 616 218 674 256
rect 616 184 628 218
rect 662 184 674 218
rect 616 146 674 184
rect 616 112 628 146
rect 662 112 674 146
rect 616 100 674 112
rect 177 54 523 66
rect 177 20 189 54
rect 223 20 261 54
rect 295 20 333 54
rect 367 20 405 54
rect 439 20 477 54
rect 511 20 523 54
rect 177 0 523 20
<< via1 >>
rect 140 506 192 542
rect 140 490 149 506
rect 149 490 183 506
rect 183 490 192 506
rect 140 472 149 478
rect 149 472 183 478
rect 183 472 192 478
rect 140 434 192 472
rect 140 426 149 434
rect 149 426 183 434
rect 183 426 192 434
rect 140 400 149 414
rect 149 400 183 414
rect 183 400 192 414
rect 140 362 192 400
rect 140 328 149 350
rect 149 328 183 350
rect 183 328 192 350
rect 140 298 192 328
rect 140 256 149 286
rect 149 256 183 286
rect 183 256 192 286
rect 140 234 192 256
rect 140 218 192 222
rect 140 184 149 218
rect 149 184 183 218
rect 183 184 192 218
rect 140 170 192 184
rect 140 146 192 158
rect 140 112 149 146
rect 149 112 183 146
rect 183 112 192 146
rect 140 106 192 112
rect 232 1082 284 1088
rect 232 1048 241 1082
rect 241 1048 275 1082
rect 275 1048 284 1082
rect 232 1036 284 1048
rect 232 1010 284 1024
rect 232 976 241 1010
rect 241 976 275 1010
rect 275 976 284 1010
rect 232 972 284 976
rect 232 938 284 960
rect 232 908 241 938
rect 241 908 275 938
rect 275 908 284 938
rect 232 866 284 896
rect 232 844 241 866
rect 241 844 275 866
rect 275 844 284 866
rect 232 794 284 832
rect 232 780 241 794
rect 241 780 275 794
rect 275 780 284 794
rect 232 760 241 768
rect 241 760 275 768
rect 275 760 284 768
rect 232 722 284 760
rect 232 716 241 722
rect 241 716 275 722
rect 275 716 284 722
rect 232 688 241 704
rect 241 688 275 704
rect 275 688 284 704
rect 232 652 284 688
rect 324 506 376 542
rect 324 490 333 506
rect 333 490 367 506
rect 367 490 376 506
rect 324 472 333 478
rect 333 472 367 478
rect 367 472 376 478
rect 324 434 376 472
rect 324 426 333 434
rect 333 426 367 434
rect 367 426 376 434
rect 324 400 333 414
rect 333 400 367 414
rect 367 400 376 414
rect 324 362 376 400
rect 324 328 333 350
rect 333 328 367 350
rect 367 328 376 350
rect 324 298 376 328
rect 324 256 333 286
rect 333 256 367 286
rect 367 256 376 286
rect 324 234 376 256
rect 324 218 376 222
rect 324 184 333 218
rect 333 184 367 218
rect 367 184 376 218
rect 324 170 376 184
rect 324 146 376 158
rect 324 112 333 146
rect 333 112 367 146
rect 367 112 376 146
rect 324 106 376 112
rect 416 1082 468 1088
rect 416 1048 425 1082
rect 425 1048 459 1082
rect 459 1048 468 1082
rect 416 1036 468 1048
rect 416 1010 468 1024
rect 416 976 425 1010
rect 425 976 459 1010
rect 459 976 468 1010
rect 416 972 468 976
rect 416 938 468 960
rect 416 908 425 938
rect 425 908 459 938
rect 459 908 468 938
rect 416 866 468 896
rect 416 844 425 866
rect 425 844 459 866
rect 459 844 468 866
rect 416 794 468 832
rect 416 780 425 794
rect 425 780 459 794
rect 459 780 468 794
rect 416 760 425 768
rect 425 760 459 768
rect 459 760 468 768
rect 416 722 468 760
rect 416 716 425 722
rect 425 716 459 722
rect 459 716 468 722
rect 416 688 425 704
rect 425 688 459 704
rect 459 688 468 704
rect 416 652 468 688
rect 508 506 560 542
rect 508 490 517 506
rect 517 490 551 506
rect 551 490 560 506
rect 508 472 517 478
rect 517 472 551 478
rect 551 472 560 478
rect 508 434 560 472
rect 508 426 517 434
rect 517 426 551 434
rect 551 426 560 434
rect 508 400 517 414
rect 517 400 551 414
rect 551 400 560 414
rect 508 362 560 400
rect 508 328 517 350
rect 517 328 551 350
rect 551 328 560 350
rect 508 298 560 328
rect 508 256 517 286
rect 517 256 551 286
rect 551 256 560 286
rect 508 234 560 256
rect 508 218 560 222
rect 508 184 517 218
rect 517 184 551 218
rect 551 184 560 218
rect 508 170 560 184
rect 508 146 560 158
rect 508 112 517 146
rect 517 112 551 146
rect 551 112 560 146
rect 508 106 560 112
<< metal2 >>
rect 0 1088 700 1094
rect 0 1036 232 1088
rect 284 1036 416 1088
rect 468 1036 700 1088
rect 0 1024 700 1036
rect 0 972 232 1024
rect 284 972 416 1024
rect 468 972 700 1024
rect 0 960 700 972
rect 0 908 232 960
rect 284 908 416 960
rect 468 908 700 960
rect 0 896 700 908
rect 0 844 232 896
rect 284 844 416 896
rect 468 844 700 896
rect 0 832 700 844
rect 0 780 232 832
rect 284 780 416 832
rect 468 780 700 832
rect 0 768 700 780
rect 0 716 232 768
rect 284 716 416 768
rect 468 716 700 768
rect 0 704 700 716
rect 0 652 232 704
rect 284 652 416 704
rect 468 652 700 704
rect 0 622 700 652
rect 0 542 700 572
rect 0 490 140 542
rect 192 490 324 542
rect 376 490 508 542
rect 560 490 700 542
rect 0 478 700 490
rect 0 426 140 478
rect 192 426 324 478
rect 376 426 508 478
rect 560 426 700 478
rect 0 414 700 426
rect 0 362 140 414
rect 192 362 324 414
rect 376 362 508 414
rect 560 362 700 414
rect 0 350 700 362
rect 0 298 140 350
rect 192 298 324 350
rect 376 298 508 350
rect 560 298 700 350
rect 0 286 700 298
rect 0 234 140 286
rect 192 234 324 286
rect 376 234 508 286
rect 560 234 700 286
rect 0 222 700 234
rect 0 170 140 222
rect 192 170 324 222
rect 376 170 508 222
rect 560 170 700 222
rect 0 158 700 170
rect 0 106 140 158
rect 192 106 324 158
rect 376 106 508 158
rect 560 106 700 158
rect 0 100 700 106
<< labels >>
flabel comment s 350 597 350 597 0 FreeSans 300 0 0 0 S
flabel comment s 350 597 350 597 0 FreeSans 300 0 0 0 S
flabel comment s 442 597 442 597 0 FreeSans 300 0 0 0 S
flabel comment s 442 597 442 597 0 FreeSans 300 0 0 0 D
flabel comment s 534 597 534 597 0 FreeSans 300 0 0 0 S
flabel comment s 166 597 166 597 0 FreeSans 300 0 0 0 S
flabel comment s 166 597 166 597 0 FreeSans 300 0 0 0 S
flabel comment s 258 597 258 597 0 FreeSans 300 0 0 0 D
flabel comment s 258 597 258 597 0 FreeSans 300 0 0 0 S
flabel metal1 s 637 674 637 674 7 FreeSans 300 90 0 0 SUBSTRATE
port 4 nsew
flabel metal1 s 309 23 391 48 0 FreeSans 300 0 0 0 GATE
port 2 nsew
flabel metal1 s 310 1144 392 1169 0 FreeSans 300 0 0 0 GATE
port 2 nsew
flabel metal1 s 51 711 51 711 7 FreeSans 300 90 0 0 SUBSTRATE
port 4 nsew
flabel metal2 s 4 817 22 887 0 FreeSans 300 90 0 0 DRAIN
port 1 nsew
flabel metal2 s 3 312 23 376 0 FreeSans 300 90 0 0 SOURCE
port 3 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 6149770
string GDS_START 6127680
<< end >>
