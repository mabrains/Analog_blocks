**.subckt Pass_transistor_TB
XM1 Vout net2 Vin Vin sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1400 m=1400 
R1 Vout net1 50k m=1
R2 net1 0 100k m=1
E1 net2 0 net1 Vref 1e6
I0 Vout 0 50m
XM2 Vout2 net4 Vin2 Vin2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=20 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1400 m=1400 
R3 Vout2 net3 50k m=1
R4 net3 0 100k m=1
I1 Vout2 0 50m
x1 net3 net4 Vref2 Ideal_opamp
**** begin user architecture code


.option wnflag=1
.option savecurrents
**.subckt test_bsource PLUS MINUS OUT
*.ipin PLUS
*.ipin MINUS
*.opin OUT
.param VDD=3.6
.param GAIN={1000/VDD*2}
VVin Vin 0 2
VVin2 Vin2 0 2
VVref Vref 0 1.2
VVref2 Vref2 0 1.2
.control
save all
save @m.xm1.msky130_fd_pr__pfet_g5v0d10v5[vds]
save @m.xm1.msky130_fd_pr__pfet_g5v0d10v5[vdsat]
save @m.xm1.msky130_fd_pr__pfet_g5v0d10v5[vgs]
save @m.xm1.msky130_fd_pr__pfet_g5v0d10v5[vth]
save @m.xm2.msky130_fd_pr__pfet_g5v0d10v5[vds]
save @m.xm2.msky130_fd_pr__pfet_g5v0d10v5[vdsat]
save @m.xm2.msky130_fd_pr__pfet_g5v0d10v5[vgs]
save @m.xm2.msky130_fd_pr__pfet_g5v0d10v5[vth]
op
show
write Pass_transistor_TB.raw
.endc




.param mc_mm_switch=0
.param mc_pr_switch=0
.include ~/mabrains/Analog_blocks/models/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_01v8__sf.corner.spice
.include ~/mabrains/Analog_blocks/models/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_01v8_lvt__sf.corner.spice
.include ~/mabrains/Analog_blocks/models/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__pfet_01v8__sf.corner.spice
.include ~/mabrains/Analog_blocks/models/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_03v3_nvt__sf.corner.spice
.include ~/mabrains/Analog_blocks/models/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_05v0_nvt__sf.corner.spice
.include ~/mabrains/Analog_blocks/models/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__esd_nfet_01v8__sf.corner.spice
.include ~/mabrains/Analog_blocks/models/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__pfet_01v8_lvt__sf.corner.spice
.include ~/mabrains/Analog_blocks/models/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__pfet_01v8_hvt__sf.corner.spice
.include ~/mabrains/Analog_blocks/models/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__esd_pfet_g5v0d10v5__sf.corner.spice
.include ~/mabrains/Analog_blocks/models/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__pfet_g5v0d10v5__sf.corner.spice
.include ~/mabrains/Analog_blocks/models/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__pfet_g5v0d16v0__sf.corner.spice
.include ~/mabrains/Analog_blocks/models/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_g5v0d10v5__sf.corner.spice
.include ~/mabrains/Analog_blocks/models/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_g5v0d16v0__sf_discrete.corner.spice
.include ~/mabrains/Analog_blocks/models/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__esd_nfet_g5v0d10v5__sf.corner.spice
.include ~/mabrains/Analog_blocks/models/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__pfet_20v0__sf_discrete.corner.spice
.include ~/mabrains/Analog_blocks/models/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_20v0__sf_discrete.corner.spice
.include ~/mabrains/Analog_blocks/models/sky130A/libs.tech/ngspice/corners/sf/nonfet.spice
* Mismatch parameters
.include ~/mabrains/Analog_blocks/models/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_01v8__mismatch.corner.spice
.include ~/mabrains/Analog_blocks/models/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__pfet_01v8__mismatch.corner.spice
.include ~/mabrains/Analog_blocks/models/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_01v8_lvt__mismatch.corner.spice
.include ~/mabrains/Analog_blocks/models/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__pfet_01v8_lvt__mismatch.corner.spice
.include ~/mabrains/Analog_blocks/models/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__pfet_01v8_hvt__mismatch.corner.spice
.include ~/mabrains/Analog_blocks/models/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_g5v0d10v5__mismatch.corner.spice
.include ~/mabrains/Analog_blocks/models/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__pfet_g5v0d10v5__mismatch.corner.spice
.include ~/mabrains/Analog_blocks/models/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_05v0_nvt__mismatch.corner.spice
.include ~/mabrains/Analog_blocks/models/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_03v3_nvt__mismatch.corner.spice
* Resistor/Capacitor
.include ~/mabrains/Analog_blocks/models/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include ~/mabrains/Analog_blocks/models/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
* Special cells
.include ~/mabrains/Analog_blocks/models/sky130A/libs.tech/ngspice/corners/sf/specialized_cells.spice
* All models
.include ~/mabrains/Analog_blocks/models/sky130A/libs.tech/ngspice/all.spice
* Corner
.include ~/mabrains/Analog_blocks/models/sky130A/libs.tech/ngspice/corners/sf/rf.spice



**** end user architecture code
**.ends

* expanding   symbol:
*+  /home/eslam/mabrains/Analog_blocks/Analog_Blocks/OTA/Schematic/Ideal_opamp/Ideal_opamp.sym # of pins=3
* sym_path:
*+ /home/eslam/mabrains/Analog_blocks/Analog_Blocks/OTA/Schematic/Ideal_opamp/Ideal_opamp.sym
* sch_path:
*+ /home/eslam/mabrains/Analog_blocks/Analog_Blocks/OTA/Schematic/Ideal_opamp/Ideal_opamp.sch
.subckt Ideal_opamp  Vp Out Vn
*.ipin Vp
*.ipin Vn
*.opin Out
V1 Vp PLUS_I 0
V2 Vn MINUS_I 0
B1 Out 0 V = 'VDD/2*(1+tanh(GAIN*(V(PLUS_I)-V(MINUS_I))))' 
.ends

** flattened .save nodes
.end
