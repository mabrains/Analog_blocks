* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre = 0.0
.param sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre = 0.0
.param sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre = 0.0
.param sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre = 0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__pfet_g5v0d10v5__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_g5v0d10v5__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_g5v0d10v5__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt  sky130_fd_pr__pfet_g5v0d10v5 d g s b
+ 
.param  l = 1 w = 1 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1 
msky130_fd_pr__pfet_g5v0d10v5 d g s b sky130_fd_pr__pfet_g5v0d10v5__model l = {l} w = {w} nf = {nf} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd} 
.model sky130_fd_pr__pfet_g5v0d10v5__model.0 pmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 9.995e-06 wmax = 1.0005e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.981+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_0+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.59804
+ k2 = {0.024041+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_0}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {68340+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_0}
+ ua = {2.1590772e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_0}
+ ub = {8.2164e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_0}
+ uc = -5.2815e-12
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_0}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.021377+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_0}
+ a0 = {0.95964+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_0}
+ keta = {-0.08587+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_0}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {1.25+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_0}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_0}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_0}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.10153677+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_0+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.1999+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_0+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_0}
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.064044+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_0}
+ etab = -0.0073156
+ dsub = 0.27967
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {1.2297+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_0}
+ pdiblc1 = 0.29403034
+ pdiblc2 = 0.0048008826
+ pdiblcb = -0.025
+ drout = 0.89960455
+ pscbe1 = 3.6263996e+8
+ pscbe2 = 1.448673e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 9.713535e-5
+ alpha1 = 0.0
+ beta0 = 54.684511
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_0}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_0}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {7.5e-009+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_0}
+ bgidl = {1.5572e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_0}
+ cgidl = {264.48+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_0}
+ egidl = 0.66526877
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.60348+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_0}
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.3724
+ ua1 = 5.52e-10
+ ub1 = -2.16e-18
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.1 pmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 1.4995e-05 wmax = 1.5005e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.9724+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_1+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.57939
+ k2 = {0.020277+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_1}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {47889+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_1}
+ ua = {1.6494295e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_1}
+ ub = {1.0975e-018+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_1}
+ uc = -5.8546e-13
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_1}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.020384+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_1}
+ a0 = {0.85515+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_1}
+ keta = {-0.084672+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_1}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.77943+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_1}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_1}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_1}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.077755783+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_1+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.3116+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_1+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_1}
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {4.2119e-005+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_1}
+ etab = 0.0
+ dsub = 0.54416
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {1.2031+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_1}
+ pdiblc1 = 0.3995264
+ pdiblc2 = 0.0015061847
+ pdiblcb = -0.025
+ drout = 0.41068941
+ pscbe1 = 2.994803e+8
+ pscbe2 = 1.4554569e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 6.7813161e-5
+ alpha1 = 0.0
+ beta0 = 50.152925
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_1}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_1}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {8.3464e-009+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_1}
+ bgidl = {1.6889e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_1}
+ cgidl = {368+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_1}
+ egidl = 0.77897916
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.6412+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_1}
+ kt2 = -0.019032
+ at = 31800.0
+ ute = -1.6069
+ ua1 = 4.1982e-10
+ ub1 = -3.8064e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.2 pmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 1.4995e-05 wmax = 1.5005e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.9885+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_2+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.59804
+ k2 = {0.024041+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_2}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {67000+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_2}
+ ua = {2.1590772e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_2}
+ ub = {9.5539e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_2}
+ uc = -5.2815e-12
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_2}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.022+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_2}
+ a0 = {0.95964+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_2}
+ keta = {-0.08587+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_2}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {1.25+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_2}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_2}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_2}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.10153677+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_2+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.1999+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_2+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_2}
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.068847+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_2}
+ etab = -0.0038503
+ dsub = 0.27967
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {1.3366+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_2}
+ pdiblc1 = 0.29403034
+ pdiblc2 = 0.0048008826
+ pdiblcb = -0.025
+ drout = 0.89960455
+ pscbe1 = 3.6263996e+8
+ pscbe2 = 1.448673e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 9.713535e-5
+ alpha1 = 0.0
+ beta0 = 54.684511
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_2}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_2}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.3668e-008+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_2}
+ bgidl = {1.6195e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_2}
+ cgidl = {316.68+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_2}
+ egidl = 0.66526877
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.60348+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_2}
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.3724
+ ua1 = 5.52e-10
+ ub1 = -2.16e-18
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.3 pmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 1.495e-06 wmax = 1.505e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.94224+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_3+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.58139
+ k2 = {0.019018+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_3}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {150350+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_3}
+ ua = {2.6796985e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_3}
+ ub = {1.7457e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_3}
+ uc = -1.4632e-12
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_3}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.020291+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_3}
+ a0 = {0.85794+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_3}
+ keta = {-0.0096207+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_3}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.13498+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_3}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_3}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_3}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.099014101+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_3+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.0709+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_3+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_3}
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_3}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.84169+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_3}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00129
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 2.1831475e+8
+ pscbe2 = 1.4985163e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.0150852e-5
+ alpha1 = 0.0
+ beta0 = 37.469254
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_3}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_3}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.22e-008+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_3}
+ bgidl = {1.5831e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_3}
+ cgidl = {576+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_3}
+ egidl = 0.89190707
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.6000+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_3}
+ kt2 = -0.019032
+ at = 10000.0
+ ute = -1.3908
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.4 pmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 1.495e-06 wmax = 1.505e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.94224+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_4+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.58139
+ k2 = {0.019018391+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_4}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {180350+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_4}
+ ua = {2.6796985e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_4}
+ ub = {1.7457e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_4}
+ uc = -3.6579e-11
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_4}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.020291+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_4}
+ a0 = {0.85794+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_4}
+ keta = {-0.0096207+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_4}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.14983+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_4}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_4}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_4}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.099014101+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_4+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.0709+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_4+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_4}
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_4}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.84169224+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_4}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00129
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 2.1831475e+8
+ pscbe2 = 1.4985163e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.0150852e-5
+ alpha1 = 0.0
+ beta0 = 37.469254
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_4}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_4}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {2e-008+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_4}
+ bgidl = {1.6008e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_4}
+ cgidl = {1200+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_4}
+ egidl = 0.89190707
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.59+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_4}
+ kt2 = -0.019032
+ at = 291500.0
+ ute = -1.4098
+ ua1 = 5.524e-10
+ ub1 = -4.2529e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.5 pmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 1.495e-06 wmax = 1.505e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.95024+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_5+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.58139
+ k2 = {0.019018391+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_5}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {180350+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_5}
+ ua = {2.6796985e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_5}
+ ub = {3.1073e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_5}
+ uc = -2.3647e-11
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_5}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.0211+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_5}
+ a0 = {0.9609+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_5}
+ keta = {-0.0096207+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_5}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.13498356+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_5}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_5}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_5}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.099014101+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_5+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.0709+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_5+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_5}
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_5}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.84169224+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_5}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00129
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 2.1831475e+8
+ pscbe2 = 1.4985163e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.0150852e-5
+ alpha1 = 0.0
+ beta0 = 37.469254
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_5}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_5}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {9.8e-009+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_5}
+ bgidl = {1.7927e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_5}
+ cgidl = {468+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_5}
+ egidl = 0.89190707
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.596+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_5}
+ kt2 = -0.019032
+ at = 341570.0
+ ute = -1.5561
+ ua1 = 2.2096e-11
+ ub1 = -3.7536e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.6 pmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 1.495e-06 wmax = 1.505e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.94153+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_6+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.5906
+ k2 = {0.030282+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_6}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {83300+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_6}
+ ua = {1.7880272e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_6}
+ ub = {1.2353e-018+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_6}
+ uc = -3.6698e-12
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_6}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.017957+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_6}
+ a0 = {0.81545+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_6}
+ keta = {-0.048114+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_6}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.84632+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_6}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_6}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_6}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.091667534+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_6+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.5024+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_6+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_6}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.059291+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_6}
+ etab = -0.013965
+ dsub = 0.27363
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {1.035+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_6}
+ pdiblc1 = 0.18699149
+ pdiblc2 = 0.0038831667
+ pdiblcb = -0.025
+ drout = 1.0
+ pscbe1 = 3.4108348e+8
+ pscbe2 = 1.4750539e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.8189581e-5
+ alpha1 = 0.0
+ beta0 = 45.963568
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_6}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_6}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {8.4723e-009+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_6}
+ bgidl = {1.6871e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_6}
+ cgidl = {500+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_6}
+ egidl = 0.64214944
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.63348+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_6}
+ kt2 = -0.019032
+ at = 5000.0
+ ute = -1.2996
+ ua1 = 5.52e-10
+ ub1 = -2.16e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.7 pmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.906+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_7+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.59627
+ k2 = {0.015964796+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_7}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {45904+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_7}
+ ua = {9.3613665e-010+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_7}
+ ub = {1.4921e-018+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_7}
+ uc = -2.2219153e-12
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_7}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.015822+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_7}
+ a0 = {0.87287+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_7}
+ keta = {-0.087434+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_7}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.70436855+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_7}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_7}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_7}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.079644655+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_7+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.2953+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_7+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_7}
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.039542+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_7}
+ etab = -0.00078616
+ dsub = 0.30791359
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {1.267944+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_7}
+ pdiblc1 = 0.32524895
+ pdiblc2 = 0.0020127014
+ pdiblcb = -0.025
+ drout = 0.99999967
+ pscbe1 = 3.1103691e+8
+ pscbe2 = 1.4418397e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.4232853e-5
+ alpha1 = 0.0
+ beta0 = 49.951734
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_7}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_7}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.8816e-009+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_7}
+ bgidl = {1.543e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_7}
+ cgidl = {360.18+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_7}
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.6380+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_7}
+ kt2 = -0.019032
+ at = 30000.0
+ ute = -1.4498
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.8 pmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.92805+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_8+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.59348
+ k2 = {0.017615423+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_8}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {21066+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_8}
+ ua = {1.6523781e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_8}
+ ub = {9.7216e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_8}
+ uc = -1.2317537e-11
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_8}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.018029+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_8}
+ a0 = {0.96928+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_8}
+ keta = {-0.11488+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_8}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.73757129+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_8}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_8}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_8}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.086157622+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_8+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.2919+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_8+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_8}
+ cit = 6.9459796e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_8}
+ etab = -0.000648
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {1.9035348+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_8}
+ pdiblc1 = 0.3909083
+ pdiblc2 = 0.00129
+ pdiblcb = -0.025
+ drout = 0.63800017
+ pscbe1 = 3.0990248e+8
+ pscbe2 = 1.4767911e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00031976739
+ alpha1 = 0.0
+ beta0 = 55.34354
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_8}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_8}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {4e-008+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_8}
+ bgidl = {1.6056e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_8}
+ cgidl = {840+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_8}
+ egidl = 1.4570704
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.615+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_8}
+ kt2 = -0.019032
+ at = 16836.0
+ ute = -1.4038
+ ua1 = 7.7336e-10
+ ub1 = -2.8009e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.9 pmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.926+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_9+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.6051
+ k2 = {0.015276967+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_9}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {120230+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_9}
+ ua = {1.9671141e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_9}
+ ub = {5.3455e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_9}
+ uc = -2.9902062e-11
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_9}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.018494+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_9}
+ a0 = {0.86595+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_9}
+ keta = {-0.0098272+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_9}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.13659769+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_9}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_9}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_9}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.097070481+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_9+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {0.99229+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_9+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_9}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_9}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.91362237+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_9}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00129
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 2.2505867e+8
+ pscbe2 = 1.5007389e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_9}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_9}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {3.36e-008+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_9}
+ bgidl = {1.4723e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_9}
+ cgidl = {492+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_9}
+ egidl = 2.0
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.576+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_9}
+ kt2 = -0.019032
+ at = 219650.0
+ ute = -1.4104
+ ua1 = 2.2096e-11
+ ub1 = -2.3998e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.10 pmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.94868+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_10+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.58485
+ k2 = {0.020475051+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_10}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {80156+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_10}
+ ua = {2.2507416e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_10}
+ ub = {3.4083e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_10}
+ uc = -4.5108582e-11
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_10}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.01919+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_10}
+ a0 = {0.90565+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_10}
+ keta = {-0.0081819+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_10}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.13283238+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_10}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_10}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_10}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.10768013+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_10+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {0.94783+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_10+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_10}
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_10}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.08353125+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_10}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0034380666
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 2.2471761e+8
+ pscbe2 = 1.4998723e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 6.4242641e-5
+ alpha1 = 0.0
+ beta0 = 39.039478
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_10}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_10}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {2e-008+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_10}
+ bgidl = {1.5204e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_10}
+ cgidl = {1400+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_10}
+ egidl = 1.5199352
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.556+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_10}
+ kt2 = -0.019032
+ at = 151090.0
+ ute = -1.5561
+ ua1 = 2.2096e-11
+ ub1 = -3.0767e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.11 pmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope2/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.89504+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_11+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.55947
+ k2 = {0.036713432+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_11}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {117570+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_11}
+ ua = {1.2669543e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_11}
+ ub = {1.2082e-018+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_11}
+ uc = -5.9494373e-12
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_11}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.016056+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_11}
+ a0 = {0.72074+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_11}
+ keta = {-0.0084885+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_11}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.11578365+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_11}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_11}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_11}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11318245+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_11+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.2536+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_11+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_11}
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.15643+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_11}
+ etab = -0.010946
+ dsub = 0.27819971
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.64077291+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_11}
+ pdiblc1 = 0.13281489
+ pdiblc2 = 0.0020780138
+ pdiblcb = -0.225
+ drout = 1.0
+ pscbe1 = 8.0e+8
+ pscbe2 = 5.6866809e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.0002497e-6
+ alpha1 = 0.0
+ beta0 = 38.089036
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_11}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_11}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.24e-008+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_11}
+ bgidl = {2.0463e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_11}
+ cgidl = {300+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_11}
+ egidl = 0.1352153
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.60348+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_11}
+ kt2 = -0.019032
+ at = 1000.0
+ ute = -1.2208
+ ua1 = 5.52e-10
+ ub1 = -2.16e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.12 pmos
* DC IV MOS Parameters
+ lmin = 5.95e-07 lmax = 6.05e-07 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.91036+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_12+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.62735
+ k2 = {0.017816539+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_12}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {74424+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_12}
+ ua = {1.2023341e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_12}
+ ub = {1.4559e-018+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_12}
+ uc = -2.7539501e-12
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_12}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.016763+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_12}
+ a0 = {0.84201+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_12}
+ keta = {-0.051484+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_12}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.72220108+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_12}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_12}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_12}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.079967669+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_12+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.473+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_12+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_12}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.017878+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_12}
+ etab = 0.0
+ dsub = 0.27181946
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {1.0998724+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_12}
+ pdiblc1 = 0.39855546
+ pdiblc2 = 0.0078480034
+ pdiblcb = -0.025
+ drout = 0.64228671
+ pscbe1 = 3.3852051e+8
+ pscbe2 = 1.4615273e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.9655204e-5
+ alpha1 = 0.0
+ beta0 = 48.175076
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_12}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_12}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {4.7e-008+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_12}
+ bgidl = {1.5488e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_12}
+ cgidl = {966+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_12}
+ egidl = 1.2131988
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.65348+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_12}
+ kt2 = -0.019032
+ at = 10000.0
+ ute = -1.3412
+ ua1 = 5.52e-10
+ ub1 = -1.8696e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.13 pmos
* DC IV MOS Parameters
+ lmin = 7.95e-07 lmax = 8.05e-07 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.88436+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_13+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.57696
+ k2 = {0.02202554+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_13}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {57942+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_13}
+ ua = {1.3736548e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_13}
+ ub = {1.2992e-018+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_13}
+ uc = -1.8899043e-12
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_13}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.016917+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_13}
+ a0 = {0.79601+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_13}
+ keta = {-0.064617+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_13}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.7357361+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_13}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_13}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_13}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.083615082+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_13+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.4934+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_13+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_13}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.0068242+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_13}
+ etab = -0.0040945
+ dsub = 0.26520582
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {1.152681+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_13}
+ pdiblc1 = 0.45413396
+ pdiblc2 = 0.0066035801
+ pdiblcb = -0.025
+ drout = 0.54609838
+ pscbe1 = 3.6891994e+8
+ pscbe2 = 1.3484359e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.2455677e-5
+ alpha1 = 0.0
+ beta0 = 47.447604
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_13}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_13}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {7.7552e-009+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_13}
+ bgidl = {1.7886e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_13}
+ cgidl = {510+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_13}
+ egidl = 0.16211671
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.6405+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_13}
+ kt2 = -0.019032
+ at = 20000.0
+ ute = -1.4798
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.14 pmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 1.9995e-05 wmax = 2.0005e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.97224+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_14+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.57939
+ k2 = {0.020277+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_14}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {47889+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_14}
+ ua = {1.6494295e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_14}
+ ub = {1.0975e-018+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_14}
+ uc = -5.8546e-13
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_14}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.020384+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_14}
+ a0 = {0.85515+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_14}
+ keta = {-0.084672+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_14}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.77943+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_14}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_14}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_14}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.077755783+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_14+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.3116+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_14+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_14}
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {2.8641e-005+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_14}
+ etab = 0.0
+ dsub = 0.54416
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {1.2031+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_14}
+ pdiblc1 = 0.3995264
+ pdiblc2 = 0.0015061847
+ pdiblcb = -0.025
+ drout = 0.41068941
+ pscbe1 = 2.994803e+8
+ pscbe2 = 1.4554569e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 6.7813161e-5
+ alpha1 = 0.0
+ beta0 = 50.152925
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_14}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_14}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.085e-008+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_14}
+ bgidl = {1.6213e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_14}
+ cgidl = {500.48+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_14}
+ egidl = 0.77897916
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.6362+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_14}
+ kt2 = -0.019032
+ at = 29800.0
+ ute = -1.6069
+ ua1 = 4.1982e-10
+ ub1 = -3.8064e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.15 pmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 1.9995e-05 wmax = 2.0005e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.9885+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_15+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.59804
+ k2 = {0.024041+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_15}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {67000+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_15}
+ ua = {2.1590772e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_15}
+ ub = {9.5539e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_15}
+ uc = -5.2815e-12
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_15}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.022232+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_15}
+ a0 = {0.95964+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_15}
+ keta = {-0.08587+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_15}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {1.25+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_15}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_15}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_15}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.10153677+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_15+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.1999+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_15+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_15}
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.080055+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_15}
+ etab = -0.0038503
+ dsub = 0.27967
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {1.3366+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_15}
+ pdiblc1 = 0.29403034
+ pdiblc2 = 0.0048008826
+ pdiblcb = -0.025
+ drout = 0.89960455
+ pscbe1 = 3.6263996e+8
+ pscbe2 = 1.448673e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 9.713535e-5
+ alpha1 = 0.0
+ beta0 = 54.684511
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_15}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_15}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.3888e-008+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_15}
+ bgidl = {1.6145e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_15}
+ cgidl = {876+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_15}
+ egidl = 0.66526877
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.61348+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_15}
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.3724
+ ua1 = 5.52e-10
+ ub1 = -2.16e-18
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.16 pmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.94424+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_16+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.57939
+ k2 = {0.020277382+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_16}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {47889+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_16}
+ ua = {1.6494295e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_16}
+ ub = {1.2762e-018+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_16}
+ uc = -5.8546e-13
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_16}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.019197+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_16}
+ a0 = {0.85515+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_16}
+ keta = {-0.084672+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_16}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.72169009+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_16}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_16}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_16}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.077755783+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_16+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.3116+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_16+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_16}
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.0087749+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_16}
+ etab = 0.0
+ dsub = 0.2989895
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {1.2031125+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_16}
+ pdiblc1 = 0.3995264
+ pdiblc2 = 0.0015061847
+ pdiblcb = -0.025
+ drout = 0.41068941
+ pscbe1 = 2.994803e+8
+ pscbe2 = 1.4554569e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 6.7813161e-5
+ alpha1 = 0.0
+ beta0 = 50.152925
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_16}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_16}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {6.0144e-009+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_16}
+ bgidl = {1.5638e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_16}
+ cgidl = {920+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_16}
+ egidl = 0.77897916
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.6300+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_16}
+ kt2 = -0.019032
+ at = 30000.0
+ ute = -1.4608
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.17 pmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.97089+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_17+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56874
+ k2 = {0.021845+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_17}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {136210+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_17}
+ ua = {2.5957213e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_17}
+ ub = {5.9095e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_17}
+ uc = 0.0
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_17}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.021802+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_17}
+ a0 = {0.92576+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_17}
+ keta = {-0.01712+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_17}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.19+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_17}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_17}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_17}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.12041324+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_17+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.2+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_17+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_17}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.1438+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_17}
+ etab = -0.015108
+ dsub = 0.29315
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.60569+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_17}
+ pdiblc1 = 0.1893326
+ pdiblc2 = 0.003828528
+ pdiblcb = -0.225
+ drout = 1.0
+ pscbe1 = 3.6834658e+8
+ pscbe2 = 1.4543145e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_17}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_17}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {9.3141e-009+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_17}
+ bgidl = {1.2201e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_17}
+ cgidl = {468.55+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_17}
+ egidl = 2.0
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.575+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_17}
+ kt2 = -0.019032
+ at = 171730.0
+ ute = -1.4498
+ ua1 = 5.524e-10
+ ub1 = -4.1218e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.18 pmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.97767+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_18+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.58606
+ k2 = {0.019966+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_18}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {124910+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_18}
+ ua = {2.9651633e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_18}
+ ub = {1.3357e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_18}
+ uc = -2.8099e-11
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_18}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.022592+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_18}
+ a0 = {0.8749+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_18}
+ keta = {-0.010964+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_18}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.15682+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_18}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_18}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_18}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.091596347+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_18+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {0.8+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_18+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_18}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_18}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.83237107+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_18}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00129
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 1.0e+8
+ pscbe2 = 4.602312e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.2543089e-5
+ alpha1 = 0.0
+ beta0 = 37.371509
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_18}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_18}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {9.4e-009+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_18}
+ bgidl = {1.8618e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_18}
+ cgidl = {660+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_18}
+ egidl = 0.16572358
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.576+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_18}
+ kt2 = -0.019032
+ at = 229660.0
+ ute = -1.5561
+ ua1 = 2.2096e-11
+ ub1 = -3.7536e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.19 pmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.97709+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_19+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.59521
+ k2 = {0.019927+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_19}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {200000+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_19}
+ ua = {2.7044348e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_19}
+ ub = {1.4379e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_19}
+ uc = -3.9972e-11
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_19}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.021226+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_19}
+ a0 = {0.89552+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_19}
+ keta = {-0.0079259+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_19}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.1318+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_19}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_19}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_19}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_19+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.0849+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_19+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_19}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_19}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.08353125+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_19}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 3.3371283e+8
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_19}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_19}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.4775e-008+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_19}
+ bgidl = {1.7757e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_19}
+ cgidl = {1000+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_19}
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.576+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_19}
+ kt2 = -0.019032
+ at = 448800.0
+ ute = -1.5361
+ ua1 = 2.2096e-11
+ ub1 = -3.6627e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.20 pmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.95089+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_20+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56874
+ k2 = {0.028835+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_20}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {130760+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_20}
+ ua = {2.5957213e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_20}
+ ub = {4.0614e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_20}
+ uc = -3.6e-11
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_20}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.020518+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_20}
+ a0 = {0.92576+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_20}
+ keta = {-0.00090104+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_20}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.19+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_20}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_20}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_20}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.12041324+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_20+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.2+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_20+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_20}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.1438+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_20}
+ etab = -0.015108
+ dsub = 0.29315
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.60569+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_20}
+ pdiblc1 = 0.1893326
+ pdiblc2 = 0.003828528
+ pdiblcb = -0.225
+ drout = 1.0
+ pscbe1 = 3.6834658e+8
+ pscbe2 = 1.4543145e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_20}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_20}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.63e-008+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_20}
+ bgidl = {1.2201e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_20}
+ cgidl = {768.42+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_20}
+ egidl = 2.0
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.58948+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_20}
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.2724
+ ua1 = 5.52e-10
+ ub1 = -2.894e-18
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.21 pmos
* DC IV MOS Parameters
+ lmin = 5.95e-07 lmax = 6.05e-07 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.93332+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_21+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.57633
+ k2 = {0.025668+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_21}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {78336+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_21}
+ ua = {2.3466113e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_21}
+ ub = {4.9371e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_21}
+ uc = -2.4658e-12
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_21}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.019791+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_21}
+ a0 = {0.84351+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_21}
+ keta = {-0.043025+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_21}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.72112+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_21}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_21}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_21}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.072821331+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_21+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.495+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_21+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_21}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.00024193+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_21}
+ etab = 0.0
+ dsub = 0.27482
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.97221+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_21}
+ pdiblc1 = 0.45695731
+ pdiblc2 = 0.011410926
+ pdiblcb = -0.025
+ drout = 0.43179535
+ pscbe1 = 4.0e+8
+ pscbe2 = 1.3503615e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.7240171e-5
+ alpha1 = 0.0
+ beta0 = 45.34673
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_21}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_21}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.1694e-008+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_21}
+ bgidl = {1.8073e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_21}
+ cgidl = {520+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_21}
+ egidl = 0.48103697
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.64548+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_21}
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.4573
+ ua1 = 5.52e-10
+ ub1 = -3.2992e-18
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.22 pmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.94824+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_22+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.57939
+ k2 = {0.020277+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_22}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {47889+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_22}
+ ua = {1.6494295e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_22}
+ ub = {1.0975e-018+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_22}
+ uc = -5.8546e-13
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_22}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.019197+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_22}
+ a0 = {0.85515+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_22}
+ keta = {-0.084672+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_22}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.77943+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_22}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_22}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_22}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.077755783+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_22+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.3116+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_22+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_22}
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.00052649+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_22}
+ etab = 0.0
+ dsub = 0.29899
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {1.2031125+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_22}
+ pdiblc1 = 0.3995264
+ pdiblc2 = 0.0015061847
+ pdiblcb = -0.025
+ drout = 0.41068941
+ pscbe1 = 2.994803e+8
+ pscbe2 = 1.4554569e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 6.7813161e-5
+ alpha1 = 0.0
+ beta0 = 50.152925
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_22}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_22}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {9.2738e-009+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_22}
+ bgidl = {1.5638e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_22}
+ cgidl = {368+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_22}
+ egidl = 0.77897916
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.6300+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_22}
+ kt2 = -0.019032
+ at = 30000.0
+ ute = -1.4608
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.23 pmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.98389+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_23+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56874
+ k2 = {0.021845+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_23}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {126210+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_23}
+ ua = {2.5957213e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_23}
+ ub = {8.9538e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_23}
+ uc = 0.0
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_23}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.023194+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_23}
+ a0 = {0.92576+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_23}
+ keta = {-0.01712+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_23}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.19+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_23}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_23}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_23}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.12041324+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_23+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.2+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_23+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_23}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.1438+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_23}
+ etab = -0.015108
+ dsub = 0.29315
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.60569082+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_23}
+ pdiblc1 = 0.1893326
+ pdiblc2 = 0.003828528
+ pdiblcb = -0.225
+ drout = 1.0
+ pscbe1 = 3.6834658e+8
+ pscbe2 = 1.4543145e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_23}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_23}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {9.7022e-009+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_23}
+ bgidl = {1.2201e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_23}
+ cgidl = {468.55+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_23}
+ egidl = 2.0
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.5750+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_23}
+ kt2 = -0.019032
+ at = 104800.0
+ ute = -1.4498
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.24 pmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.98767+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_24+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.58606
+ k2 = {0.019966+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_24}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {124910+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_24}
+ ua = {2.9651633e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_24}
+ ub = {2.244e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_24}
+ uc = -2.8099e-11
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_24}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.023496+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_24}
+ a0 = {0.8749+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_24}
+ keta = {-0.010964+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_24}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.15682+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_24}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_24}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_24}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.091596347+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_24+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {0.8+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_24+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_24}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_24}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.83237107+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_24}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00129
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 1.0e+8
+ pscbe2 = 4.602312e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.2543089e-5
+ alpha1 = 0.0
+ beta0 = 37.371509
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_24}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_24}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {7.896e-009+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_24}
+ bgidl = {1.8618e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_24}
+ cgidl = {660+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_24}
+ egidl = 0.16572358
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.576+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_24}
+ kt2 = -0.019032
+ at = 235700.0
+ ute = -1.5561
+ ua1 = 2.2096e-11
+ ub1 = -3.8766e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.25 pmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.99209+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_25+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.59521
+ k2 = {0.019927+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_25}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {200000+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_25}
+ ua = {2.7044348e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_25}
+ ub = {3.9379e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_25}
+ uc = -3.9972e-11
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_25}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.0225+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_25}
+ a0 = {0.89552+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_25}
+ keta = {-0.0079259+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_25}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.1318+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_25}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_25}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_25}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_25+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.0849+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_25+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_25}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_25}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.08353125+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_25}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 3.3371283e+8
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_25}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_25}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.5366e-008+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_25}
+ bgidl = {1.7047e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_25}
+ cgidl = {1000+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_25}
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.576+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_25}
+ kt2 = -0.019032
+ at = 448800.0
+ ute = -1.5361
+ ua1 = 2.2096e-11
+ ub1 = -3.6627e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.26 pmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.98229+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_26+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.58637
+ k2 = {0.02619+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_26}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {73540+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_26}
+ ua = {2.8298029e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_26}
+ ub = {5.993e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_26}
+ uc = -9.8477e-12
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_26}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.02333+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_26}
+ a0 = {0.79883+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_26}
+ keta = {-0.075644+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_26}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {1.25+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_26}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_26}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_26}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.13295587+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_26+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.3232+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_26+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_26}
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.040327+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_26}
+ etab = -0.010229
+ dsub = 0.29048905
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {1.184192+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_26}
+ pdiblc1 = 0.39269218
+ pdiblc2 = 0.0079692374
+ pdiblcb = -0.025
+ drout = 0.72266506
+ pscbe1 = 3.1758291e+8
+ pscbe2 = 1.4459233e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.4081425e-5
+ alpha1 = 0.0
+ beta0 = 50.534039
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_26}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_26}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.1634e-008+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_26}
+ bgidl = {1.6718e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_26}
+ cgidl = {400+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_26}
+ egidl = 0.67432849
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.58348+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_26}
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.3724
+ ua1 = 5.52e-10
+ ub1 = -2.894e-18
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.27 pmos
* DC IV MOS Parameters
+ lmin = 5.95e-07 lmax = 6.05e-07 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.96559+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_27+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56924
+ k2 = {0.025929+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_27}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {60844+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_27}
+ ua = {4.0655985e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_27}
+ ub = {-5.6854e-021+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_27}
+ uc = -4.527e-12
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_27}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.027729+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_27}
+ a0 = {0.80598+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_27}
+ keta = {-0.096905+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_27}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {1.25+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_27}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_27}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_27}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.10586774+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_27+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.3874+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_27+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_27}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.023711+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_27}
+ etab = 0.0
+ dsub = 0.30839886
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {1.2669585+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_27}
+ pdiblc1 = 0.56716046
+ pdiblc2 = 0.0054000816
+ pdiblcb = -0.025
+ drout = 0.89134169
+ pscbe1 = 3.8734436e+8
+ pscbe2 = 1.4665318e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.1782526e-5
+ alpha1 = 0.0
+ beta0 = 52.761864
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_27}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_27}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {6.5211e-009+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_27}
+ bgidl = {1.7072e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_27}
+ cgidl = {230+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_27}
+ egidl = 0.76686217
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.61848+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_27}
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.4273
+ ua1 = 5.52e-10
+ ub1 = -3.2992e-18
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.28 pmos
* DC IV MOS Parameters
+ lmin = 7.95e-07 lmax = 8.05e-07 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.93332+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_28+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.57633
+ k2 = {0.025668+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_28}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {61200+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_28}
+ ua = {2.3466113e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_28}
+ ub = {7.4804e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_28}
+ uc = -2.4658e-12
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_28}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.021512+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_28}
+ a0 = {0.84351+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_28}
+ keta = {-0.06519+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_28}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.72112+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_28}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_28}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_28}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.072821331+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_28+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.495+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_28+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_28}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.00071157+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_28}
+ etab = -0.00053192
+ dsub = 0.27482351
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.97220765+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_28}
+ pdiblc1 = 0.45695731
+ pdiblc2 = 0.011410926
+ pdiblcb = -0.025
+ drout = 0.43179535
+ pscbe1 = 4.0e+8
+ pscbe2 = 1.3503615e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.7240171e-5
+ alpha1 = 0.0
+ beta0 = 45.34673
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_28}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_28}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.6706e-008+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_28}
+ bgidl = {1.8073e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_28}
+ cgidl = {520+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_28}
+ egidl = 0.48103697
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.6405+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_28}
+ kt2 = -0.019032
+ at = 25000.0
+ ute = -1.4798
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.29 pmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.96224+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_29+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.57939
+ k2 = {0.020277+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_29}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {47889+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_29}
+ ua = {1.6494295e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_29}
+ ub = {1.0975e-018+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_29}
+ uc = -5.8546e-13
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_29}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.0196+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_29}
+ a0 = {0.85515+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_29}
+ keta = {-0.084672+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_29}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.77943+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_29}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_29}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_29}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.077755783+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_29+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.3116+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_29+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_29}
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {4.2119e-005+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_29}
+ etab = 0.0
+ dsub = 0.54416
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {1.2031125+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_29}
+ pdiblc1 = 0.3995264
+ pdiblc2 = 0.0015061847
+ pdiblcb = -0.025
+ drout = 0.41068941
+ pscbe1 = 2.994803e+8
+ pscbe2 = 1.4554569e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 6.7813161e-5
+ alpha1 = 0.0
+ beta0 = 50.152925
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_29}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_29}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {8.3464e-009+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_29}
+ bgidl = {1.6889e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_29}
+ cgidl = {368+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_29}
+ egidl = 0.77897916
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.6300+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_29}
+ kt2 = -0.019032
+ at = 30000.0
+ ute = -1.4608
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.30 pmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.98989+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_30+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.56874
+ k2 = {0.021845+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_30}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {116210+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_30}
+ ua = {2.5957213e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_30}
+ ub = {8.9538e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_30}
+ uc = 0.0
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_30}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.023594+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_30}
+ a0 = {0.92576+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_30}
+ keta = {-0.01712+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_30}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.19+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_30}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_30}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_30}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.12041324+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_30+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.2+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_30+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_30}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.1438+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_30}
+ etab = -0.015108
+ dsub = 0.29315
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.60569082+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_30}
+ pdiblc1 = 0.1893326
+ pdiblc2 = 0.003828528
+ pdiblcb = -0.225
+ drout = 1.0
+ pscbe1 = 3.6834658e+8
+ pscbe2 = 1.4543145e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_30}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_30}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {7.1796e-009+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_30}
+ bgidl = {1.2201e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_30}
+ cgidl = {468.55+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_30}
+ egidl = 2.0
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.5650+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_30}
+ kt2 = -0.019032
+ at = 150800.0
+ ute = -1.4000
+ ua1 = 5.524e-10
+ ub1 = -3.6627e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.31 pmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.99467+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_31+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.58606
+ k2 = {0.019966+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_31}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {100010+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_31}
+ ua = {2.9651633e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_31}
+ ub = {2.244e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_31}
+ uc = -2.8099e-11
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_31}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.024036+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_31}
+ a0 = {0.8749+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_31}
+ keta = {-0.010964+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_31}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.15682+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_31}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_31}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_31}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.091596347+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_31+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {0.8+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_31+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_31}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_31}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.83237107+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_31}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00129
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 1.0e+8
+ pscbe2 = 4.602312e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.2543089e-5
+ alpha1 = 0.0
+ beta0 = 37.371509
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_31}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_31}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {8.2118e-009+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_31}
+ bgidl = {1.9363e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_31}
+ cgidl = {462+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_31}
+ egidl = 0.16572358
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.566+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_31}
+ kt2 = -0.019032
+ at = 181310.0
+ ute = -1.5561
+ ua1 = 2.2096e-11
+ ub1 = -3.6920e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.32 pmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-1+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_32+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.59521
+ k2 = {0.019927+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_32}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {200000+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_32}
+ ua = {2.7044348e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_32}
+ ub = {3.9379e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_32}
+ uc = -3.9972e-11
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_32}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.0229+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_32}
+ a0 = {0.89552+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_32}
+ keta = {-0.0079259+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_32}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.1318+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_32}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_32}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_32}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.093204657+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_32+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.0849+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_32+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_32}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_32}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.08353125+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_32}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029407877
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 3.3371283e+8
+ pscbe2 = 1.5000958e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0667189e-5
+ alpha1 = 0.0
+ beta0 = 38.266046
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_32}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_32}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {7.3657e-009+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_32}
+ bgidl = {1.7047e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_32}
+ cgidl = {700+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_32}
+ egidl = 0.69350825
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.57573+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_32}
+ kt2 = -0.019032
+ at = 430000.0
+ ute = -1.3864
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.33 pmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.9675+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_33+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.59804
+ k2 = {0.024041+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_33}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {67000+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_33}
+ ua = {2.1590772e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_33}
+ ub = {9.5539e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_33}
+ uc = -5.2815e-12
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_33}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.021377+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_33}
+ a0 = {0.95964+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_33}
+ keta = {-0.08587+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_33}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {1.25+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_33}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_33}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_33}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.10153677+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_33+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.1999+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_33+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_33}
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.080055+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_33}
+ etab = -0.0038503
+ dsub = 0.27967
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {1.3366321+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_33}
+ pdiblc1 = 0.29403034
+ pdiblc2 = 0.0048008826
+ pdiblcb = -0.025
+ drout = 0.89960455
+ pscbe1 = 3.6263996e+8
+ pscbe2 = 1.448673e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 9.713535e-5
+ alpha1 = 0.0
+ beta0 = 54.684511
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_33}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_33}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.02e-008+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_33}
+ bgidl = {1.5572e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_33}
+ cgidl = {174+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_33}
+ egidl = 0.66526877
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.60348+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_33}
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.3724
+ ua1 = 5.52e-10
+ ub1 = -2.16e-18
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.34 pmos
* DC IV MOS Parameters
+ lmin = 7.95e-07 lmax = 8.05e-07 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.949+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_34+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.57633
+ k2 = {0.025668+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_34}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {61200+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_34}
+ ua = {2.3466113e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_34}
+ ub = {7.4804e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_34}
+ uc = -2.4658e-12
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_34}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.022+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_34}
+ a0 = {0.84351+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_34}
+ keta = {-0.06519+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_34}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.72112+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_34}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_34}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_34}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.072821331+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_34+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.495+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_34+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_34}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {5.6926e-005+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_34}
+ etab = -0.00021277
+ dsub = 0.27482
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.97220765+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_34}
+ pdiblc1 = 0.45695731
+ pdiblc2 = 0.011410926
+ pdiblcb = -0.025
+ drout = 0.43179535
+ pscbe1 = 4.0e+8
+ pscbe2 = 1.3503615e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.7240171e-5
+ alpha1 = 0.0
+ beta0 = 45.34673
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_34}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_34}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.136e-008+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_34}
+ bgidl = {1.8073e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_34}
+ cgidl = {520+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_34}
+ egidl = 0.48103697
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.6435+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_34}
+ kt2 = -0.019032
+ at = 25000.0
+ ute = -1.4798
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.35 pmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.90360217+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_35+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.58237463
+ k2 = {0.021666466+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_35}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {89566+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_35}
+ ua = {1.7625428e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_35}
+ ub = {5.4082628e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_35}
+ uc = -4.2959383e-12
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_35}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.018653409+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_35}
+ a0 = {0.63337751+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_35}
+ keta = {-0.012595257+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_35}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.128125+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_35}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_35}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_35}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.088381148+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_35+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.4655+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_35+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_35}
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.28744+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_35}
+ etab = -0.00077252
+ dsub = 0.26831464
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.97281896+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_35}
+ pdiblc1 = 0.42058379
+ pdiblc2 = 0.0011725831
+ pdiblcb = -0.025
+ drout = 0.87592071
+ pscbe1 = 3.089798e+8
+ pscbe2 = 1.4883743e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.053402e-5
+ alpha1 = 0.0
+ beta0 = 40.210566
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_35}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_35}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5e-008+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_35}
+ bgidl = {1.7848738e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_35}
+ cgidl = {1000+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_35}
+ egidl = 0.76372321
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.6400+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_35}
+ kt2 = -0.019032
+ at = 10000.0
+ ute = -1.4498
+ ua1 = 5.524e-10
+ ub1 = -2.8959e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.36 pmos
* DC IV MOS Parameters
+ lmin = 1.9995e-05 lmax = 2.0005e-05 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.95807+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_36+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.60281
+ k2 = {0.018238228+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_36}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {26719+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_36}
+ ua = {1.5847414e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_36}
+ ub = {7.8391e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_36}
+ uc = -4.1711723e-11
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_36}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.018506+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_36}
+ a0 = {0.90435+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_36}
+ keta = {-0.0042037+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_36}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.10781371+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_36}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_36}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_36}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.12217944+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_36+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {0.8+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_36+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_36}
+ cit = 9.1876579e-8
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_36}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.08353125+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_36}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00129
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 2.25e+8
+ pscbe2 = 1.5e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_36}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_36}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1e-008+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_36}
+ bgidl = {1.2463e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_36}
+ cgidl = {1400+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_36}
+ egidl = 2.0
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.55573+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_36}
+ kt2 = -0.019032
+ at = 46800.0
+ ute = -1.4448
+ ua1 = 7.0656e-10
+ ub1 = -3.145e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.37 pmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.95955+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_37+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.59139
+ k2 = {0.019352451+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_37}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {130850+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_37}
+ ua = {1.9590891e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_37}
+ ub = {5.3943007e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_37}
+ uc = -1.1497139e-11
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_37}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.020158+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_37}
+ a0 = {0.88+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_37}
+ keta = {-0.009+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_37}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.10+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_37}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_37}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_37}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.10401589+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_37+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.0056+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_37+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_37}
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.49+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_37}
+ etab = -1.0565
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {1.8727984+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_37}
+ pdiblc1 = 0.58340637
+ pdiblc2 = 0.00129
+ pdiblcb = -0.025
+ drout = 0.31028214
+ pscbe1 = 2.9284027e+8
+ pscbe2 = 1.4741685e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.7693836e-6
+ alpha1 = 0.0
+ beta0 = 35.270704
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_37}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_37}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {6.86e-008+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_37}
+ bgidl = {1.5689515e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_37}
+ cgidl = {1152+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_37}
+ egidl = 1.4760927
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.588+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_37}
+ kt2 = -0.019032
+ at = 184000.0
+ ute = -1.35
+ ua1 = 5.524e-10
+ ub1 = -3.2036e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.38 pmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.96107+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_38+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.59047
+ k2 = {0.018746757+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_38}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {120230+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_38}
+ ua = {2.1146882e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_38}
+ ub = {2.5096855e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_38}
+ uc = -2.7456539e-11
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_38}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.020131+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_38}
+ a0 = {0.81+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_38}
+ keta = {-0.0050598+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_38}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.11483891+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_38}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_38}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_38}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.10968052+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_38+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.005+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_38+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_38}
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_38}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {1.2961212+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_38}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00129
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 2.2500144e+8
+ pscbe2 = 1.5000011e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.206037e-5
+ alpha1 = 0.0
+ beta0 = 36.963614
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_38}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_38}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {6.37e-008+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_38}
+ bgidl = {1.5860386e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_38}
+ cgidl = {1200+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_38}
+ egidl = 1.3291649
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.566+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_38}
+ kt2 = -0.019032
+ at = 219650.0
+ ute = -1.4424
+ ua1 = 2.2096e-11
+ ub1 = -2.3998e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.39 pmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.9723+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_39+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.55533
+ k2 = {0.030745+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_39}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {80156+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_39}
+ ua = {2.2137527e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_39}
+ ub = {2.7518e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_39}
+ uc = -3.1546e-11
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_39}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.020541+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_39}
+ a0 = {0.88+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_39}
+ keta = {-0.0051528+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_39}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.11911+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_39}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_39}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_39}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.12715703+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_39+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.134+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_39+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_39}
+ cit = 2.5e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_39}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.083531+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_39}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0056422857
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 2.25e+8
+ pscbe2 = 1.5e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_39}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_39}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {7e-008+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_39}
+ bgidl = {1.3e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_39}
+ cgidl = {1485+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_39}
+ egidl = 2.0
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.546+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_39}
+ kt2 = -0.019032
+ at = 151090.0
+ ute = -1.5561
+ ua1 = 2.2096e-11
+ ub1 = -3.0767e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.40 pmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.93514+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_40+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.5044
+ k2 = {0.047795+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_40}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {96000+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_40}
+ ua = {2.520839e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_40}
+ ub = {-3.95e-021+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_40}
+ uc = -7.0465e-12
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_40}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.020095+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_40}
+ a0 = {0.023438+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_40}
+ keta = {-0.0087101+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_40}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.024023+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_40}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_40}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_40}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.08150653+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_40+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.8602+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_40+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_40}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.0042715+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_40}
+ etab = -0.021343
+ dsub = 0.27992
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {1.0922+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_40}
+ pdiblc1 = 0.38852895
+ pdiblc2 = 0.0069782586
+ pdiblcb = -0.025
+ drout = 0.82656681
+ pscbe1 = 3.6230113e+8
+ pscbe2 = 1.4700248e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0979853e-5
+ alpha1 = 0.0
+ beta0 = 43.428559
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_40}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_40}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {4.144e-008+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_40}
+ bgidl = {1.671e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_40}
+ cgidl = {767.95+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_40}
+ egidl = 1.1526517
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.64948+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_40}
+ kt2 = -0.019032
+ at = 18000.0
+ ute = -1.3624
+ ua1 = 5.52e-10
+ ub1 = -2.894e-18
+ uc1 = -4.1496e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.41 pmos
* DC IV MOS Parameters
+ lmin = 5.95e-07 lmax = 6.05e-07 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.90453619+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_41+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.53447619
+ k2 = {0.039396842+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_41}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {85096.792+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_41}
+ ua = {1.173516e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_41}
+ ub = {1.222731e-018+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_41}
+ uc = -4.6607993e-12
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_41}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.016303299+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_41}
+ a0 = {0.63343726+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_41}
+ keta = {-0.019041557+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_41}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.43242187+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_41}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_41}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_41}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11136124+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_41+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.3719842+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_41+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_41}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.094454882+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_41}
+ etab = -0.035896073
+ dsub = 0.29420499
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {1.0997509+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_41}
+ pdiblc1 = 0.35412617
+ pdiblc2 = 0.0032399298
+ pdiblcb = -0.025
+ drout = 0.71796338
+ pscbe1 = 3.8500909e+8
+ pscbe2 = 1.3804759e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.9848596e-5
+ alpha1 = 0.0
+ beta0 = 45.089194
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_41}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_41}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {8e-008+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_41}
+ bgidl = {1.5810321e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_41}
+ cgidl = {1908.2+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_41}
+ egidl = 1.3390402
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.60348+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_41}
+ kt2 = -0.019032
+ at = 10000.0
+ ute = -1.2412
+ ua1 = 5.52e-10
+ ub1 = -1.8696e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.42 pmos
* DC IV MOS Parameters
+ lmin = 7.95e-07 lmax = 8.05e-07 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.9264+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_42+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.52566309
+ k2 = {0.035643+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_42}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {77067+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_42}
+ ua = {1.5643566e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_42}
+ ub = {6.5919e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_42}
+ uc = -4.3553868e-12
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_42}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.018908+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_42}
+ a0 = {0.76528248+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_42}
+ keta = {-0.029626108+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_42}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.40595436+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_42}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_42}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_42}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11007505+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_42+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.3820472+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_42+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_42}
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.49+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_42}
+ etab = -6.25e-6
+ dsub = 0.46919791
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.99477438+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_42}
+ pdiblc1 = 0.40166422
+ pdiblc2 = 0.0064917125
+ pdiblcb = -0.025
+ drout = 0.51082388
+ pscbe1 = 3.0891221e+8
+ pscbe2 = 1.4440738e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_42}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_42}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {6.824e-007+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_42}
+ bgidl = {1.5947033e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_42}
+ cgidl = {5748.2+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_42}
+ egidl = 2.0
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.6175+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_42}
+ kt2 = -0.019032
+ at = 10000.0
+ ute = -1.4798
+ ua1 = 5.524e-10
+ ub1 = -2.8959e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.43 pmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 7.45e-07 wmax = 7.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.88639+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_43+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.55984
+ k2 = {0.026386144+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_43}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {69528+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_43}
+ ua = {2.0341039e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_43}
+ ub = {5.878e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_43}
+ uc = -2.7970035e-12
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_43}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.018442+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_43}
+ a0 = {0.73934+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_43}
+ keta = {-0.032622+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_43}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.43242187+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_43}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_43}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_43}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.075734118+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_43+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.5401+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_43+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_43}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.036111+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_43}
+ etab = -0.0043407
+ dsub = 0.31595571
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {1.1707598+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_43}
+ pdiblc1 = 0.54661982
+ pdiblc2 = 0.0020306546
+ pdiblcb = -0.025
+ drout = 0.42584153
+ pscbe1 = 2.7813655e+8
+ pscbe2 = 1.4513967e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_43}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_43}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.056e-010+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_43}
+ bgidl = {1.0285e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_43}
+ cgidl = {994.06+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_43}
+ egidl = 0.90967406
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.6480+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_43}
+ kt2 = -0.019032
+ at = 30000.0
+ ute = -1.4498
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.44 pmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 7.45e-07 wmax = 7.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.904+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_44+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.55984
+ k2 = {0.026386144+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_44}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {38200+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_44}
+ ua = {2.0341039e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_44}
+ ub = {6.4658e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_44}
+ uc = -2.7970035e-12
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_44}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.01918+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_44}
+ a0 = {0.73934+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_44}
+ keta = {-0.037189+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_44}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.43242187+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_44}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_44}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_44}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.075734118+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_44+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.5401+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_44+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_44}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.06+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_44}
+ etab = 0.0
+ dsub = 0.31595571
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {1.1707598+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_44}
+ pdiblc1 = 0.54661982
+ pdiblc2 = 0.0020306546
+ pdiblcb = -0.025
+ drout = 0.42584153
+ pscbe1 = 2.7813655e+8
+ pscbe2 = 1.4513967e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_44}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_44}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {1.056e-010+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_44}
+ bgidl = {1.0285e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_44}
+ cgidl = {1670+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_44}
+ egidl = 0.90967406
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.6480+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_44}
+ kt2 = -0.019032
+ at = 34800.0
+ ute = -1.4498
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.45 pmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 7.45e-07 wmax = 7.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.93527+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_45+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.57102
+ k2 = {0.023085+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_45}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {180350+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_45}
+ ua = {2.334849e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_45}
+ ub = {3.4026e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_45}
+ uc = -3.2639e-11
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_45}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.020132+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_45}
+ a0 = {0.87668+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_45}
+ keta = {-0.0076977+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_45}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.1244+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_45}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_45}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_45}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.10903374+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_45+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.0655+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_45+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_45}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.08+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_45}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.99495+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_45}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00129
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 2.2560035e+8
+ pscbe2 = 1.4994384e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.8978653e-5
+ alpha1 = 0.0
+ beta0 = 37.686511
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_45}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_45}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {3.08e-008+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_45}
+ bgidl = {1.7019e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_45}
+ cgidl = {1200+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_45}
+ egidl = 1.0890786
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.566+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_45}
+ kt2 = -0.019032
+ at = 351440.0
+ ute = -1.4104
+ ua1 = 2.2096e-11
+ ub1 = -2.3998e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.46 pmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 7.45e-07 wmax = 7.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.92036+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_46+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.53224
+ k2 = {0.046095+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_46}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {80727+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_46}
+ ua = {1.8760013e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_46}
+ ub = {1.0003e-018+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_46}
+ uc = -5.0888e-12
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_46}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.017891+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_46}
+ a0 = {0.68242+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_46}
+ keta = {-0.04781+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_46}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.98885+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_46}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_46}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_46}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.099269478+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_46+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.7634+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_46+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_46}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.068197+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_46}
+ etab = -0.0043723
+ dsub = 0.26967
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {1.0392+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_46}
+ pdiblc1 = 0.18044532
+ pdiblc2 = 0.0037051928
+ pdiblcb = -0.025
+ drout = 1.0
+ pscbe1 = 4.0e+8
+ pscbe2 = 1.4741409e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.9436447e-5
+ alpha1 = 0.0
+ beta0 = 46.62143
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_46}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_46}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {3.32e-008+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_46}
+ bgidl = {1.7842e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_46}
+ cgidl = {840+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_46}
+ egidl = 0.92927294
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.64848+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_46}
+ kt2 = -0.019032
+ at = 5000.0
+ ute = -1.3696
+ ua1 = 5.52e-10
+ ub1 = -2.6784e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.47 pmos
* DC IV MOS Parameters
+ lmin = 7.95e-07 lmax = 8.05e-07 wmin = 7.45e-07 wmax = 7.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.88639+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_47+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.55984
+ k2 = {0.026386144+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_47}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {75574+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_47}
+ ua = {2.0341039e-009+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_47}
+ ub = {5.878e-019+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_47}
+ uc = -2.7970035e-12
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_47}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.019002+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_47}
+ a0 = {0.73934+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_47}
+ keta = {-0.032622+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_47}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.43242187+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_47}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_47}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_47}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.075734118+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_47+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.5401+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_47+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_47}
+ cit = 1.0e-5
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.036111+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_47}
+ etab = -0.0043407
+ dsub = 0.31595571
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {1.1707598+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_47}
+ pdiblc1 = 0.54661982
+ pdiblc2 = 0.0020306546
+ pdiblcb = -0.025
+ drout = 0.42584153
+ pscbe1 = 2.7813655e+8
+ pscbe2 = 1.4513967e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_47}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_47}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {2.4e-010+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_47}
+ bgidl = {1.0285e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_47}
+ cgidl = {994.06+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_47}
+ egidl = 0.90967406
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.6475+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_47}
+ kt2 = -0.019032
+ at = 10000.0
+ ute = -1.4798
+ ua1 = 5.524e-10
+ ub1 = -3.5909e-18
+ uc1 = -1.092e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_g5v0d10v5__model.48 pmos
* DC IV MOS Parameters
+ lmin = 5.95e-07 lmax = 6.05e-07 wmin = 6.95e-07 wmax = 7.05e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.175e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {4.5375e-008+sky130_fd_pr__pfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {1.2277e-008+sky130_fd_pr__pfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.7338e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.37
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.175e-008*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(1.175e-08*sky130_fd_pr__pfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__pfet_g5v0d10v5__toxe_slope3/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__pfet_g5v0d10v5__rshp_mult}
* Threshold Voltage Parameters
+ vth0 = {-0.87115+sky130_fd_pr__pfet_g5v0d10v5__vth0_diff_48+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.57069
+ k2 = {0.030351152+sky130_fd_pr__pfet_g5v0d10v5__k2_diff_48}
+ k3 = -2.2405
+ dvt0 = 4.657
+ dvt1 = 0.34864
+ dvt2 = -0.030206
+ dvt0w = -2.2
+ dvt1w = 1016300.0
+ dvt2w = 0.0
+ w0 = 0.0
+ k3b = -0.172
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {68461+sky130_fd_pr__pfet_g5v0d10v5__vsat_diff_48}
+ ua = {9.5685789e-010+sky130_fd_pr__pfet_g5v0d10v5__ua_diff_48}
+ ub = {1.6857e-018+sky130_fd_pr__pfet_g5v0d10v5__ub_diff_48}
+ uc = -2.8451032e-12
+ rdsw = {788.47+sky130_fd_pr__pfet_g5v0d10v5__rdsw_diff_48}
+ prwb = 0.053538
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.015405+sky130_fd_pr__pfet_g5v0d10v5__u0_diff_48}
+ a0 = {0.81031+sky130_fd_pr__pfet_g5v0d10v5__a0_diff_48}
+ keta = {-0.073162+sky130_fd_pr__pfet_g5v0d10v5__keta_diff_48}
+ a1 = 0.0
+ a2 = 0.5
+ ags = {0.9538163+sky130_fd_pr__pfet_g5v0d10v5__ags_diff_48}
+ b0 = {0+sky130_fd_pr__pfet_g5v0d10v5__b0_diff_48}
+ b1 = {0+sky130_fd_pr__pfet_g5v0d10v5__b1_diff_48}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.10729755+sky130_fd_pr__pfet_g5v0d10v5__voff_diff_48+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.2484+sky130_fd_pr__pfet_g5v0d10v5__nfactor_diff_48+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_g5v0d10v5__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__pfet_g5v0d10v5__tvoff_diff_48}
+ cit = 5.0e-6
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.020883+sky130_fd_pr__pfet_g5v0d10v5__eta0_diff_48}
+ etab = 0.0
+ dsub = 0.29051085
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {1.2193396+sky130_fd_pr__pfet_g5v0d10v5__pclm_diff_48}
+ pdiblc1 = 0.59952915
+ pdiblc2 = 0.0045454479
+ pdiblcb = -0.025
+ drout = 0.99912731
+ pscbe1 = 4.0e+8
+ pscbe2 = 1.4479847e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.4267536e-5
+ alpha1 = 0.0
+ beta0 = 49.499633
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {0+sky130_fd_pr__pfet_g5v0d10v5__pdits_diff_48}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__pfet_g5v0d10v5__pditsd_diff_48}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {2.91e-008+sky130_fd_pr__pfet_g5v0d10v5__agidl_diff_48}
+ bgidl = {1.7407e009+sky130_fd_pr__pfet_g5v0d10v5__bgidl_diff_48}
+ cgidl = {800+sky130_fd_pr__pfet_g5v0d10v5__cgidl_diff_48}
+ egidl = 0.95326514
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.175e-8
* Temperature Effects Parameters
+ kt1 = {-0.60348+sky130_fd_pr__pfet_g5v0d10v5__kt1_diff_48}
+ kt2 = -0.019032
+ at = 10000.0
+ ute = -1.3412
+ ua1 = 5.52e-10
+ ub1 = -1.8696e-18
+ uc1 = -3.7128e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0000000e+40
+ noib = 8.5300000e+24
+ noic = 8.4000000e+7
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 4.02e-12
+ xtis = 10.0
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.00096
+ tcjsw = 3.0e-5
+ tcjswg = 0.0
+ cgdo = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgso = {1.9771e-010*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cgdl = {1.0005e-011*sky130_fd_pr__pfet_g5v0d10v5__overlap_mult}
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {4.4983e-008+sky130_fd_pr__pfet_g5v0d10v5__dlc_diff+sky130_fd_pr__pfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__pfet_g5v0d10v5__dwc_diff}
+ vfbcv = -0.1446893
+ acde = 0.401
+ moin = 15.773
+ noff = 4.0
+ voffcv = 0.0
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.00077547*sky130_fd_pr__pfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.33956
+ pbs = 0.6587
+ cjsws = {9.8717e-011*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.24676
+ pbsws = 1.0
+ cjswgs = {1.46e-010*sky130_fd_pr__pfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.81
+ pbswgs = 3.0
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+sky130_fd_pr__pfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.ends sky130_fd_pr__pfet_g5v0d10v5
