**.subckt Bandgap1.8v_2_meas_post
x1 Vdd Vref 0 Bandgap 
**** begin user architecture code

.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/cells/nfet_01v8/sky130_fd_pr__nfet_01v8__tt.corner.spice
.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/cells/nfet_01v8_lvt/sky130_fd_pr__nfet_01v8_lvt__tt.corner.spice
.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/cells/pfet_01v8/sky130_fd_pr__pfet_01v8__tt.corner.spice
.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/cells/nfet_03v3_nvt/sky130_fd_pr__nfet_03v3_nvt__tt.corner.spice
.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/cells/nfet_05v0_nvt/sky130_fd_pr__nfet_05v0_nvt__tt.corner.spice
.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/cells/esd_nfet_01v8/sky130_fd_pr__esd_nfet_01v8__tt.corner.spice
.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/cells/pfet_01v8_lvt/sky130_fd_pr__pfet_01v8_lvt__tt.corner.spice
.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/cells/pfet_01v8_hvt/sky130_fd_pr__pfet_01v8_hvt__tt.corner.spice
.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/cells/esd_pfet_g5v0d10v5/sky130_fd_pr__esd_pfet_g5v0d10v5__tt.corner.spice
.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/cells/pfet_g5v0d10v5/sky130_fd_pr__pfet_g5v0d10v5__tt.corner.spice
.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/cells/pfet_g5v0d16v0/sky130_fd_pr__pfet_g5v0d16v0__tt.corner.spice
.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/cells/nfet_g5v0d10v5/sky130_fd_pr__nfet_g5v0d10v5__tt.corner.spice
.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/cells/nfet_g5v0d16v0/sky130_fd_pr__nfet_g5v0d16v0__tt_discrete.corner.spice
.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/cells/esd_nfet_g5v0d10v5/sky130_fd_pr__esd_nfet_g5v0d10v5__tt.corner.spice
.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/models/corners/tt/nonfet.spice
* Mismatch parameters
.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/cells/nfet_01v8/sky130_fd_pr__nfet_01v8__mismatch.corner.spice
.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/cells/pfet_01v8/sky130_fd_pr__pfet_01v8__mismatch.corner.spice
.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/cells/nfet_01v8_lvt/sky130_fd_pr__nfet_01v8_lvt__mismatch.corner.spice
.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/cells/pfet_01v8_lvt/sky130_fd_pr__pfet_01v8_lvt__mismatch.corner.spice
.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/cells/pfet_01v8_hvt/sky130_fd_pr__pfet_01v8_hvt__mismatch.corner.spice
.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/cells/nfet_g5v0d10v5/sky130_fd_pr__nfet_g5v0d10v5__mismatch.corner.spice
.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/cells/pfet_g5v0d10v5/sky130_fd_pr__pfet_g5v0d10v5__mismatch.corner.spice
.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/cells/nfet_05v0_nvt/sky130_fd_pr__nfet_05v0_nvt__mismatch.corner.spice
.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/cells/nfet_03v3_nvt/sky130_fd_pr__nfet_03v3_nvt__mismatch.corner.spice
* Resistor
.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/models/r+c/res_typical__cap_typical.spice
.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/models/r+c/res_typical__cap_typical__lin.spice
* Special cells
.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/models/corners/tt/specialized_cells.spice
* All models
.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/models/all.spice
* Corner
.include ~/Analog_blocks/models/skywater-pdk/libraries/sky130_fd_pr/latest/models/corners/tt/rf.spice



************************************************
*Source initialization
************************************************
Vsup Vdd 0 DC 0 AC 0
************************************************
*Temp variation
************************************************
.control
alter Vsup DC = 1.8
dc temp -40 120 1
show
plot vref
meas DC Vref_27 FIND Vref AT=27
meas DC Vref_neg40 FIND Vref AT=-40
meas DC Vref_120 FIND Vref AT=120
.endc
************************************************
*Supply variation
************************************************
.control
dc Vsup 0 3 0.5
plot vdd vref
meas DC Vref_nom FIND Vref AT=1.8
meas DC Vref_Sup_pos10per FIND Vref AT=1.62
meas DC Vref_Sup_neg10per FIND Vref AT=1.98
.endc
************************************************
*PSRR analysis
************************************************
.control
alter Vsup DC = 1.8
alter Vsup AC = 1
ac dec 10 1 100MEG
plot db(vref)
meas ac PSR_1k FIND vdb(Vref) AT=1k
meas ac PSR_1M FIND vdb(vref) AT=1Meg
.endc
************************************************
*Transient analysis
************************************************
.control
alter @Vsup[pwl] = [ 0 0 100u 0 200u 3 500u 3 ]
tran 100u 500u
plot vdd vref
.endc
************************************************

**** end user architecture code
**.ends

* expanding   symbol:
.subckt Bandgap VDD Vref GND
*.ipin VDD
*.ipin GND
*.opin Vref
XM0 G1011.t87 G1011.t86 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM1 G1011.t92 D6.t10 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
XM2 GND D6.t11 G1011.t89 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
XM3 D5.t3 G1011.t98 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XQ4 GND GND VBJTS GND sky130_fd_pr__pnp_05v5_W0p68L0p68 
XM5 VDD G1011.t84 G1011.t85 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM6 VDD G1011.t82 G1011.t83 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM7 D9.t5 G4 D5.t5 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=500000u
XM8 G1011.t90 D6.t12 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
XM9 GND D6.t13 G1011.t97 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
XR1694 G3.t0 Vref.t4 GND sky130_fd_pr__res_xhigh_po_1p41 w=1.41e+06u l=1.8e+06u
XM11 VDD G1011.t99 D5.t2 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM12 VDD G1011.t100 Vref.t3 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
XM13 VDD G1011.t80 G1011.t81 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XQ14 GND GND G4 GND sky130_fd_pr__pnp_05v5_W0p68L0p68 
XM15 GND D9.t12 D9.t13 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
XM16 D5.t15 G3.t1 D6.t5 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=500000u
XM17 G1011.t79 G1011.t78 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM18 VDD G1011.t76 G1011.t77 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM19 VDD G1011.t74 G1011.t75 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM20 VDD G1011.t72 G1011.t73 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM21 VDD G1011.t70 G1011.t71 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XQ22 GND GND VBJTS GND sky130_fd_pr__pnp_05v5_W0p68L0p68 
XM23 VDD G1011.t68 G1011.t69 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM24 G1011.t67 G1011.t66 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM25 G1011.t65 G1011.t64 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XQ26 GND GND VBJTS GND sky130_fd_pr__pnp_05v5_W0p68L0p68 
XM27 G1011.t96 D6.t14 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
XM28 G1011.t63 G1011.t62 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM29 D6.t3 G3.t2 D5.t13 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=500000u
XM30 G1011.t61 G1011.t60 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM31 G1011.t59 G1011.t58 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM32 G1011.t94 D6.t15 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
XM33 D6.t6 D9.t14 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
XR1695 a_523_n9665# a_n7_n8873# GND sky130_fd_pr__res_xhigh_po_1p41 w=1.41e+06u l=1.8e+06u
XM35 G1011.t57 G1011.t56 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XR1696 a_2643_n9665# a_3173_n8873# GND sky130_fd_pr__res_xhigh_po_1p41 w=1.41e+06u l=1.8e+06u
XM37 VDD G1011.t54 G1011.t55 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM38 D5.t11 G3.t3 D6.t1 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=500000u
XM39 VDD G1011.t52 G1011.t53 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM40 D1011.t2 G1011.t101 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=1e+06u
XM41 VDD G1011.t50 G1011.t51 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM42 GND D9.t10 D9.t11 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
XM43 GND D6.t16 G1011.t93 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
XM44 Vref.t2 G1011.t102 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
XM45 G4 D1011.t3 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=1e+06u
XM46 G1011.t49 G1011.t48 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XQ47 GND GND VBJTS GND sky130_fd_pr__pnp_05v5_W0p68L0p68 
XM48 G1011.t47 G1011.t46 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM49 VDD G1011.t44 G1011.t45 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM50 D9.t9 D9.t8 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
XM51 VDD G1011.t103 D2.t3 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
XR1697 G3.t0 a_n7_n8873# GND sky130_fd_pr__res_xhigh_po_1p41 w=1.41e+06u l=1.8e+06u
XM53 D2.t2 G1011.t104 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
XR1698 G4 a_3173_n8873# GND sky130_fd_pr__res_xhigh_po_1p41 w=1.41e+06u l=1.8e+06u
XM55 D5.t14 G3.t4 D6.t4 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=500000u
XM56 GND D9.t15 D6.t7 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
XM57 G1011.t43 G1011.t42 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM58 VDD D1011.t4 G4 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=1e+06u
XM59 G1011.t41 G1011.t40 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM60 D6.t8 D9.t16 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
XM61 VDD G1011.t105 D1011.t1 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=1e+06u
XM62 VDD G1011.t106 Vref.t1 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
XM63 G1011.t39 G1011.t38 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM64 D6.t2 G3.t5 D5.t12 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=500000u
XM65 D5.t4 G4 D9.t4 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=500000u
XM66 D1011.t0 G1011.t107 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=2e+07u
XQ67 GND GND VBJTS GND sky130_fd_pr__pnp_05v5_W0p68L0p68 
XR1699 a_2643_n9665# a_2113_n8873# GND sky130_fd_pr__res_xhigh_po_1p41 w=1.41e+06u l=1.8e+06u
XM69 G1011.t37 G1011.t36 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM70 G1011.t35 G1011.t34 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM71 GND D9.t17 D6.t9 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
XM72 D5.t9 G4 D9.t3 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=500000u
XM73 D2.t1 G1011.t108 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
XM74 D6.t0 G3.t6 D5.t10 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=500000u
XM75 VDD G1011.t32 G1011.t33 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM76 VDD G1011.t30 G1011.t31 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM77 G1011.t29 G1011.t28 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XQ78 GND GND VBJTS GND sky130_fd_pr__pnp_05v5_W0p68L0p68 
XM79 VDD G1011.t109 D2.t0 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
XM80 G1011.t27 G1011.t26 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM81 G1011.t25 G1011.t24 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM82 G1011.t23 G1011.t22 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XQ83 GND GND VBJTS GND sky130_fd_pr__pnp_05v5_W0p68L0p68 
XM84 VDD G1011.t20 G1011.t21 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM85 Vref.t0 G1011.t110 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
XR1700 VBJTS a_1053_n8873# GND sky130_fd_pr__res_xhigh_po_1p41 w=1.41e+06u l=1.8e+06u
XR1701 D2.t4 a_2113_n8873# GND sky130_fd_pr__res_xhigh_po_1p41 w=1.41e+06u l=1.8e+06u
XM88 VDD G1011.t18 G1011.t19 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM89 VDD G1011.t16 G1011.t17 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM90 VDD G1011.t14 G1011.t15 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM91 D9.t7 D9.t6 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
XM92 D9.t2 G4 D5.t8 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=500000u
XM93 G1011.t13 G1011.t12 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM94 G1011.t11 G1011.t10 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM95 VDD G1011.t111 D5.t1 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM96 D9.t1 G4 D5.t7 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=500000u
XQ97 GND GND VBJTS GND sky130_fd_pr__pnp_05v5_W0p68L0p68 
XM98 D5.t0 G1011.t112 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM99 GND D6.t17 G1011.t91 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
XM100 VDD G1011.t8 G1011.t9 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM101 VDD G1011.t6 G1011.t7 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM102 G1011.t95 D6.t18 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
XR1702 a_523_n9665# a_1053_n8873# GND sky130_fd_pr__res_xhigh_po w=1.41e+06u l=1.8e+06u
XM104 D5.t6 G4 D9.t0 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=500000u
XM105 VDD G1011.t4 G1011.t5 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM106 GND D6.t19 G1011.t88 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u
XM107 G1011.t3 G1011.t2 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XM108 VDD G1011.t0 G1011.t1 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
XR0 G1011.n98 G1011.t101 517.956
XR1 G1011.n183 G1011.t105 482
XR2 G1011.t105 G1011.n182 482
XR3 G1011.n206 G1011.t108 361.93
XR4 G1011.n200 G1011.t109 361.93
XR5 G1011.n206 G1011.t103 361.501
XR6 G1011.n207 G1011.t102 361.501
XR7 G1011.n208 G1011.t100 361.501
XR8 G1011.n201 G1011.t106 361.501
XR9 G1011.n200 G1011.t104 361.501
XR10 G1011.n51 G1011.t110 293.262
XR11 G1011.n224 G1011.t68 168.915
XR12 G1011.n236 G1011.t86 168.915
XR13 G1011.n235 G1011.t30 168.701
XR14 G1011.n277 G1011.t34 168.701
XR15 G1011.n276 G1011.t70 168.701
XR16 G1011.n293 G1011.t56 168.701
XR17 G1011.n292 G1011.t32 168.701
XR18 G1011.n309 G1011.t36 168.701
XR19 G1011.n308 G1011.t72 168.701
XR20 G1011.n325 G1011.t10 168.701
XR21 G1011.n324 G1011.t18 168.701
XR22 G1011.n341 G1011.t64 168.701
XR23 G1011.n340 G1011.t74 168.701
XR24 G1011.n357 G1011.t12 168.701
XR25 G1011.n356 G1011.t44 168.701
XR26 G1011.n373 G1011.t48 168.701
XR27 G1011.n372 G1011.t20 168.701
XR28 G1011.n389 G1011.t28 168.701
XR29 G1011.n388 G1011.t52 168.701
XR30 G1011.n405 G1011.t58 168.701
XR31 G1011.n404 G1011.t6 168.701
XR32 G1011.n423 G1011.t66 168.701
XR33 G1011.n422 G1011.t76 168.701
XR34 G1011.n421 G1011.t98 168.701
XR35 G1011.n420 G1011.t111 168.701
XR36 G1011.n439 G1011.t112 168.701
XR37 G1011.n440 G1011.t99 168.701
XR38 G1011.n441 G1011.t38 168.701
XR39 G1011.n438 G1011.t4 168.701
XR40 G1011.n457 G1011.t2 168.701
XR41 G1011.n456 G1011.t80 168.701
XR42 G1011.n473 G1011.t42 168.701
XR43 G1011.n472 G1011.t8 168.701
XR44 G1011.n489 G1011.t62 168.701
XR45 G1011.n488 G1011.t54 168.701
XR46 G1011.n505 G1011.t26 168.701
XR47 G1011.n504 G1011.t0 168.701
XR48 G1011.n521 G1011.t60 168.701
XR49 G1011.n520 G1011.t50 168.701
XR50 G1011.n537 G1011.t24 168.701
XR51 G1011.n536 G1011.t84 168.701
XR52 G1011.n553 G1011.t46 168.701
XR53 G1011.n552 G1011.t16 168.701
XR54 G1011.n217 G1011.t22 168.701
XR55 G1011.n219 G1011.t82 168.701
XR56 G1011.n220 G1011.t40 168.701
XR57 G1011.n222 G1011.t14 168.701
XR58 G1011.n223 G1011.t78 168.701
XR59 G1011.n53 G1011.n285 152
XR60 G1011.n280 G1011.n279 152
XR61 G1011.n53 G1011.n284 152
XR62 G1011.n288 G1011.n287 152
XR63 G1011.n52 G1011.n282 152
XR64 G1011.n52 G1011.n281 152
XR65 G1011.n55 G1011.n301 152
XR66 G1011.n296 G1011.n295 152
XR67 G1011.n55 G1011.n300 152
XR68 G1011.n304 G1011.n303 152
XR69 G1011.n54 G1011.n298 152
XR70 G1011.n54 G1011.n297 152
XR71 G1011.n57 G1011.n317 152
XR72 G1011.n312 G1011.n311 152
XR73 G1011.n57 G1011.n316 152
XR74 G1011.n320 G1011.n319 152
XR75 G1011.n56 G1011.n314 152
XR76 G1011.n56 G1011.n313 152
XR77 G1011.n59 G1011.n333 152
XR78 G1011.n328 G1011.n327 152
XR79 G1011.n59 G1011.n332 152
XR80 G1011.n336 G1011.n335 152
XR81 G1011.n58 G1011.n330 152
XR82 G1011.n58 G1011.n329 152
XR83 G1011.n61 G1011.n349 152
XR84 G1011.n344 G1011.n343 152
XR85 G1011.n61 G1011.n348 152
XR86 G1011.n352 G1011.n351 152
XR87 G1011.n60 G1011.n346 152
XR88 G1011.n60 G1011.n345 152
XR89 G1011.n63 G1011.n365 152
XR90 G1011.n360 G1011.n359 152
XR91 G1011.n63 G1011.n364 152
XR92 G1011.n368 G1011.n367 152
XR93 G1011.n62 G1011.n362 152
XR94 G1011.n62 G1011.n361 152
XR95 G1011.n65 G1011.n381 152
XR96 G1011.n376 G1011.n375 152
XR97 G1011.n65 G1011.n380 152
XR98 G1011.n384 G1011.n383 152
XR99 G1011.n64 G1011.n378 152
XR100 G1011.n64 G1011.n377 152
XR101 G1011.n67 G1011.n397 152
XR102 G1011.n392 G1011.n391 152
XR103 G1011.n67 G1011.n396 152
XR104 G1011.n400 G1011.n399 152
XR105 G1011.n66 G1011.n394 152
XR106 G1011.n66 G1011.n393 152
XR107 G1011.n69 G1011.n413 152
XR108 G1011.n408 G1011.n407 152
XR109 G1011.n69 G1011.n412 152
XR110 G1011.n416 G1011.n415 152
XR111 G1011.n68 G1011.n410 152
XR112 G1011.n68 G1011.n409 152
XR113 G1011.n71 G1011.n431 152
XR114 G1011.n426 G1011.n425 152
XR115 G1011.n71 G1011.n430 152
XR116 G1011.n434 G1011.n433 152
XR117 G1011.n70 G1011.n428 152
XR118 G1011.n70 G1011.n427 152
XR119 G1011.n73 G1011.n449 152
XR120 G1011.n444 G1011.n443 152
XR121 G1011.n73 G1011.n448 152
XR122 G1011.n452 G1011.n451 152
XR123 G1011.n72 G1011.n446 152
XR124 G1011.n72 G1011.n445 152
XR125 G1011.n75 G1011.n465 152
XR126 G1011.n460 G1011.n459 152
XR127 G1011.n75 G1011.n464 152
XR128 G1011.n468 G1011.n467 152
XR129 G1011.n74 G1011.n462 152
XR130 G1011.n74 G1011.n461 152
XR131 G1011.n77 G1011.n481 152
XR132 G1011.n476 G1011.n475 152
XR133 G1011.n77 G1011.n480 152
XR134 G1011.n484 G1011.n483 152
XR135 G1011.n76 G1011.n478 152
XR136 G1011.n76 G1011.n477 152
XR137 G1011.n79 G1011.n497 152
XR138 G1011.n492 G1011.n491 152
XR139 G1011.n79 G1011.n496 152
XR140 G1011.n500 G1011.n499 152
XR141 G1011.n78 G1011.n494 152
XR142 G1011.n78 G1011.n493 152
XR143 G1011.n81 G1011.n513 152
XR144 G1011.n508 G1011.n507 152
XR145 G1011.n81 G1011.n512 152
XR146 G1011.n516 G1011.n515 152
XR147 G1011.n80 G1011.n510 152
XR148 G1011.n80 G1011.n509 152
XR149 G1011.n83 G1011.n529 152
XR150 G1011.n524 G1011.n523 152
XR151 G1011.n83 G1011.n528 152
XR152 G1011.n532 G1011.n531 152
XR153 G1011.n82 G1011.n526 152
XR154 G1011.n82 G1011.n525 152
XR155 G1011.n85 G1011.n545 152
XR156 G1011.n540 G1011.n539 152
XR157 G1011.n85 G1011.n544 152
XR158 G1011.n548 G1011.n547 152
XR159 G1011.n84 G1011.n542 152
XR160 G1011.n84 G1011.n541 152
XR161 G1011.n87 G1011.n561 152
XR162 G1011.n556 G1011.n555 152
XR163 G1011.n87 G1011.n560 152
XR164 G1011.n564 G1011.n563 152
XR165 G1011.n86 G1011.n558 152
XR166 G1011.n86 G1011.n557 152
XR167 G1011.n89 G1011.n574 152
XR168 G1011.n569 G1011.n568 152
XR169 G1011.n89 G1011.n573 152
XR170 G1011.n577 G1011.n576 152
XR171 G1011.n88 G1011.n571 152
XR172 G1011.n88 G1011.n570 152
XR173 G1011.n91 G1011.n582 152
XR174 G1011.n216 G1011.n215 152
XR175 G1011.n91 G1011.n581 152
XR176 G1011.n584 G1011.n583 152
XR177 G1011.n90 G1011.n212 152
XR178 G1011.n90 G1011.n213 152
XR179 G1011.n92 G1011.n227 152
XR180 G1011.n93 G1011.n230 152
XR181 G1011.n92 G1011.n228 152
XR182 G1011.n226 G1011.n225 152
XR183 G1011.n234 G1011.n233 152
XR184 G1011.n93 G1011.n231 152
XR185 G1011.n95 G1011.n243 152
XR186 G1011.n95 G1011.n242 152
XR187 G1011.n94 G1011.n240 152
XR188 G1011.n94 G1011.n239 152
XR189 G1011.n238 G1011.n237 152
XR190 G1011.n246 G1011.n245 152
XR191 G1011.n3 G1011.t90 131.509
XR192 G1011.n270 G1011.t91 131.056
XR193 G1011.n251 G1011.n250 91.699
XR194 G1011.n256 G1011.n255 91.699
XR195 G1011.n261 G1011.n260 91.699
XR196 G1011.n266 G1011.n265 91.699
XR197 G1011.n250 G1011.t88 39.357
XR198 G1011.n250 G1011.t94 39.357
XR199 G1011.n255 G1011.t89 39.357
XR200 G1011.n255 G1011.t95 39.357
XR201 G1011.n260 G1011.t93 39.357
XR202 G1011.n260 G1011.t96 39.357
XR203 G1011.n265 G1011.t97 39.357
XR204 G1011.n265 G1011.t92 39.357
XR205 G1011.n113 G1011.n112 29.029
XR206 G1011.n121 G1011.n120 29.029
XR207 G1011.n232 G1011.t69 27.695
XR208 G1011.n232 G1011.t79 27.695
XR209 G1011.n286 G1011.t71 27.695
XR210 G1011.n286 G1011.t35 27.695
XR211 G1011.n302 G1011.t33 27.695
XR212 G1011.n302 G1011.t57 27.695
XR213 G1011.n318 G1011.t73 27.695
XR214 G1011.n318 G1011.t37 27.695
XR215 G1011.n334 G1011.t19 27.695
XR216 G1011.n334 G1011.t11 27.695
XR217 G1011.n350 G1011.t75 27.695
XR218 G1011.n350 G1011.t65 27.695
XR219 G1011.n366 G1011.t45 27.695
XR220 G1011.n366 G1011.t13 27.695
XR221 G1011.n382 G1011.t21 27.695
XR222 G1011.n382 G1011.t49 27.695
XR223 G1011.n398 G1011.t53 27.695
XR224 G1011.n398 G1011.t29 27.695
XR225 G1011.n414 G1011.t7 27.695
XR226 G1011.n414 G1011.t59 27.695
XR227 G1011.n432 G1011.t77 27.695
XR228 G1011.n432 G1011.t67 27.695
XR229 G1011.n450 G1011.t5 27.695
XR230 G1011.n450 G1011.t39 27.695
XR231 G1011.n466 G1011.t81 27.695
XR232 G1011.n466 G1011.t3 27.695
XR233 G1011.n482 G1011.t9 27.695
XR234 G1011.n482 G1011.t43 27.695
XR235 G1011.n498 G1011.t55 27.695
XR236 G1011.n498 G1011.t63 27.695
XR237 G1011.n514 G1011.t1 27.695
XR238 G1011.n514 G1011.t27 27.695
XR239 G1011.n530 G1011.t51 27.695
XR240 G1011.n530 G1011.t61 27.695
XR241 G1011.n546 G1011.t85 27.695
XR242 G1011.n546 G1011.t25 27.695
XR243 G1011.n562 G1011.t17 27.695
XR244 G1011.n562 G1011.t47 27.695
XR245 G1011.n575 G1011.t83 27.695
XR246 G1011.n575 G1011.t23 27.695
XR247 G1011.n214 G1011.t15 27.695
XR248 G1011.n214 G1011.t41 27.695
XR249 G1011.n244 G1011.t31 27.695
XR250 G1011.n244 G1011.t87 27.695
XR251 G1011.n124 G1011.n123 26.727
XR252 G1011.n124 G1011.n122 21.301
XR253 G1011.n114 G1011.n113 15
XR254 G1011.n136 G1011.n135 15
XR255 G1011.n152 G1011.n151 15
XR256 G1011.n126 G1011.n125 15
XR257 G1011.n129 G1011.n128 15
XR258 G1011.n160 G1011.n159 15
XR259 G1011.n158 G1011.n157 15
XR260 G1011.n150 G1011.n149 15
XR261 G1011.n144 G1011.n143 15
XR262 G1011.n142 G1011.n141 15
XR263 G1011.n134 G1011.n133 15
XR264 G1011.n106 G1011.n105 15
XR265 G1011.n108 G1011.n107 15
XR266 G1011.n116 G1011.n115 15
XR267 G1011.n181 G1011.n180 15
XR268 G1011.n174 G1011.n173 15
XR269 G1011.n185 G1011.n184 15
XR270 G1011.n190 G1011.n189 15
XR271 G1011.n161 G1011.n160 12.917
XR272 G1011.n153 G1011.n152 12.917
XR273 G1011.n145 G1011.n144 12.917
XR274 G1011.n137 G1011.n136 12.917
XR275 G1011.n106 G1011.n104 12.917
XR276 G1011.n114 G1011.n111 12.917
XR277 G1011.n122 G1011.n119 12.917
XR278 G1011.n230 G1011.n229 12.558
XR279 G1011.n284 G1011.n283 12.558
XR280 G1011.n300 G1011.n299 12.558
XR281 G1011.n316 G1011.n315 12.558
XR282 G1011.n332 G1011.n331 12.558
XR283 G1011.n348 G1011.n347 12.558
XR284 G1011.n364 G1011.n363 12.558
XR285 G1011.n380 G1011.n379 12.558
XR286 G1011.n396 G1011.n395 12.558
XR287 G1011.n412 G1011.n411 12.558
XR288 G1011.n430 G1011.n429 12.558
XR289 G1011.n448 G1011.n447 12.558
XR290 G1011.n464 G1011.n463 12.558
XR291 G1011.n480 G1011.n479 12.558
XR292 G1011.n496 G1011.n495 12.558
XR293 G1011.n512 G1011.n511 12.558
XR294 G1011.n528 G1011.n527 12.558
XR295 G1011.n544 G1011.n543 12.558
XR296 G1011.n560 G1011.n559 12.558
XR297 G1011.n573 G1011.n572 12.558
XR298 G1011.n212 G1011.n211 12.558
XR299 G1011.n242 G1011.n241 12.558
XR300 G1011.n233 G1011.n232 12.256
XR301 G1011.n215 G1011.n214 12.256
XR302 G1011.n287 G1011.n286 12.256
XR303 G1011.n303 G1011.n302 12.256
XR304 G1011.n319 G1011.n318 12.256
XR305 G1011.n335 G1011.n334 12.256
XR306 G1011.n351 G1011.n350 12.256
XR307 G1011.n367 G1011.n366 12.256
XR308 G1011.n383 G1011.n382 12.256
XR309 G1011.n399 G1011.n398 12.256
XR310 G1011.n415 G1011.n414 12.256
XR311 G1011.n433 G1011.n432 12.256
XR312 G1011.n451 G1011.n450 12.256
XR313 G1011.n467 G1011.n466 12.256
XR314 G1011.n483 G1011.n482 12.256
XR315 G1011.n499 G1011.n498 12.256
XR316 G1011.n515 G1011.n514 12.256
XR317 G1011.n531 G1011.n530 12.256
XR318 G1011.n547 G1011.n546 12.256
XR319 G1011.n563 G1011.n562 12.256
XR320 G1011.n576 G1011.n575 12.256
XR321 G1011.n245 G1011.n244 12.256
XR322 G1011.n182 G1011.n174 8.944
XR323 G1011.n182 G1011.n181 8.944
XR324 G1011.n184 G1011.n183 8.944
XR325 G1011.n122 G1011.n121 7.5
XR326 G1011.n133 G1011.n132 6.025
XR327 G1011.n167 G1011.n166 5.741
XR328 G1011.n210 G1011.n209 5.54
XR329 G1011.n117 G1011.n116 5.382
XR330 G1011.n118 G1011.n117 5.382
XR331 G1011.n129 G1011.n126 5.023
XR332 G1011.n162 G1011.n161 5.023
XR333 G1011.n141 G1011.n140 4.929
XR334 G1011.n179 G1011.n178 4.696
XR335 G1011.n192 G1011.n191 4.696
XR336 G1011.n109 G1011.n108 4.664
XR337 G1011.n110 G1011.n109 4.664
XR338 G1011.n50 G1011.n167 4.5
XR339 G1011.n0 G1011.n162 4.5
XR340 G1011.n172 G1011.n171 4.5
XR341 G1011.n196 G1011.n195 4.5
XR342 G1011.n187 G1011.n186 4.5
XR343 G1011.n160 G1011.n158 4.305
XR344 G1011.n154 G1011.n153 4.305
XR345 G1011.n173 G1011.n172 4.305
XR346 G1011.n186 G1011.n185 4.305
XR347 G1011.n28 G1011.n272 4.298
XR348 G1011.n134 G1011.n131 3.947
XR349 G1011.n149 G1011.n148 3.834
XR350 G1011.n165 G1011.n164 3.781
XR351 G1011.n152 G1011.n150 3.588
XR352 G1011.n146 G1011.n145 3.588
XR353 G1011.n2 G1011.n202 3.41
XR354 G1011.n49 G1011.n208 3.509
XR355 G1011.n198 G1011.n197 3.41
XR356 G1011.n142 G1011.n139 3.229
XR357 G1011.n139 G1011.n138 3.229
XR358 G1011.n144 G1011.n142 2.87
XR359 G1011.n138 G1011.n137 2.87
XR360 G1011.n157 G1011.n156 2.738
XR361 G1011.n150 G1011.n147 2.511
XR362 G1011.n147 G1011.n146 2.511
XR363 G1011.n1 G1011.n0 2.263
XR364 G1011.n1 G1011.n50 2.247
XR365 G1011.n1 G1011.n102 2.241
XR366 G1011.n136 G1011.n134 2.152
XR367 G1011.n104 G1011.n103 2.152
XR368 G1011.n158 G1011.n155 1.794
XR369 G1011.n155 G1011.n154 1.794
XR370 G1011.n289 G1011.n288 1.704
XR371 G1011.n305 G1011.n304 1.704
XR372 G1011.n321 G1011.n320 1.704
XR373 G1011.n337 G1011.n336 1.704
XR374 G1011.n353 G1011.n352 1.704
XR375 G1011.n369 G1011.n368 1.704
XR376 G1011.n385 G1011.n384 1.704
XR377 G1011.n401 G1011.n400 1.704
XR378 G1011.n417 G1011.n416 1.704
XR379 G1011.n435 G1011.n434 1.704
XR380 G1011.n453 G1011.n452 1.704
XR381 G1011.n469 G1011.n468 1.704
XR382 G1011.n485 G1011.n484 1.704
XR383 G1011.n501 G1011.n500 1.704
XR384 G1011.n517 G1011.n516 1.704
XR385 G1011.n533 G1011.n532 1.704
XR386 G1011.n549 G1011.n548 1.704
XR387 G1011.n565 G1011.n564 1.704
XR388 G1011.n578 G1011.n577 1.704
XR389 G1011.n585 G1011.n584 1.704
XR390 G1011.n247 G1011.n246 1.704
XR391 G1011.n128 G1011.n127 1.643
XR392 G1011 G1011.n587 1.635
XR393 G1011.n172 G1011.n100 1.467
XR394 G1011.n186 G1011.n99 1.467
XR395 G1011.n108 G1011.n106 1.435
XR396 G1011.n111 G1011.n110 1.435
XR397 G1011.n130 G1011.n129 1.076
XR398 G1011.n162 G1011.n130 1.076
XR399 G1011.n180 G1011.n179 1.076
XR400 G1011.n191 G1011.n190 1.076
XR401 G1011.n587 G1011.n234 1.014
XR402 G1011.n8 G1011.n580 0.857
XR403 G1011.n9 G1011.n567 0.857
XR404 G1011.n10 G1011.n551 0.857
XR405 G1011.n11 G1011.n535 0.857
XR406 G1011.n12 G1011.n519 0.857
XR407 G1011.n13 G1011.n503 0.857
XR408 G1011.n14 G1011.n487 0.857
XR409 G1011.n15 G1011.n471 0.857
XR410 G1011.n16 G1011.n455 0.857
XR411 G1011.n17 G1011.n437 0.857
XR412 G1011.n18 G1011.n419 0.857
XR413 G1011.n19 G1011.n403 0.857
XR414 G1011.n20 G1011.n387 0.857
XR415 G1011.n21 G1011.n371 0.857
XR416 G1011.n22 G1011.n355 0.857
XR417 G1011.n23 G1011.n339 0.857
XR418 G1011.n24 G1011.n323 0.857
XR419 G1011.n25 G1011.n307 0.857
XR420 G1011.n26 G1011.n291 0.857
XR421 G1011.n27 G1011.n275 0.857
XR422 G1011.n28 G1011.n248 0.856
XR423 G1011.n28 G1011.n273 0.856
XR424 G1011.n3 G1011.n249 0.856
XR425 G1011.n4 G1011.n254 0.856
XR426 G1011.n5 G1011.n259 0.856
XR427 G1011.n6 G1011.n264 0.856
XR428 G1011.n7 G1011.n269 0.856
XR429 G1011.n7 G1011.n271 0.856
XR430 G1011.n5 G1011.n262 0.856
XR431 G1011.n3 G1011.n252 0.856
XR432 G1011.n27 G1011.n290 0.856
XR433 G1011.n26 G1011.n306 0.856
XR434 G1011.n25 G1011.n322 0.856
XR435 G1011.n24 G1011.n338 0.856
XR436 G1011.n23 G1011.n354 0.856
XR437 G1011.n22 G1011.n370 0.856
XR438 G1011.n21 G1011.n386 0.856
XR439 G1011.n20 G1011.n402 0.856
XR440 G1011.n19 G1011.n418 0.856
XR441 G1011.n18 G1011.n436 0.856
XR442 G1011.n17 G1011.n454 0.856
XR443 G1011.n16 G1011.n470 0.856
XR444 G1011.n15 G1011.n486 0.856
XR445 G1011.n14 G1011.n502 0.856
XR446 G1011.n13 G1011.n518 0.856
XR447 G1011.n12 G1011.n534 0.856
XR448 G1011.n11 G1011.n550 0.856
XR449 G1011.n10 G1011.n566 0.856
XR450 G1011.n9 G1011.n579 0.856
XR451 G1011.n8 G1011.n586 0.856
XR452 G1011.n6 G1011.n267 0.856
XR453 G1011.n4 G1011.n257 0.856
XR454 G1011.n209 G1011.n49 0.746
XR455 G1011.n210 G1011.n198 1.007
XR456 G1011.n116 G1011.n114 0.717
XR457 G1011.n119 G1011.n118 0.717
XR458 G1011.n176 G1011.n175 0.717
XR459 G1011.n195 G1011.n194 0.717
XR460 G1011.n170 G1011.n169 0.589
XR461 G1011.n123 G1011.t107 0.506
XR462 G1011.n5 G1011.n258 0.448
XR463 G1011.n51 G1011.n201 0.432
XR464 G1011.n223 G1011.n222 0.429
XR465 G1011.n220 G1011.n219 0.429
XR466 G1011.n441 G1011.n440 0.429
XR467 G1011.n440 G1011.n439 0.429
XR468 G1011.n421 G1011.n420 0.429
XR469 G1011.n422 G1011.n421 0.429
XR470 G1011.n208 G1011.n207 0.429
XR471 G1011.n207 G1011.n206 0.429
XR472 G1011.n201 G1011.n200 0.429
XR473 G1011.n167 G1011.n165 0.358
XR474 G1011.n177 G1011.n176 0.358
XR475 G1011.n194 G1011.n193 0.358
XR476 G1011.n178 G1011.n177 0.326
XR477 G1011.n193 G1011.n192 0.326
XR478 G1011.n38 G1011.n18 0.262
XR479 G1011.n280 G1011.n278 0.241
XR480 G1011.n296 G1011.n294 0.241
XR481 G1011.n312 G1011.n310 0.241
XR482 G1011.n328 G1011.n326 0.241
XR483 G1011.n344 G1011.n342 0.241
XR484 G1011.n360 G1011.n358 0.241
XR485 G1011.n376 G1011.n374 0.241
XR486 G1011.n392 G1011.n390 0.241
XR487 G1011.n408 G1011.n406 0.241
XR488 G1011.n426 G1011.n424 0.241
XR489 G1011.n444 G1011.n442 0.241
XR490 G1011.n460 G1011.n458 0.241
XR491 G1011.n476 G1011.n474 0.241
XR492 G1011.n492 G1011.n490 0.241
XR493 G1011.n508 G1011.n506 0.241
XR494 G1011.n524 G1011.n522 0.241
XR495 G1011.n540 G1011.n538 0.241
XR496 G1011.n556 G1011.n554 0.241
XR497 G1011.n221 G1011.n216 0.241
XR498 G1011.n226 G1011.n224 0.241
XR499 G1011.n238 G1011.n236 0.241
XR500 G1011.n224 G1011.n223 0.214
XR501 G1011.n222 G1011.n221 0.214
XR502 G1011.n221 G1011.n220 0.214
XR503 G1011.n219 G1011.n218 0.214
XR504 G1011.n218 G1011.n217 0.214
XR505 G1011.n554 G1011.n552 0.214
XR506 G1011.n554 G1011.n553 0.214
XR507 G1011.n538 G1011.n536 0.214
XR508 G1011.n538 G1011.n537 0.214
XR509 G1011.n522 G1011.n520 0.214
XR510 G1011.n522 G1011.n521 0.214
XR511 G1011.n506 G1011.n504 0.214
XR512 G1011.n506 G1011.n505 0.214
XR513 G1011.n490 G1011.n488 0.214
XR514 G1011.n490 G1011.n489 0.214
XR515 G1011.n474 G1011.n472 0.214
XR516 G1011.n474 G1011.n473 0.214
XR517 G1011.n458 G1011.n456 0.214
XR518 G1011.n458 G1011.n457 0.214
XR519 G1011.n442 G1011.n438 0.214
XR520 G1011.n442 G1011.n441 0.214
XR521 G1011.n424 G1011.n422 0.214
XR522 G1011.n424 G1011.n423 0.214
XR523 G1011.n406 G1011.n404 0.214
XR524 G1011.n406 G1011.n405 0.214
XR525 G1011.n390 G1011.n388 0.214
XR526 G1011.n390 G1011.n389 0.214
XR527 G1011.n374 G1011.n372 0.214
XR528 G1011.n374 G1011.n373 0.214
XR529 G1011.n358 G1011.n356 0.214
XR530 G1011.n358 G1011.n357 0.214
XR531 G1011.n342 G1011.n340 0.214
XR532 G1011.n342 G1011.n341 0.214
XR533 G1011.n326 G1011.n324 0.214
XR534 G1011.n326 G1011.n325 0.214
XR535 G1011.n310 G1011.n308 0.214
XR536 G1011.n310 G1011.n309 0.214
XR537 G1011.n294 G1011.n292 0.214
XR538 G1011.n294 G1011.n293 0.214
XR539 G1011.n278 G1011.n276 0.214
XR540 G1011.n278 G1011.n277 0.214
XR541 G1011.n236 G1011.n235 0.214
XR542 G1011.n53 G1011.n52 0.19
XR543 G1011.n55 G1011.n54 0.19
XR544 G1011.n57 G1011.n56 0.19
XR545 G1011.n59 G1011.n58 0.19
XR546 G1011.n61 G1011.n60 0.19
XR547 G1011.n63 G1011.n62 0.19
XR548 G1011.n65 G1011.n64 0.19
XR549 G1011.n67 G1011.n66 0.19
XR550 G1011.n69 G1011.n68 0.19
XR551 G1011.n71 G1011.n70 0.19
XR552 G1011.n73 G1011.n72 0.19
XR553 G1011.n75 G1011.n74 0.19
XR554 G1011.n77 G1011.n76 0.19
XR555 G1011.n79 G1011.n78 0.19
XR556 G1011.n81 G1011.n80 0.19
XR557 G1011.n83 G1011.n82 0.19
XR558 G1011.n85 G1011.n84 0.19
XR559 G1011.n87 G1011.n86 0.19
XR560 G1011.n89 G1011.n88 0.19
XR561 G1011.n93 G1011.n92 0.19
XR562 G1011.n95 G1011.n94 0.19
XR563 G1011.n198 G1011.n97 0.113
XR564 G1011.n0 G1011.n124 20.061
XR565 G1011 G1011.n210 0.102
XR566 G1011.n587 G1011.n8 0.099
XR567 G1011.n197 G1011.n196 0.085
XR568 G1011.n4 G1011.n253 0.077
XR569 G1011.n35 G1011.n15 0.077
XR570 G1011.n39 G1011.n19 0.077
XR571 G1011.n6 G1011.n263 0.076
XR572 G1011.n7 G1011.n268 0.076
XR573 G1011.n29 G1011.n9 0.076
XR574 G1011.n30 G1011.n10 0.076
XR575 G1011.n31 G1011.n11 0.076
XR576 G1011.n32 G1011.n12 0.076
XR577 G1011.n33 G1011.n13 0.076
XR578 G1011.n34 G1011.n14 0.076
XR579 G1011.n36 G1011.n16 0.076
XR580 G1011.n37 G1011.n17 0.076
XR581 G1011.n40 G1011.n20 0.076
XR582 G1011.n41 G1011.n21 0.076
XR583 G1011.n42 G1011.n22 0.076
XR584 G1011.n43 G1011.n23 0.076
XR585 G1011.n44 G1011.n24 0.076
XR586 G1011.n45 G1011.n25 0.076
XR587 G1011.n46 G1011.n26 0.076
XR588 G1011.n47 G1011.n27 0.076
XR589 G1011.n48 G1011.n274 0.076
XR590 G1011.n271 G1011.n270 0.052
XR591 G1011.n262 G1011.n261 0.052
XR592 G1011.n252 G1011.n251 0.052
XR593 G1011.n257 G1011.n256 0.052
XR594 G1011.n267 G1011.n266 0.052
XR595 G1011.n586 G1011.n585 0.052
XR596 G1011.n579 G1011.n578 0.052
XR597 G1011.n566 G1011.n565 0.052
XR598 G1011.n550 G1011.n549 0.052
XR599 G1011.n534 G1011.n533 0.052
XR600 G1011.n518 G1011.n517 0.052
XR601 G1011.n502 G1011.n501 0.052
XR602 G1011.n486 G1011.n485 0.052
XR603 G1011.n470 G1011.n469 0.052
XR604 G1011.n454 G1011.n453 0.052
XR605 G1011.n436 G1011.n435 0.052
XR606 G1011.n418 G1011.n417 0.052
XR607 G1011.n402 G1011.n401 0.052
XR608 G1011.n386 G1011.n385 0.052
XR609 G1011.n370 G1011.n369 0.052
XR610 G1011.n354 G1011.n353 0.052
XR611 G1011.n338 G1011.n337 0.052
XR612 G1011.n322 G1011.n321 0.052
XR613 G1011.n306 G1011.n305 0.052
XR614 G1011.n290 G1011.n289 0.052
XR615 G1011.n248 G1011.n247 0.052
XR616 G1011.n246 G1011.n95 0.045
XR617 G1011.n94 G1011.n238 0.045
XR618 G1011.n234 G1011.n93 0.045
XR619 G1011.n92 G1011.n226 0.045
XR620 G1011.n584 G1011.n91 0.045
XR621 G1011.n216 G1011.n90 0.045
XR622 G1011.n577 G1011.n89 0.045
XR623 G1011.n88 G1011.n569 0.045
XR624 G1011.n564 G1011.n87 0.045
XR625 G1011.n86 G1011.n556 0.045
XR626 G1011.n548 G1011.n85 0.045
XR627 G1011.n84 G1011.n540 0.045
XR628 G1011.n532 G1011.n83 0.045
XR629 G1011.n82 G1011.n524 0.045
XR630 G1011.n516 G1011.n81 0.045
XR631 G1011.n80 G1011.n508 0.045
XR632 G1011.n500 G1011.n79 0.045
XR633 G1011.n78 G1011.n492 0.045
XR634 G1011.n484 G1011.n77 0.045
XR635 G1011.n76 G1011.n476 0.045
XR636 G1011.n468 G1011.n75 0.045
XR637 G1011.n74 G1011.n460 0.045
XR638 G1011.n452 G1011.n73 0.045
XR639 G1011.n72 G1011.n444 0.045
XR640 G1011.n434 G1011.n71 0.045
XR641 G1011.n70 G1011.n426 0.045
XR642 G1011.n416 G1011.n69 0.045
XR643 G1011.n68 G1011.n408 0.045
XR644 G1011.n400 G1011.n67 0.045
XR645 G1011.n66 G1011.n392 0.045
XR646 G1011.n384 G1011.n65 0.045
XR647 G1011.n64 G1011.n376 0.045
XR648 G1011.n368 G1011.n63 0.045
XR649 G1011.n62 G1011.n360 0.045
XR650 G1011.n352 G1011.n61 0.045
XR651 G1011.n60 G1011.n344 0.045
XR652 G1011.n336 G1011.n59 0.045
XR653 G1011.n58 G1011.n328 0.045
XR654 G1011.n320 G1011.n57 0.045
XR655 G1011.n56 G1011.n312 0.045
XR656 G1011.n304 G1011.n55 0.045
XR657 G1011.n54 G1011.n296 0.045
XR658 G1011.n288 G1011.n53 0.045
XR659 G1011.n52 G1011.n280 0.045
XR660 G1011.n49 G1011.n205 0.039
XR661 G1011.n202 G1011.n51 0.033
XR662 G1011.n204 G1011.n203 0.029
XR663 G1011.n50 G1011.n163 0.029
XR664 G1011.n205 G1011.n204 0.028
XR665 G1011.n50 G1011.n168 0.025
XR666 G1011.n2 G1011.n199 0.021
XR667 G1011.n171 G1011.n170 2.275
XR668 G1011.n196 G1011.n188 0.02
XR669 G1011.n171 G1011.n101 0.019
XR670 G1011.n187 G1011.n98 0.019
XR671 G1011.n274 G1011.n28 0.018
XR672 G1011.n272 G1011.n7 0.018
XR673 G1011.n263 G1011.n5 0.018
XR674 G1011.n253 G1011.n3 0.018
XR675 G1011.n197 G1011.n187 0.017
XR676 G1011.n203 G1011.n2 0.017
XR677 G1011.n27 G1011.n48 0.017
XR678 G1011.n26 G1011.n47 0.017
XR679 G1011.n25 G1011.n46 0.017
XR680 G1011.n24 G1011.n45 0.017
XR681 G1011.n23 G1011.n44 0.017
XR682 G1011.n22 G1011.n43 0.017
XR683 G1011.n21 G1011.n42 0.017
XR684 G1011.n20 G1011.n41 0.017
XR685 G1011.n19 G1011.n40 0.017
XR686 G1011.n18 G1011.n39 0.017
XR687 G1011.n17 G1011.n38 0.017
XR688 G1011.n16 G1011.n37 0.017
XR689 G1011.n15 G1011.n36 0.017
XR690 G1011.n14 G1011.n35 0.017
XR691 G1011.n13 G1011.n34 0.017
XR692 G1011.n12 G1011.n33 0.017
XR693 G1011.n11 G1011.n32 0.017
XR694 G1011.n10 G1011.n31 0.017
XR695 G1011.n9 G1011.n30 0.017
XR696 G1011.n8 G1011.n29 0.017
XR697 G1011.n268 G1011.n6 0.017
XR698 G1011.n258 G1011.n4 0.017
XR699 G1011.n169 G1011.n1 0.017
XR700 G1011.n97 G1011.n96 0.012
XR701 D6.n33 D6.t17 136.836
XR702 D6.n6 D6.t12 136.836
XR703 D6.n33 D6.t10 136.407
XR704 D6.n34 D6.t13 136.407
XR705 D6.n35 D6.t14 136.407
XR706 D6.n8 D6.t11 136.407
XR707 D6.n7 D6.t15 136.407
XR708 D6.n6 D6.t19 136.407
XR709 D6.n38 D6.n37 92.376
XR710 D6.n41 D6.n42 92.376
XR711 D6.n5 D6.t16 65.516
XR712 D6.n9 D6.t18 65.516
XR713 D6.n37 D6.t9 39.357
XR714 D6.n37 D6.t8 39.357
XR715 D6.n42 D6.t7 39.357
XR716 D6.n42 D6.t6 39.357
XR717 D6.n14 D6.n13 5.741
XR718 D6.n22 D6.n21 5.741
XR719 D6.n31 D6.n30 5.741
XR720 D6.n2 D6.n15 4.5
XR721 D6.n19 D6.n23 4.5
XR722 D6.n27 D6.n32 4.5
XR723 D6.n27 D6.n26 3.648
XR724 D6.n2 D6.n11 3.648
XR725 D6.n19 D6.n18 3.648
XR726 D6.n4 D6.n1 3.5
XR727 D6.n3 D6.n2 3.234
XR728 D6.n1 D6.n27 3.229
XR729 D6.n18 D6.n17 2.666
XR730 D6.n11 D6.n10 2.666
XR731 D6.n26 D6.n25 2.666
XR732 D6.n38 D6.n36 2.383
XR733 D6.n11 D6.t1 1.846
XR734 D6.n11 D6.t2 1.846
XR735 D6.n18 D6.t4 1.846
XR736 D6.n18 D6.t3 1.846
XR737 D6.n26 D6.t5 1.846
XR738 D6.n26 D6.t0 1.846
XR739 D6.n3 D6.n16 1.711
XR740 D6.n1 D6.n24 1.711
XR741 D6.n0 D6.n19 2.67
XR742 D6 D6.n40 1.084
XR743 D6.n4 D6.n39 0.856
XR744 D6.n35 D6.n34 0.429
XR745 D6.n34 D6.n33 0.429
XR746 D6.n7 D6.n6 0.429
XR747 D6.n8 D6.n7 0.429
XR748 D6.n15 D6.n14 0.358
XR749 D6.n13 D6.n12 0.358
XR750 D6.n23 D6.n22 0.358
XR751 D6.n21 D6.n20 0.358
XR752 D6.n32 D6.n31 0.358
XR753 D6.n30 D6.n29 0.358
XR754 D6.n9 D6.n8 0.349
XR755 D6.n40 D6.n41 0.056
XR756 D6.n39 D6.n38 0.056
XR757 D6.n36 D6.n5 1.619
XR758 D6.n9 D6.n41 4
XR759 D6.n5 D6.n35 0.349
XR760 D6.n1 D6.n0 0.1
XR761 D6.n0 D6.n3 0.09
XR762 D6 D6.n4 0.048
XR763 D6.n27 D6.n28 0.041
XR764 D5.n0 D5.n8 32.825
XR765 D5.n11 D5.n10 32.371
XR766 D5.n8 D5.t2 27.695
XR767 D5.n8 D5.t0 27.695
XR768 D5.n10 D5.t1 27.695
XR769 D5.n10 D5.t3 27.695
XR770 D5.n33 D5.n32 6.05
XR771 D5.n27 D5.n29 6
XR772 D5.n29 D5.n28 3.947
XR773 D5.n32 D5.n31 3.947
XR774 D5.n35 D5.n34 3.171
XR775 D5.n18 D5.n17 3.171
XR776 D5.n25 D5.n24 3.171
XR777 D5.n16 D5.n15 3.171
XR778 D5.n14 D5.n13 3.171
XR779 D5.n33 D5.n35 4.419
XR780 D5.n30 D5.n25 4.419
XR781 D5.n23 D5.n22 1.882
XR782 D5.n18 D5.t5 1.846
XR783 D5.n18 D5.t6 1.846
XR784 D5.n21 D5.t7 1.846
XR785 D5.n21 D5.t11 1.846
XR786 D5.n25 D5.t12 1.846
XR787 D5.n25 D5.t14 1.846
XR788 D5.n16 D5.t13 1.846
XR789 D5.n16 D5.t15 1.846
XR790 D5.n14 D5.t8 1.846
XR791 D5.n14 D5.t9 1.846
XR792 D5.n35 D5.t10 1.846
XR793 D5.n35 D5.t4 1.846
XR794 D5.n6 D5.n5 1.748
XR795 D5.n6 D5.n18 6.114
XR796 D5.n4 D5.n16 6.114
XR797 D5.n3 D5.n14 6.114
XR798 D5.n27 D5.n26 1.604
XR799 D5.n21 D5.n20 1.516
XR800 D5.n19 D5.n23 1.512
XR801 D5 D5.n3 1.446
XR802 D5.n1 D5.n19 1.271
XR803 D5.n7 D5.n33 1.131
XR804 D5.n2 D5.n30 1.131
XR805 D5.n22 D5.n21 1.016
XR806 D5.n0 D5.n12 0.856
XR807 D5.n0 D5.n9 0.856
XR808 D5 D5.n0 0.708
XR809 D5.n4 D5.n2 0.099
XR810 D5.n7 D5.n4 0.092
XR811 D5.n3 D5.n7 0.091
XR812 D5.n1 D5.n6 0.09
XR813 D5.n2 D5.n1 0.084
XR814 D5.n12 D5.n11 0.052
XR815 D5.n30 D5.n27 0.05
XR816 D9.n154 D9.t15 136.6
XR817 D9.n152 D9.t16 136.6
XR818 D9.n147 D9.t10 136.407
XR819 D9.n148 D9.t8 136.407
XR820 D9.n151 D9.t6 136.407
XR821 D9.n152 D9.t17 136.407
XR822 D9.n153 D9.t12 136.407
XR823 D9.n154 D9.t14 136.407
XR824 D9.n115 D9.t3 122.45
XR825 D9.n44 D9.t5 122.45
XR826 D9.n42 D9.t5 111.965
XR827 D9.n140 D9.n150 92.998
XR828 D9.n143 D9.n155 92.998
XR829 D9.n131 D9.n130 49.396
XR830 D9.n60 D9.n59 49.396
XR831 D9.n124 D9.n123 42.81
XR832 D9.n53 D9.n52 42.81
XR833 D9.n150 D9.t13 39.357
XR834 D9.n150 D9.t9 39.357
XR835 D9.n155 D9.t11 39.357
XR836 D9.n155 D9.t7 39.357
XR837 D9.n45 D9.n44 22.786
XR838 D9.n116 D9.n115 22.786
XR839 D9.n115 D9.n114 19.893
XR840 D9.n44 D9.n43 19.893
XR841 D9.n132 D9.n131 15
XR842 D9.n125 D9.n124 15
XR843 D9.n134 D9.n133 15
XR844 D9.n122 D9.n121 15
XR845 D9.n54 D9.n53 15
XR846 D9.n61 D9.n60 15
XR847 D9.n51 D9.n50 15
XR848 D9.n63 D9.n62 15
XR849 D9.n135 D9.n134 12.917
XR850 D9.n64 D9.n63 12.917
XR851 D9.n114 D9.n113 7.5
XR852 D9.n43 D9.n42 7.5
XR853 D9.n85 D9.n83 6.614
XR854 D9.n101 D9.n99 6.614
XR855 D9 D9.n137 5.428
XR856 D9.n132 D9.n129 5.382
XR857 D9.n129 D9.n128 5.382
XR858 D9.n61 D9.n58 5.382
XR859 D9.n58 D9.n57 5.382
XR860 D9.n82 D9.n80 4.664
XR861 D9.n98 D9.n96 4.664
XR862 D9.n126 D9.n125 4.664
XR863 D9.n136 D9.n126 4.664
XR864 D9.n55 D9.n54 4.664
XR865 D9.n65 D9.n55 4.664
XR866 D9.n10 D9.n82 4.5
XR867 D9.n9 D9.n36 4.5
XR868 D9.n12 D9.n29 4.5
XR869 D9.n13 D9.n98 4.5
XR870 D9.n16 D9.n136 4.5
XR871 D9.n15 D9.n24 4.5
XR872 D9.n7 D9.n71 4.5
XR873 D9.n8 D9.n65 4.5
XR874 D9.n36 D9.n34 3.947
XR875 D9.n29 D9.n27 3.947
XR876 D9.n24 D9.n22 3.947
XR877 D9.n71 D9.n69 3.947
XR878 D9.n87 D9.n86 3.882
XR879 D9.n103 D9.n102 3.882
XR880 D9.n69 D9.n68 3.695
XR881 D9.n22 D9.n21 3.695
XR882 D9.n138 D9.n146 2.879
XR883 D9.n144 D9.n149 2.878
XR884 D9.n36 D9.n35 2.152
XR885 D9.n29 D9.n28 2.152
XR886 D9.n24 D9.n23 2.152
XR887 D9.n71 D9.n70 2.152
XR888 D9.n85 D9.t0 1.846
XR889 D9.n85 D9.t1 1.846
XR890 D9.n101 D9.t4 1.846
XR891 D9.n101 D9.t2 1.846
XR892 D9.n6 D9.n14 1.704
XR893 D9.n5 D9.n17 1.704
XR894 D9.n2 D9.n11 1.704
XR895 D9.n0 D9.n18 1.704
XR896 D9.n1 D9.n31 1.703
XR897 D9.n6 D9.n90 1.703
XR898 D9.n5 D9.n106 1.703
XR899 D9.n0 D9.n72 1.703
XR900 D9.n1 D9.n30 1.702
XR901 D9.n6 D9.n89 1.702
XR902 D9.n5 D9.n107 1.702
XR903 D9.n0 D9.n73 1.702
XR904 D9.n11 D9.n10 1.5
XR905 D9.n1 D9.n9 3.204
XR906 D9.n4 D9.n12 3.204
XR907 D9.n14 D9.n13 1.5
XR908 D9.n17 D9.n16 1.5
XR909 D9.n3 D9.n15 3.204
XR910 D9.n0 D9.n7 3.204
XR911 D9.n18 D9.n8 1.5
XR912 D9.n82 D9.n81 1.435
XR913 D9.n98 D9.n97 1.435
XR914 D9.n125 D9.n122 1.435
XR915 D9.n136 D9.n135 1.435
XR916 D9.n54 D9.n51 1.435
XR917 D9.n65 D9.n64 1.435
XR918 D9.n141 D9.n142 0.856
XR919 D9.n134 D9.n132 0.717
XR920 D9.n128 D9.n127 0.717
XR921 D9.n63 D9.n61 0.717
XR922 D9.n57 D9.n56 0.717
XR923 D9.n4 D9.n2 0.355
XR924 D9.n86 D9.n85 0.302
XR925 D9.n102 D9.n101 0.302
XR926 D9.n85 D9.n84 0.207
XR927 D9.n101 D9.n100 0.207
XR928 D9.n153 D9.n154 0.193
XR929 D9.n147 D9.n148 0.193
XR930 D9.n151 D9.n152 0.193
XR931 D9 D9.n141 0.114
XR932 D9.n146 D9.n151 0.099
XR933 D9.n149 D9.n153 0.096
XR934 D9.n146 D9.n147 0.094
XR935 D9.n1 D9.n74 0.076
XR936 D9.n3 D9.n105 0.076
XR937 D9.n48 D9.n47 0.072
XR938 D9.n119 D9.n118 0.072
XR939 D9.n142 D9.n143 0.056
XR940 D9.n143 D9.n145 0.052
XR941 D9.n140 D9.n139 0.052
XR942 D9.n47 D9.n46 0.04
XR943 D9.n118 D9.n117 0.04
XR944 D9.n18 D9.n38 0.035
XR945 D9.n17 D9.n109 0.035
XR946 D9.n14 D9.n92 0.035
XR947 D9.n11 D9.n76 0.035
XR948 D9.n49 D9.n48 0.025
XR949 D9.n88 D9.n87 0.025
XR950 D9.n104 D9.n103 0.025
XR951 D9.n120 D9.n119 0.025
XR952 D9.n139 D9.n144 0.025
XR953 D9.n145 D9.n138 0.025
XR954 D9.n8 D9.n41 0.018
XR955 D9.n10 D9.n79 0.018
XR956 D9.n13 D9.n95 0.018
XR957 D9.n16 D9.n112 0.018
XR958 D9.n7 D9.n67 0.017
XR959 D9.n9 D9.n33 0.017
XR960 D9.n12 D9.n26 0.017
XR961 D9.n15 D9.n20 0.017
XR962 D9.n41 D9.n40 0.015
XR963 D9.n79 D9.n78 0.015
XR964 D9.n95 D9.n94 0.015
XR965 D9.n112 D9.n111 0.015
XR966 D9.n67 D9.n66 0.012
XR967 D9.n33 D9.n32 0.012
XR968 D9.n26 D9.n25 0.012
XR969 D9.n20 D9.n19 0.012
XR970 D9.n16 D9.n120 0.007
XR971 D9.n13 D9.n104 0.007
XR972 D9.n10 D9.n88 0.007
XR973 D9.n8 D9.n49 0.007
XR974 D9.n40 D9.n39 0.006
XR975 D9.n78 D9.n77 0.006
XR976 D9.n76 D9.n75 0.006
XR977 D9.n94 D9.n93 0.006
XR978 D9.n92 D9.n91 0.006
XR979 D9.n111 D9.n110 0.006
XR980 D9.n109 D9.n108 0.006
XR981 D9.n38 D9.n37 0.006
XR982 D9.n141 D9.n140 1.287
XR983 D9.n2 D9.n1 0.016
XR984 D9.n74 D9.n0 0.012
XR985 D9.n105 D9.n6 0.008
XR986 D9.n137 D9.n5 0.008
XR987 D9.n6 D9.n4 0.008
XR988 D9.n5 D9.n3 0.008
XR989 D9.n46 D9.n45 0.005
XR990 D9.n117 D9.n116 0.005
XR991 G3.n1 G3.t6 843.93
XR992 G3.n1 G3.t1 843.501
XR993 G3.n1 G3.t2 843.501
XR994 G3.n0 G3.t4 843.501
XR995 G3.n0 G3.t5 843.501
XR996 G3.n0 G3.t3 772.29
XR997 G3.n0 G3.t0 7.354
XR998 G3.n1 G3.n0 1.475
XR999 Vref.n36 Vref.n0 9.09
XR1000 Vref.n22 Vref.n21 6.614
XR1001 Vref.n7 Vref.n6 6.614
XR1002 Vref.n22 Vref.n20 6.489
XR1003 Vref.n7 Vref.n5 6.489
XR1004 Vref.n8 Vref.n7 6.208
XR1005 Vref.n4 Vref.n22 6.208
XR1006 Vref.n7 Vref.t1 5.539
XR1007 Vref.n7 Vref.t0 5.539
XR1008 Vref.n22 Vref.t3 5.539
XR1009 Vref.n22 Vref.t2 5.539
XR1010 Vref.n8 Vref.n11 4.5
XR1011 Vref.n14 Vref.n17 4.5
XR1012 Vref.n28 Vref.n32 4.5
XR1013 Vref.n4 Vref.n25 4.5
XR1014 Vref.n17 Vref.n15 3.947
XR1015 Vref.n32 Vref.n30 3.947
XR1016 Vref.n11 Vref.n9 3.229
XR1017 Vref.n25 Vref.n23 3.229
XR1018 Vref.n11 Vref.n10 2.87
XR1019 Vref.n25 Vref.n24 2.87
XR1020 Vref.n17 Vref.n16 2.152
XR1021 Vref.n32 Vref.n31 2.152
XR1022 Vref.n0 Vref.n35 1.704
XR1023 Vref.n1 Vref.n26 1.704
XR1024 Vref.n0 Vref.n3 1.704
XR1025 Vref.n0 Vref.n8 3.208
XR1026 Vref.n1 Vref.n2 1.704
XR1027 Vref.n3 Vref.n14 1.5
XR1028 Vref.n2 Vref.n28 1.5
XR1029 Vref Vref.n36 1.214
XR1030 Vref.n36 Vref.t4 0.265
XR1031 Vref.n3 Vref.n12 0.031
XR1032 Vref.n2 Vref.n33 0.031
XR1033 Vref.n14 Vref.n18 0.027
XR1034 Vref.n28 Vref.n29 0.027
XR1035 Vref.n12 Vref.n13 0.009
XR1036 Vref.n33 Vref.n34 0.009
XR1037 Vref.n1 Vref.n4 3.208
XR1038 Vref.n0 Vref.n1 0.099
XR1039 Vref.n3 Vref.n19 0.036
XR1040 Vref.n2 Vref.n27 0.036
XR1041 D1011.n10 D1011.t3 517.997
XR1042 D1011.n12 D1011.t4 482
XR1043 D1011.n506 D1011.n505 152
XR1044 D1011.n495 D1011.n494 152
XR1045 D1011.n484 D1011.n483 152
XR1046 D1011.n473 D1011.n472 152
XR1047 D1011.n462 D1011.n461 152
XR1048 D1011.n5 D1011.n451 152
XR1049 D1011.n6 D1011.n438 152
XR1050 D1011.n428 D1011.n427 152
XR1051 D1011.n417 D1011.n416 152
XR1052 D1011.n406 D1011.n405 152
XR1053 D1011.n404 D1011.n403 152
XR1054 D1011.n413 D1011.n412 152
XR1055 D1011.n415 D1011.n414 152
XR1056 D1011.n424 D1011.n423 152
XR1057 D1011.n426 D1011.n425 152
XR1058 D1011.n435 D1011.n434 152
XR1059 D1011.n437 D1011.n436 152
XR1060 D1011.n6 D1011.n444 152
XR1061 D1011.n5 D1011.n450 152
XR1062 D1011.n453 D1011.n452 152
XR1063 D1011.n460 D1011.n459 152
XR1064 D1011.n464 D1011.n463 152
XR1065 D1011.n471 D1011.n470 152
XR1066 D1011.n475 D1011.n474 152
XR1067 D1011.n482 D1011.n481 152
XR1068 D1011.n486 D1011.n485 152
XR1069 D1011.n493 D1011.n492 152
XR1070 D1011.n497 D1011.n496 152
XR1071 D1011.n504 D1011.n503 152
XR1072 D1011.n90 D1011.n89 152
XR1073 D1011.n101 D1011.n100 152
XR1074 D1011.n112 D1011.n111 152
XR1075 D1011.n4 D1011.n122 152
XR1076 D1011.n3 D1011.n135 152
XR1077 D1011.n146 D1011.n145 152
XR1078 D1011.n157 D1011.n156 152
XR1079 D1011.n168 D1011.n167 152
XR1080 D1011.n179 D1011.n178 152
XR1081 D1011.n190 D1011.n189 152
XR1082 D1011.n88 D1011.n87 152
XR1083 D1011.n99 D1011.n98 152
XR1084 D1011.n110 D1011.n109 152
XR1085 D1011.n121 D1011.n120 152
XR1086 D1011.n137 D1011.n136 152
XR1087 D1011.n148 D1011.n147 152
XR1088 D1011.n159 D1011.n158 152
XR1089 D1011.n170 D1011.n169 152
XR1090 D1011.n181 D1011.n180 152
XR1091 D1011.n97 D1011.n96 152
XR1092 D1011.n108 D1011.n107 152
XR1093 D1011.n119 D1011.n118 152
XR1094 D1011.n4 D1011.n128 152
XR1095 D1011.n3 D1011.n134 152
XR1096 D1011.n144 D1011.n143 152
XR1097 D1011.n155 D1011.n154 152
XR1098 D1011.n166 D1011.n165 152
XR1099 D1011.n177 D1011.n176 152
XR1100 D1011.n188 D1011.n187 152
XR1101 D1011.n74 D1011.t2 122.45
XR1102 D1011.n390 D1011.t1 122.45
XR1103 D1011.n72 D1011.t2 111.965
XR1104 D1011.n552 D1011.n551 76
XR1105 D1011.n236 D1011.n235 76
XR1106 D1011.n26 D1011.t0 62.054
XR1107 D1011.n525 D1011.n524 49.396
XR1108 D1011.n544 D1011.n543 49.396
XR1109 D1011.n383 D1011.n382 49.396
XR1110 D1011.n209 D1011.n208 49.396
XR1111 D1011.n228 D1011.n227 49.396
XR1112 D1011.n67 D1011.n66 49.396
XR1113 D1011.n517 D1011.n516 42.81
XR1114 D1011.n536 D1011.n535 42.81
XR1115 D1011.n375 D1011.n374 42.81
XR1116 D1011.n201 D1011.n200 42.81
XR1117 D1011.n220 D1011.n219 42.81
XR1118 D1011.n59 D1011.n58 42.81
XR1119 D1011.n318 D1011.n317 36.224
XR1120 D1011.n501 D1011.n500 36.224
XR1121 D1011.n367 D1011.n366 36.224
XR1122 D1011.n267 D1011.n266 36.224
XR1123 D1011.n185 D1011.n184 36.224
XR1124 D1011.n51 D1011.n50 36.224
XR1125 D1011.n326 D1011.n325 29.637
XR1126 D1011.n490 D1011.n489 29.637
XR1127 D1011.n359 D1011.n358 29.637
XR1128 D1011.n275 D1011.n274 29.637
XR1129 D1011.n174 D1011.n173 29.637
XR1130 D1011.n43 D1011.n42 29.637
XR1131 D1011.n334 D1011.n333 23.051
XR1132 D1011.n479 D1011.n478 23.051
XR1133 D1011.n410 D1011.n409 23.051
XR1134 D1011.n283 D1011.n282 23.051
XR1135 D1011.n163 D1011.n162 23.051
XR1136 D1011.n94 D1011.n93 23.051
XR1137 D1011.n75 D1011.n74 22.786
XR1138 D1011.n391 D1011.n390 22.786
XR1139 D1011.n390 D1011.n389 19.893
XR1140 D1011.n74 D1011.n73 19.893
XR1141 D1011.n342 D1011.n341 16.465
XR1142 D1011.n468 D1011.n467 16.465
XR1143 D1011.n421 D1011.n420 16.465
XR1144 D1011.n291 D1011.n290 16.465
XR1145 D1011.n152 D1011.n151 16.465
XR1146 D1011.n105 D1011.n104 16.465
XR1147 D1011.n20 D1011.n19 15
XR1148 D1011.n14 D1011.n13 15
XR1149 D1011.n384 D1011.n383 15
XR1150 D1011.n376 D1011.n375 15
XR1151 D1011.n368 D1011.n367 15
XR1152 D1011.n360 D1011.n359 15
XR1153 D1011.n411 D1011.n410 15
XR1154 D1011.n422 D1011.n421 15
XR1155 D1011.n433 D1011.n432 15
XR1156 D1011.n443 D1011.n442 15
XR1157 D1011.n449 D1011.n448 15
XR1158 D1011.n458 D1011.n457 15
XR1159 D1011.n469 D1011.n468 15
XR1160 D1011.n480 D1011.n479 15
XR1161 D1011.n491 D1011.n490 15
XR1162 D1011.n502 D1011.n501 15
XR1163 D1011.n537 D1011.n536 15
XR1164 D1011.n545 D1011.n544 15
XR1165 D1011.n526 D1011.n525 15
XR1166 D1011.n518 D1011.n517 15
XR1167 D1011.n319 D1011.n318 15
XR1168 D1011.n327 D1011.n326 15
XR1169 D1011.n335 D1011.n334 15
XR1170 D1011.n343 D1011.n342 15
XR1171 D1011.n351 D1011.n350 15
XR1172 D1011.n312 D1011.n311 15
XR1173 D1011.n582 D1011.n581 15
XR1174 D1011.n381 D1011.n380 15
XR1175 D1011.n373 D1011.n372 15
XR1176 D1011.n365 D1011.n364 15
XR1177 D1011.n357 D1011.n356 15
XR1178 D1011.n408 D1011.n407 15
XR1179 D1011.n419 D1011.n418 15
XR1180 D1011.n430 D1011.n429 15
XR1181 D1011.n440 D1011.n439 15
XR1182 D1011.n446 D1011.n445 15
XR1183 D1011.n455 D1011.n454 15
XR1184 D1011.n466 D1011.n465 15
XR1185 D1011.n477 D1011.n476 15
XR1186 D1011.n488 D1011.n487 15
XR1187 D1011.n499 D1011.n498 15
XR1188 D1011.n534 D1011.n533 15
XR1189 D1011.n542 D1011.n541 15
XR1190 D1011.n523 D1011.n522 15
XR1191 D1011.n515 D1011.n514 15
XR1192 D1011.n321 D1011.n320 15
XR1193 D1011.n329 D1011.n328 15
XR1194 D1011.n337 D1011.n336 15
XR1195 D1011.n345 D1011.n344 15
XR1196 D1011.n353 D1011.n352 15
XR1197 D1011.n309 D1011.n308 15
XR1198 D1011.n579 D1011.n578 15
XR1199 D1011.n33 D1011.n32 15
XR1200 D1011.n261 D1011.n260 15
XR1201 D1011.n300 D1011.n299 15
XR1202 D1011.n292 D1011.n291 15
XR1203 D1011.n284 D1011.n283 15
XR1204 D1011.n276 D1011.n275 15
XR1205 D1011.n268 D1011.n267 15
XR1206 D1011.n202 D1011.n201 15
XR1207 D1011.n210 D1011.n209 15
XR1208 D1011.n229 D1011.n228 15
XR1209 D1011.n221 D1011.n220 15
XR1210 D1011.n186 D1011.n185 15
XR1211 D1011.n175 D1011.n174 15
XR1212 D1011.n164 D1011.n163 15
XR1213 D1011.n153 D1011.n152 15
XR1214 D1011.n142 D1011.n141 15
XR1215 D1011.n133 D1011.n132 15
XR1216 D1011.n127 D1011.n126 15
XR1217 D1011.n117 D1011.n116 15
XR1218 D1011.n106 D1011.n105 15
XR1219 D1011.n95 D1011.n94 15
XR1220 D1011.n44 D1011.n43 15
XR1221 D1011.n52 D1011.n51 15
XR1222 D1011.n60 D1011.n59 15
XR1223 D1011.n68 D1011.n67 15
XR1224 D1011.n30 D1011.n29 15
XR1225 D1011.n258 D1011.n257 15
XR1226 D1011.n65 D1011.n64 15
XR1227 D1011.n57 D1011.n56 15
XR1228 D1011.n49 D1011.n48 15
XR1229 D1011.n41 D1011.n40 15
XR1230 D1011.n92 D1011.n91 15
XR1231 D1011.n103 D1011.n102 15
XR1232 D1011.n114 D1011.n113 15
XR1233 D1011.n124 D1011.n123 15
XR1234 D1011.n130 D1011.n129 15
XR1235 D1011.n139 D1011.n138 15
XR1236 D1011.n150 D1011.n149 15
XR1237 D1011.n161 D1011.n160 15
XR1238 D1011.n172 D1011.n171 15
XR1239 D1011.n183 D1011.n182 15
XR1240 D1011.n218 D1011.n217 15
XR1241 D1011.n226 D1011.n225 15
XR1242 D1011.n207 D1011.n206 15
XR1243 D1011.n199 D1011.n198 15
XR1244 D1011.n270 D1011.n269 15
XR1245 D1011.n278 D1011.n277 15
XR1246 D1011.n286 D1011.n285 15
XR1247 D1011.n294 D1011.n293 15
XR1248 D1011.n302 D1011.n301 15
XR1249 D1011.n577 D1011.n576 13.878
XR1250 D1011.n28 D1011.n27 13.878
XR1251 D1011.n354 D1011.n353 12.917
XR1252 D1011.n346 D1011.n345 12.917
XR1253 D1011.n338 D1011.n337 12.917
XR1254 D1011.n330 D1011.n329 12.917
XR1255 D1011.n322 D1011.n321 12.917
XR1256 D1011.n523 D1011.n521 12.917
XR1257 D1011.n531 D1011.n529 12.917
XR1258 D1011.n550 D1011.n548 12.917
XR1259 D1011.n542 D1011.n540 12.917
XR1260 D1011.n534 D1011.n532 12.917
XR1261 D1011.n365 D1011.n363 12.917
XR1262 D1011.n373 D1011.n371 12.917
XR1263 D1011.n381 D1011.n379 12.917
XR1264 D1011.n389 D1011.n387 12.917
XR1265 D1011.n303 D1011.n302 12.917
XR1266 D1011.n295 D1011.n294 12.917
XR1267 D1011.n287 D1011.n286 12.917
XR1268 D1011.n279 D1011.n278 12.917
XR1269 D1011.n271 D1011.n270 12.917
XR1270 D1011.n207 D1011.n205 12.917
XR1271 D1011.n215 D1011.n213 12.917
XR1272 D1011.n234 D1011.n232 12.917
XR1273 D1011.n226 D1011.n224 12.917
XR1274 D1011.n218 D1011.n216 12.917
XR1275 D1011.n49 D1011.n47 12.917
XR1276 D1011.n57 D1011.n55 12.917
XR1277 D1011.n65 D1011.n63 12.917
XR1278 D1011.n73 D1011.n71 12.917
XR1279 D1011.n551 D1011.n531 12.2
XR1280 D1011.n551 D1011.n550 12.2
XR1281 D1011.n235 D1011.n215 12.2
XR1282 D1011.n235 D1011.n234 12.2
XR1283 D1011.n350 D1011.n349 9.879
XR1284 D1011.n457 D1011.n456 9.879
XR1285 D1011.n432 D1011.n431 9.879
XR1286 D1011.n299 D1011.n298 9.879
XR1287 D1011.n141 D1011.n140 9.879
XR1288 D1011.n116 D1011.n115 9.879
XR1289 D1011.n13 D1011.n12 8.944
XR1290 D1011.n389 D1011.n388 7.5
XR1291 D1011.n550 D1011.n549 7.5
XR1292 D1011.n531 D1011.n530 7.5
XR1293 D1011.n73 D1011.n72 7.5
XR1294 D1011.n234 D1011.n233 7.5
XR1295 D1011.n215 D1011.n214 7.5
XR1296 D1011.n2 D1011.n577 5.741
XR1297 D1011.n582 D1011.n579 5.741
XR1298 D1011.n312 D1011.n309 5.741
XR1299 D1011.n355 D1011.n354 5.741
XR1300 D1011.n449 D1011.n446 5.741
XR1301 D1011.n443 D1011.n440 5.741
XR1302 D1011.n35 D1011.n28 5.741
XR1303 D1011.n33 D1011.n30 5.741
XR1304 D1011.n261 D1011.n258 5.741
XR1305 D1011.n304 D1011.n303 5.741
XR1306 D1011.n133 D1011.n130 5.741
XR1307 D1011.n127 D1011.n124 5.741
XR1308 D1011.n527 D1011.n526 5.382
XR1309 D1011.n528 D1011.n527 5.382
XR1310 D1011.n547 D1011.n546 5.382
XR1311 D1011.n546 D1011.n545 5.382
XR1312 D1011.n385 D1011.n384 5.382
XR1313 D1011.n386 D1011.n385 5.382
XR1314 D1011.n211 D1011.n210 5.382
XR1315 D1011.n212 D1011.n211 5.382
XR1316 D1011.n231 D1011.n230 5.382
XR1317 D1011.n230 D1011.n229 5.382
XR1318 D1011.n69 D1011.n68 5.382
XR1319 D1011.n70 D1011.n69 5.382
XR1320 D1011.n353 D1011.n351 5.023
XR1321 D1011.n347 D1011.n346 5.023
XR1322 D1011.n458 D1011.n455 5.023
XR1323 D1011.n433 D1011.n430 5.023
XR1324 D1011.n302 D1011.n300 5.023
XR1325 D1011.n296 D1011.n295 5.023
XR1326 D1011.n142 D1011.n139 5.023
XR1327 D1011.n117 D1011.n114 5.023
XR1328 D1011.n22 D1011.n21 4.696
XR1329 D1011.n519 D1011.n518 4.664
XR1330 D1011.n520 D1011.n519 4.664
XR1331 D1011.n539 D1011.n538 4.664
XR1332 D1011.n538 D1011.n537 4.664
XR1333 D1011.n377 D1011.n376 4.664
XR1334 D1011.n378 D1011.n377 4.664
XR1335 D1011.n203 D1011.n202 4.664
XR1336 D1011.n204 D1011.n203 4.664
XR1337 D1011.n223 D1011.n222 4.664
XR1338 D1011.n222 D1011.n221 4.664
XR1339 D1011.n61 D1011.n60 4.664
XR1340 D1011.n62 D1011.n61 4.664
XR1341 D1011.n18 D1011.n17 4.585
XR1342 D1011.n16 D1011.n15 4.5
XR1343 D1011.n307 D1011.n355 4.5
XR1344 D1011.n39 D1011.n304 4.5
XR1345 D1011.n15 D1011.n14 4.305
XR1346 D1011.n345 D1011.n343 4.305
XR1347 D1011.n339 D1011.n338 4.305
XR1348 D1011.n469 D1011.n466 4.305
XR1349 D1011.n422 D1011.n419 4.305
XR1350 D1011.n294 D1011.n292 4.305
XR1351 D1011.n288 D1011.n287 4.305
XR1352 D1011.n153 D1011.n150 4.305
XR1353 D1011.n106 D1011.n103 4.305
XR1354 D1011.n319 D1011.n316 3.947
XR1355 D1011.n316 D1011.n315 3.947
XR1356 D1011.n503 D1011.n502 3.947
XR1357 D1011.n369 D1011.n368 3.947
XR1358 D1011.n370 D1011.n369 3.947
XR1359 D1011.n268 D1011.n265 3.947
XR1360 D1011.n265 D1011.n264 3.947
XR1361 D1011.n187 D1011.n186 3.947
XR1362 D1011.n53 D1011.n52 3.947
XR1363 D1011.n54 D1011.n53 3.947
XR1364 D1011.n337 D1011.n335 3.588
XR1365 D1011.n331 D1011.n330 3.588
XR1366 D1011.n480 D1011.n477 3.588
XR1367 D1011.n411 D1011.n408 3.588
XR1368 D1011.n286 D1011.n284 3.588
XR1369 D1011.n280 D1011.n279 3.588
XR1370 D1011.n164 D1011.n161 3.588
XR1371 D1011.n95 D1011.n92 3.588
XR1372 D1011.n8 D1011.n18 3.41
XR1373 D1011.n581 D1011.n580 3.293
XR1374 D1011.n311 D1011.n310 3.293
XR1375 D1011.n448 D1011.n447 3.293
XR1376 D1011.n442 D1011.n441 3.293
XR1377 D1011.n32 D1011.n31 3.293
XR1378 D1011.n260 D1011.n259 3.293
XR1379 D1011.n132 D1011.n131 3.293
XR1380 D1011.n126 D1011.n125 3.293
XR1381 D1011.n327 D1011.n324 3.229
XR1382 D1011.n324 D1011.n323 3.229
XR1383 D1011.n492 D1011.n491 3.229
XR1384 D1011.n361 D1011.n360 3.229
XR1385 D1011.n362 D1011.n361 3.229
XR1386 D1011.n276 D1011.n273 3.229
XR1387 D1011.n273 D1011.n272 3.229
XR1388 D1011.n176 D1011.n175 3.229
XR1389 D1011.n45 D1011.n44 3.229
XR1390 D1011.n46 D1011.n45 3.229
XR1391 D1011.n329 D1011.n327 2.87
XR1392 D1011.n323 D1011.n322 2.87
XR1393 D1011.n491 D1011.n488 2.87
XR1394 D1011.n360 D1011.n357 2.87
XR1395 D1011.n363 D1011.n362 2.87
XR1396 D1011.n278 D1011.n276 2.87
XR1397 D1011.n272 D1011.n271 2.87
XR1398 D1011.n175 D1011.n172 2.87
XR1399 D1011.n44 D1011.n41 2.87
XR1400 D1011.n47 D1011.n46 2.87
XR1401 D1011.n335 D1011.n332 2.511
XR1402 D1011.n332 D1011.n331 2.511
XR1403 D1011.n481 D1011.n480 2.511
XR1404 D1011.n412 D1011.n411 2.511
XR1405 D1011.n284 D1011.n281 2.511
XR1406 D1011.n281 D1011.n280 2.511
XR1407 D1011.n165 D1011.n164 2.511
XR1408 D1011.n96 D1011.n95 2.511
XR1409 D1011.n321 D1011.n319 2.152
XR1410 D1011.n315 D1011.n314 2.152
XR1411 D1011.n502 D1011.n499 2.152
XR1412 D1011.n368 D1011.n365 2.152
XR1413 D1011.n371 D1011.n370 2.152
XR1414 D1011.n270 D1011.n268 2.152
XR1415 D1011.n264 D1011.n263 2.152
XR1416 D1011.n186 D1011.n183 2.152
XR1417 D1011.n52 D1011.n49 2.152
XR1418 D1011.n55 D1011.n54 2.152
XR1419 D1011.n343 D1011.n340 1.794
XR1420 D1011.n340 D1011.n339 1.794
XR1421 D1011.n470 D1011.n469 1.794
XR1422 D1011.n423 D1011.n422 1.794
XR1423 D1011.n292 D1011.n289 1.794
XR1424 D1011.n289 D1011.n288 1.794
XR1425 D1011.n154 D1011.n153 1.794
XR1426 D1011.n107 D1011.n106 1.794
XR1427 D1011.n1 D1011.n586 1.706
XR1428 D1011.n1 D1011.n575 1.704
XR1429 D1011.n0 D1011.n36 1.704
XR1430 D1011.n0 D1011.n306 1.704
XR1431 D1011.n0 D1011.n35 7.708
XR1432 D1011.n1 D1011.n574 1.7
XR1433 D1011.n0 D1011.n587 1.7
XR1434 D1011.n573 D1011.n307 1.5
XR1435 D1011.n305 D1011.n39 1.5
XR1436 D1011.n15 D1011.n11 1.467
XR1437 D1011.n518 D1011.n515 1.435
XR1438 D1011.n521 D1011.n520 1.435
XR1439 D1011.n540 D1011.n539 1.435
XR1440 D1011.n537 D1011.n534 1.435
XR1441 D1011.n376 D1011.n373 1.435
XR1442 D1011.n379 D1011.n378 1.435
XR1443 D1011.n202 D1011.n199 1.435
XR1444 D1011.n205 D1011.n204 1.435
XR1445 D1011.n224 D1011.n223 1.435
XR1446 D1011.n221 D1011.n218 1.435
XR1447 D1011.n60 D1011.n57 1.435
XR1448 D1011.n63 D1011.n62 1.435
XR1449 D1011.n26 D1011.n25 1.32
XR1450 D1011.n21 D1011.n20 1.076
XR1451 D1011.n351 D1011.n348 1.076
XR1452 D1011.n348 D1011.n347 1.076
XR1453 D1011.n459 D1011.n458 1.076
XR1454 D1011.n434 D1011.n433 1.076
XR1455 D1011.n300 D1011.n297 1.076
XR1456 D1011.n297 D1011.n296 1.076
XR1457 D1011.n143 D1011.n142 1.076
XR1458 D1011.n118 D1011.n117 1.076
XR1459 D1011.n25 D1011.n8 0.747
XR1460 D1011.n17 D1011.n24 0.717
XR1461 D1011.n526 D1011.n523 0.717
XR1462 D1011.n529 D1011.n528 0.717
XR1463 D1011.n548 D1011.n547 0.717
XR1464 D1011.n545 D1011.n542 0.717
XR1465 D1011.n384 D1011.n381 0.717
XR1466 D1011.n387 D1011.n386 0.717
XR1467 D1011.n210 D1011.n207 0.717
XR1468 D1011.n213 D1011.n212 0.717
XR1469 D1011.n232 D1011.n231 0.717
XR1470 D1011.n229 D1011.n226 0.717
XR1471 D1011.n68 D1011.n65 0.717
XR1472 D1011.n71 D1011.n70 0.717
XR1473 D1011.n24 D1011.n23 0.358
XR1474 D1011.n2 D1011.n583 0.358
XR1475 D1011.n583 D1011.n582 0.358
XR1476 D1011.n313 D1011.n312 0.358
XR1477 D1011.n355 D1011.n313 0.358
XR1478 D1011.n450 D1011.n449 0.358
XR1479 D1011.n444 D1011.n443 0.358
XR1480 D1011.n35 D1011.n34 0.358
XR1481 D1011.n34 D1011.n33 0.358
XR1482 D1011.n262 D1011.n261 0.358
XR1483 D1011.n304 D1011.n262 0.358
XR1484 D1011.n134 D1011.n133 0.358
XR1485 D1011.n128 D1011.n127 0.358
XR1486 D1011.n23 D1011.n22 0.326
XR1487 D1011.n237 D1011.n236 0.19
XR1488 D1011.n236 D1011.n197 0.19
XR1489 D1011.n3 D1011.n4 0.19
XR1490 D1011.n553 D1011.n552 0.19
XR1491 D1011.n552 D1011.n513 0.19
XR1492 D1011.n5 D1011.n6 0.19
XR1493 D1011.n255 D1011.n254 0.144
XR1494 D1011.n252 D1011.n251 0.144
XR1495 D1011.n249 D1011.n248 0.144
XR1496 D1011.n246 D1011.n245 0.144
XR1497 D1011.n243 D1011.n242 0.144
XR1498 D1011.n240 D1011.n239 0.144
XR1499 D1011.n195 D1011.n194 0.144
XR1500 D1011.n192 D1011.n191 0.144
XR1501 D1011.n188 D1011.n181 0.144
XR1502 D1011.n177 D1011.n170 0.144
XR1503 D1011.n166 D1011.n159 0.144
XR1504 D1011.n155 D1011.n148 0.144
XR1505 D1011.n144 D1011.n137 0.144
XR1506 D1011.n121 D1011.n119 0.144
XR1507 D1011.n110 D1011.n108 0.144
XR1508 D1011.n99 D1011.n97 0.144
XR1509 D1011.n88 D1011.n86 0.144
XR1510 D1011.n84 D1011.n83 0.144
XR1511 D1011.n81 D1011.n80 0.144
XR1512 D1011.n78 D1011.n77 0.144
XR1513 D1011.n571 D1011.n570 0.144
XR1514 D1011.n568 D1011.n567 0.144
XR1515 D1011.n565 D1011.n564 0.144
XR1516 D1011.n562 D1011.n561 0.144
XR1517 D1011.n559 D1011.n558 0.144
XR1518 D1011.n556 D1011.n555 0.144
XR1519 D1011.n511 D1011.n510 0.144
XR1520 D1011.n508 D1011.n507 0.144
XR1521 D1011.n504 D1011.n497 0.144
XR1522 D1011.n493 D1011.n486 0.144
XR1523 D1011.n482 D1011.n475 0.144
XR1524 D1011.n471 D1011.n464 0.144
XR1525 D1011.n460 D1011.n453 0.144
XR1526 D1011.n437 D1011.n435 0.144
XR1527 D1011.n426 D1011.n424 0.144
XR1528 D1011.n415 D1011.n413 0.144
XR1529 D1011.n404 D1011.n402 0.144
XR1530 D1011.n400 D1011.n399 0.144
XR1531 D1011.n397 D1011.n396 0.144
XR1532 D1011.n394 D1011.n393 0.144
XR1533 D1011.n8 D1011.n7 0.113
XR1534 D1011.n39 D1011.n256 0.148
XR1535 D1011.n307 D1011.n572 0.148
XR1536 D1011 D1011.n26 0.059
XR1537 D1011.n239 D1011.n238 0.04
XR1538 D1011.n196 D1011.n195 0.04
XR1539 D1011.n77 D1011.n76 0.04
XR1540 D1011.n555 D1011.n554 0.04
XR1541 D1011.n512 D1011.n511 0.04
XR1542 D1011.n393 D1011.n392 0.04
XR1543 D1011.n256 D1011.n255 0.038
XR1544 D1011.n148 D1011.n146 0.038
XR1545 D1011.n112 D1011.n110 0.038
XR1546 D1011.n572 D1011.n571 0.038
XR1547 D1011.n464 D1011.n462 0.038
XR1548 D1011.n428 D1011.n426 0.038
XR1549 D1011.n242 D1011.n241 0.035
XR1550 D1011.n193 D1011.n192 0.035
XR1551 D1011.n80 D1011.n79 0.035
XR1552 D1011.n558 D1011.n557 0.035
XR1553 D1011.n509 D1011.n508 0.035
XR1554 D1011.n396 D1011.n395 0.035
XR1555 D1011.n253 D1011.n252 0.032
XR1556 D1011.n159 D1011.n157 0.032
XR1557 D1011.n101 D1011.n99 0.032
XR1558 D1011.n569 D1011.n568 0.032
XR1559 D1011.n475 D1011.n473 0.032
XR1560 D1011.n417 D1011.n415 0.032
XR1561 D1011.n586 D1011.n584 0.031
XR1562 D1011.n306 D1011.n37 0.031
XR1563 D1011.n245 D1011.n244 0.029
XR1564 D1011.n190 D1011.n188 0.029
XR1565 D1011.n83 D1011.n82 0.029
XR1566 D1011.n561 D1011.n560 0.029
XR1567 D1011.n506 D1011.n504 0.029
XR1568 D1011.n399 D1011.n398 0.029
XR1569 D1011.n250 D1011.n249 0.027
XR1570 D1011.n170 D1011.n168 0.027
XR1571 D1011.n90 D1011.n88 0.027
XR1572 D1011.n566 D1011.n565 0.027
XR1573 D1011.n486 D1011.n484 0.027
XR1574 D1011.n406 D1011.n404 0.027
XR1575 D1011.n248 D1011.n247 0.024
XR1576 D1011.n179 D1011.n177 0.024
XR1577 D1011.n86 D1011.n85 0.024
XR1578 D1011.n564 D1011.n563 0.024
XR1579 D1011.n495 D1011.n493 0.024
XR1580 D1011.n402 D1011.n401 0.024
XR1581 D1011.n247 D1011.n246 0.021
XR1582 D1011.n181 D1011.n179 0.021
XR1583 D1011.n85 D1011.n84 0.021
XR1584 D1011.n563 D1011.n562 0.021
XR1585 D1011.n497 D1011.n495 0.021
XR1586 D1011.n401 D1011.n400 0.021
XR1587 D1011.n251 D1011.n250 0.019
XR1588 D1011.n168 D1011.n166 0.019
XR1589 D1011.n97 D1011.n90 0.019
XR1590 D1011.n567 D1011.n566 0.019
XR1591 D1011.n484 D1011.n482 0.019
XR1592 D1011.n413 D1011.n406 0.019
XR1593 D1011.n16 D1011.n10 0.019
XR1594 D1011.n18 D1011.n16 0.017
XR1595 D1011.n244 D1011.n243 0.016
XR1596 D1011.n191 D1011.n190 0.016
XR1597 D1011.n82 D1011.n81 0.016
XR1598 D1011.n560 D1011.n559 0.016
XR1599 D1011.n507 D1011.n506 0.016
XR1600 D1011.n398 D1011.n397 0.016
XR1601 D1011.n574 D1011.n573 0.014
XR1602 D1011.n254 D1011.n253 0.013
XR1603 D1011.n157 D1011.n155 0.013
XR1604 D1011.n108 D1011.n101 0.013
XR1605 D1011.n570 D1011.n569 0.013
XR1606 D1011.n473 D1011.n471 0.013
XR1607 D1011.n424 D1011.n417 0.013
XR1608 D1011.n7 D1011.n9 0.012
XR1609 D1011.n241 D1011.n240 0.01
XR1610 D1011.n194 D1011.n193 0.01
XR1611 D1011.n79 D1011.n78 0.01
XR1612 D1011.n557 D1011.n556 0.01
XR1613 D1011.n510 D1011.n509 0.01
XR1614 D1011.n395 D1011.n394 0.01
XR1615 D1011.n584 D1011.n585 0.009
XR1616 D1011.n37 D1011.n38 0.009
XR1617 D1011.n146 D1011.n144 0.008
XR1618 D1011.n119 D1011.n112 0.008
XR1619 D1011.n462 D1011.n460 0.008
XR1620 D1011.n435 D1011.n428 0.008
XR1621 D1011.n306 D1011.n305 0.007
XR1622 D1011.n238 D1011.n237 0.005
XR1623 D1011.n197 D1011.n196 0.005
XR1624 D1011.n76 D1011.n75 0.005
XR1625 D1011.n554 D1011.n553 0.005
XR1626 D1011.n513 D1011.n512 0.005
XR1627 D1011.n392 D1011.n391 0.005
XR1628 D1011.n1 D1011.n2 7.71
XR1629 D1011.n0 D1011.n1 0.144
XR1630 D1011 D1011.n0 0.111
XR1631 D1011.n6 D1011.n437 0.045
XR1632 D1011.n453 D1011.n5 0.045
XR1633 D1011.n4 D1011.n121 0.045
XR1634 D1011.n137 D1011.n3 0.045
XR1635 D2.n1 D2.n6 10.626
XR1636 D2.n0 D2.n31 10.626
XR1637 D2.n24 D2.n23 9.733
XR1638 D2.n42 D2.n41 9.733
XR1639 D2.n20 D2.n19 6.189
XR1640 D2.n36 D2.n35 6.189
XR1641 D2.n9 D2.n7 5.741
XR1642 D2.n22 D2.n21 5.741
XR1643 D2.n37 D2.n34 5.741
XR1644 D2.n46 D2.n45 5.741
XR1645 D2.n6 D2.t0 5.539
XR1646 D2.n6 D2.t2 5.539
XR1647 D2.n31 D2.t3 5.539
XR1648 D2.n31 D2.t1 5.539
XR1649 D2.n18 D2.n22 4.5
XR1650 D2.n1 D2.n9 4.5
XR1651 D2.n0 D2.n37 4.5
XR1652 D2.n40 D2.n46 4.5
XR1653 D2.n30 D2.t4 3.35
XR1654 D2.n15 D2.n3 1.704
XR1655 D2.n28 D2.n27 1.704
XR1656 D2.n14 D2.n13 1.704
XR1657 D2.n52 D2.n30 1.704
XR1658 D2.n49 D2.n48 1.704
XR1659 D2.n15 D2.n2 1.701
XR1660 D2.n51 D2.n50 1.701
XR1661 D2.n26 D2.n18 1.5
XR1662 D2.n12 D2.n1 1.5
XR1663 D2.n47 D2.n40 1.5
XR1664 D2.n9 D2.n8 0.358
XR1665 D2.n22 D2.n20 0.358
XR1666 D2.n37 D2.n36 0.358
XR1667 D2.n46 D2.n44 0.358
XR1668 D2 D2.n29 0.131
XR1669 D2 D2.n53 0.131
XR1670 D2.n12 D2.n4 0.034
XR1671 D2.n1 D2.n10 0.033
XR1672 D2.n0 D2.n32 0.033
XR1673 D2.n27 D2.n16 0.032
XR1674 D2.n48 D2.n38 0.032
XR1675 D2.n40 D2.n43 0.025
XR1676 D2.n18 D2.n25 0.025
XR1677 D2.n16 D2.n17 0.007
XR1678 D2.n38 D2.n39 0.007
XR1679 D2.n27 D2.n26 0.006
XR1680 D2.n48 D2.n47 0.006
XR1681 D2.n29 D2.n28 0.004
XR1682 D2.n52 D2.n51 0.004
XR1683 D2.n28 D2.n15 0.004
XR1684 D2.n15 D2.n14 0.004
XR1685 D2.n53 D2.n52 0.004
XR1686 D2.n51 D2.n49 0.004
XR1687 D2.n32 D2.n33 0.003
XR1688 D2.n43 D2.n42 0.003
XR1689 D2.n10 D2.n11 0.003
XR1690 D2.n25 D2.n24 0.003
XR1691 D2.n13 D2.n12 0.003
XR1692 D2.n4 D2.n5 0.003
XR1693 D2.n30 D2.n0 1.503
XC0 G1011 D5 3.59fF
XC1 VDD G4 8.61fF
XC2 a_2113_n8873# a_1053_n8873# 0.19fF
XC3 a_523_n9665# a_1053_n8873# 0.06fF
XC4 D1011 VDD 9.50fF
XC5 a_3173_n8873# G4 0.06fF
XC6 G1011 G4 0.52fF
XC7 a_2113_n8873# a_2643_n9665# 0.06fF
XC8 D1011 G1011 1.18fF
XC9 VDD D9 2.15fF
XC10 D5 G4 1.32fF
XC11 D2 a_2643_n9665# 0.19fF
XC12 D2 Vref 1.22fF
XC13 VDD D6 0.17fF
XC14 G1011 D9 1.86fF
XC15 Vref VDD 4.10fF
XC16 D1011 G4 0.93fF
XC17 a_n7_n8873# a_1053_n8873# 0.19fF
XC18 a_2643_n9665# a_3173_n8873# 0.06fF
XC19 D5 D9 13.43fF
XC20 G1011 D6 2.55fF
XC21 Vref G1011 3.12fF
XC22 VBJTS a_523_n9665# 0.19fF
XC23 VBJTS D2 0.25fF
XC24 D5 D6 13.15fF
XC25 G4 D9 1.16fF
XC26 Vref a_n7_n8873# 0.19fF
XC27 Vref D5 1.25fF
XC28 a_2113_n8873# D2 0.06fF
XC29 a_2643_n9665# G4 0.19fF
XC30 G4 D6 0.45fF
XC31 Vref G4 0.10fF
XC32 D2 VDD 5.09fF
XC33 a_2113_n8873# a_3173_n8873# 0.19fF
XC34 D9 D6 7.65fF
XC35 D2 G1011 1.35fF
XC36 VBJTS G4 1.92fF
XC37 a_n7_n8873# a_523_n9665# 0.06fF
XC38 VDD G1011 33.26fF
XC39 VDD D5 2.20fF
XC40 D2 G4 1.01fF
XC41 VBJTS a_1053_n8873# 0.06fF
XC42 D1011 GND 4.56fF
XC43 a_3173_n8873# GND 2.22fF
XC44 a_2643_n9665# GND 1.51fF
XC45 D2 GND 1.66fF
XC46 a_2113_n8873# GND 1.86fF
XC47 VBJTS GND 18.00fF
XC48 a_1053_n8873# GND 1.86fF
XC49 a_523_n9665# GND 1.51fF
XC50 a_n7_n8873# GND 1.86fF
XC51 Vref GND 8.86fF
XC52 D6 GND 13.83fF
XC53 D9 GND 12.96fF
XC54 G4 GND 9.61fF
XC55 D5 GND 7.29fF
XC56 G1011 GND 52.29fF
XC57 VDD GND 121.12fF
XC58 D2.n0 GND 0.11fF
XC59 D2.n1 GND 0.11fF
XC60 D2.n2 GND 0.01fF
XC61 D2.n3 GND 0.01fF
XC62 D2.t0 GND 0.06fF
XC63 D2.t2 GND 0.06fF
XC64 D2.n6 GND 0.22fF
XC65 D2.n14 GND 0.02fF
XC66 D2.n15 GND 0.02fF
XC67 D2.n18 GND 0.02fF
XC68 D2.n23 GND 0.01fF
XC69 D2.n24 GND 0.09fF
XC70 D2.n29 GND 0.16fF
XC71 D2.t4 GND 2.71fF
XC72 D2.n30 GND 0.40fF
XC73 D2.t3 GND 0.06fF
XC74 D2.t1 GND 0.06fF
XC75 D2.n31 GND 0.22fF
XC76 D2.n40 GND 0.02fF
XC77 D2.n41 GND 0.01fF
XC78 D2.n42 GND 0.09fF
XC79 D2.n49 GND 0.02fF
XC80 D2.n50 GND 0.01fF
XC81 D2.n51 GND 0.02fF
XC82 D2.n53 GND 0.16fF
XC83 D1011.n0 GND 0.28fF
XC84 D1011.n1 GND 0.20fF
XC85 D1011.n2 GND 0.02fF
XC86 D1011.t0 GND 0.12fF
XC87 D1011.n7 GND 0.01fF
XC88 D1011.n8 GND 0.02fF
XC89 D1011.t3 GND 2.06fF
XC90 D1011.n10 GND 0.81fF
XC91 D1011.n11 GND 0.02fF
XC92 D1011.t4 GND 2.01fF
XC93 D1011.n12 GND 0.70fF
XC94 D1011.n13 GND 0.02fF
XC95 D1011.n18 GND 0.03fF
XC96 D1011.n19 GND 0.02fF
XC97 D1011.n25 GND 0.19fF
XC98 D1011.n26 GND 3.35fF
XC99 D1011.n27 GND 0.03fF
XC100 D1011.n35 GND 0.02fF
XC101 D1011.n36 GND 0.01fF
XC102 D1011.n39 GND 0.02fF
XC103 D1011.n74 GND 0.06fF
XC104 D1011.n75 GND 0.91fF
XC105 D1011.n214 GND 0.01fF
XC106 D1011.n233 GND 0.01fF
XC107 D1011.n236 GND 0.01fF
XC108 D1011.n307 GND 0.02fF
XC109 D1011.n390 GND 0.06fF
XC110 D1011.n391 GND 0.91fF
XC111 D1011.n530 GND 0.01fF
XC112 D1011.n549 GND 0.01fF
XC113 D1011.n552 GND 0.01fF
XC114 D1011.n575 GND 0.01fF
XC115 D1011.n576 GND 0.03fF
XC116 Vref.n0 GND 2.04fF
XC117 Vref.n1 GND 0.17fF
XC118 Vref.n4 GND 0.22fF
XC119 Vref.t4 GND 2.20fF
XC120 Vref.t1 GND 0.07fF
XC121 Vref.n6 GND 0.01fF
XC122 Vref.t0 GND 0.07fF
XC123 Vref.n7 GND 0.29fF
XC124 Vref.n8 GND 0.22fF
XC125 Vref.n14 GND 0.02fF
XC126 Vref.n18 GND 0.03fF
XC127 Vref.n19 GND 0.01fF
XC128 Vref.t3 GND 0.07fF
XC129 Vref.t2 GND 0.07fF
XC130 Vref.n21 GND 0.01fF
XC131 Vref.n22 GND 0.29fF
XC132 Vref.n26 GND 0.02fF
XC133 Vref.n27 GND 0.01fF
XC134 Vref.n28 GND 0.02fF
XC135 Vref.n29 GND 0.03fF
XC136 Vref.n35 GND 0.02fF
XC137 Vref.n36 GND 6.62fF
XC138 G3.n0 GND 0.46fF
XC139 G3.n1 GND 0.29fF
XC140 G3.t0 GND 1.53fF
XC141 G3.t3 GND 0.25fF
XC142 G3.t5 GND 0.26fF
XC143 G3.t4 GND 0.26fF
XC144 G3.t2 GND 0.26fF
XC145 G3.t1 GND 0.26fF
XC146 G3.t6 GND 0.26fF
XC147 D9.n0 GND 0.11fF
XC148 D9.n1 GND 0.30fF
XC149 D9.n2 GND 1.03fF
XC150 D9.n3 GND 0.26fF
XC151 D9.n4 GND 1.04fF
XC152 D9.n5 GND 0.04fF
XC153 D9.n6 GND 0.04fF
XC154 D9.n7 GND 0.05fF
XC155 D9.n9 GND 0.05fF
XC156 D9.n11 GND 0.02fF
XC157 D9.n12 GND 0.05fF
XC158 D9.n14 GND 0.02fF
XC159 D9.n15 GND 0.05fF
XC160 D9.n17 GND 0.02fF
XC161 D9.n18 GND 0.02fF
XC162 D9.n19 GND 1.70fF
XC163 D9.n21 GND 0.13fF
XC164 D9.n25 GND 0.52fF
XC165 D9.n27 GND 0.01fF
XC166 D9.n30 GND 0.03fF
XC167 D9.n31 GND 0.03fF
XC168 D9.n32 GND 0.52fF
XC169 D9.n34 GND 0.01fF
XC170 D9.n38 GND 0.01fF
XC171 D9.t5 GND 0.03fF
XC172 D9.n42 GND 0.03fF
XC173 D9.n43 GND 0.02fF
XC174 D9.n44 GND 0.16fF
XC175 D9.n45 GND 2.01fF
XC176 D9.n47 GND 0.01fF
XC177 D9.n48 GND 0.02fF
XC178 D9.n50 GND 0.02fF
XC179 D9.n52 GND 0.02fF
XC180 D9.n59 GND 0.02fF
XC181 D9.n62 GND 0.02fF
XC182 D9.n66 GND 1.70fF
XC183 D9.n68 GND 0.13fF
XC184 D9.n72 GND 0.03fF
XC185 D9.n73 GND 0.03fF
XC186 D9.n74 GND 0.24fF
XC187 D9.n76 GND 0.01fF
XC188 D9.n81 GND 0.01fF
XC189 D9.t0 GND 0.45fF
XC190 D9.n84 GND 0.04fF
XC191 D9.t1 GND 0.45fF
XC192 D9.n85 GND 2.11fF
XC193 D9.n86 GND 0.04fF
XC194 D9.n87 GND 0.59fF
XC195 D9.n89 GND 0.03fF
XC196 D9.n90 GND 0.03fF
XC197 D9.n92 GND 0.01fF
XC198 D9.n97 GND 0.01fF
XC199 D9.t4 GND 0.45fF
XC200 D9.n100 GND 0.04fF
XC201 D9.t2 GND 0.45fF
XC202 D9.n101 GND 2.11fF
XC203 D9.n102 GND 0.04fF
XC204 D9.n103 GND 0.59fF
XC205 D9.n105 GND 0.24fF
XC206 D9.n106 GND 0.03fF
XC207 D9.n107 GND 0.03fF
XC208 D9.n109 GND 0.01fF
XC209 D9.t3 GND 0.03fF
XC210 D9.n113 GND 0.03fF
XC211 D9.n114 GND 0.02fF
XC212 D9.n115 GND 0.16fF
XC213 D9.n116 GND 2.01fF
XC214 D9.n118 GND 0.01fF
XC215 D9.n119 GND 0.02fF
XC216 D9.n121 GND 0.02fF
XC217 D9.n123 GND 0.02fF
XC218 D9.n130 GND 0.02fF
XC219 D9.n133 GND 0.02fF
XC220 D9.n137 GND 1.90fF
XC221 D9.n138 GND 0.68fF
XC222 D9.n139 GND 0.03fF
XC223 D9.n140 GND 0.69fF
XC224 D9.n141 GND 0.88fF
XC225 D9.n142 GND 0.06fF
XC226 D9.n143 GND 0.61fF
XC227 D9.n144 GND 0.68fF
XC228 D9.n145 GND 0.03fF
XC229 D9.n146 GND 0.46fF
XC230 D9.n147 GND 0.17fF
XC231 D9.t10 GND 0.08fF
XC232 D9.n148 GND 0.17fF
XC233 D9.t8 GND 0.08fF
XC234 D9.n149 GND 0.46fF
XC235 D9.n150 GND 0.06fF
XC236 D9.t9 GND 0.01fF
XC237 D9.t13 GND 0.01fF
XC238 D9.n151 GND 0.17fF
XC239 D9.t6 GND 0.08fF
XC240 D9.n152 GND 0.39fF
XC241 D9.t17 GND 0.08fF
XC242 D9.t16 GND 0.08fF
XC243 D9.n153 GND 0.17fF
XC244 D9.t12 GND 0.08fF
XC245 D9.n154 GND 0.39fF
XC246 D9.t14 GND 0.08fF
XC247 D9.t15 GND 0.08fF
XC248 D9.n155 GND 0.06fF
XC249 D9.t7 GND 0.01fF
XC250 D9.t11 GND 0.01fF
XC251 D5.n0 GND 2.74fF
XC252 D5.n1 GND 0.45fF
XC253 D5.n2 GND 0.47fF
XC254 D5.n3 GND 2.96fF
XC255 D5.n4 GND 1.00fF
XC256 D5.n5 GND 0.06fF
XC257 D5.n6 GND 0.78fF
XC258 D5.n7 GND 0.45fF
XC259 D5.t2 GND 0.03fF
XC260 D5.t0 GND 0.03fF
XC261 D5.n8 GND 0.14fF
XC262 D5.n9 GND 0.06fF
XC263 D5.t1 GND 0.03fF
XC264 D5.t3 GND 0.03fF
XC265 D5.n10 GND 0.13fF
XC266 D5.n11 GND 0.42fF
XC267 D5.n12 GND 0.05fF
XC268 D5.t8 GND 0.39fF
XC269 D5.n13 GND 0.01fF
XC270 D5.t9 GND 0.39fF
XC271 D5.n14 GND 2.51fF
XC272 D5.t13 GND 0.39fF
XC273 D5.n15 GND 0.01fF
XC274 D5.t15 GND 0.39fF
XC275 D5.n16 GND 2.51fF
XC276 D5.t5 GND 0.39fF
XC277 D5.n17 GND 0.01fF
XC278 D5.t6 GND 0.39fF
XC279 D5.n18 GND 2.51fF
XC280 D5.n19 GND 0.26fF
XC281 D5.t7 GND 0.39fF
XC282 D5.n20 GND 0.02fF
XC283 D5.t11 GND 0.39fF
XC284 D5.n21 GND 2.17fF
XC285 D5.n22 GND 0.01fF
XC286 D5.n23 GND 0.59fF
XC287 D5.t12 GND 0.39fF
XC288 D5.n24 GND 0.01fF
XC289 D5.t14 GND 0.39fF
XC290 D5.n25 GND 2.39fF
XC291 D5.n26 GND 0.09fF
XC292 D5.n27 GND 0.12fF
XC293 D5.n29 GND 0.02fF
XC294 D5.n30 GND 0.44fF
XC295 D5.n32 GND 0.02fF
XC296 D5.n33 GND 0.65fF
XC297 D5.t10 GND 0.39fF
XC298 D5.n34 GND 0.01fF
XC299 D5.t4 GND 0.39fF
XC300 D5.n35 GND 2.39fF
XC301 D6.n0 GND 0.73fF
XC302 D6.n1 GND 3.05fF
XC303 D6.n2 GND 0.92fF
XC304 D6.n3 GND 0.68fF
XC305 D6.n4 GND 2.75fF
XC306 D6.n5 GND 0.41fF
XC307 D6.t12 GND 0.10fF
XC308 D6.t19 GND 0.10fF
XC309 D6.n6 GND 0.28fF
XC310 D6.t15 GND 0.10fF
XC311 D6.n7 GND 0.15fF
XC312 D6.t11 GND 0.10fF
XC313 D6.n8 GND 0.14fF
XC314 D6.t18 GND 0.04fF
XC315 D6.n9 GND 1.59fF
XC316 D6.t1 GND 0.57fF
XC317 D6.n10 GND 0.02fF
XC318 D6.t2 GND 0.57fF
XC319 D6.n11 GND 3.26fF
XC320 D6.n15 GND 0.02fF
XC321 D6.n16 GND 0.04fF
XC322 D6.t4 GND 0.57fF
XC323 D6.n17 GND 0.02fF
XC324 D6.t3 GND 0.57fF
XC325 D6.n18 GND 3.26fF
XC326 D6.n19 GND 1.14fF
XC327 D6.n23 GND 0.02fF
XC328 D6.n24 GND 0.04fF
XC329 D6.t5 GND 0.57fF
XC330 D6.n25 GND 0.02fF
XC331 D6.t0 GND 0.57fF
XC332 D6.n26 GND 3.26fF
XC333 D6.n27 GND 0.91fF
XC334 D6.n28 GND 0.02fF
XC335 D6.n32 GND 0.02fF
XC336 D6.t14 GND 0.10fF
XC337 D6.t13 GND 0.10fF
XC338 D6.t10 GND 0.10fF
XC339 D6.t17 GND 0.10fF
XC340 D6.n33 GND 0.28fF
XC341 D6.n34 GND 0.15fF
XC342 D6.n35 GND 0.14fF
XC343 D6.t16 GND 0.04fF
XC344 D6.n36 GND 1.98fF
XC345 D6.t9 GND 0.02fF
XC346 D6.t8 GND 0.02fF
XC347 D6.n37 GND 0.08fF
XC348 D6.n38 GND 1.39fF
XC349 D6.n39 GND 0.08fF
XC350 D6.n40 GND 0.27fF
XC351 D6.n41 GND 2.19fF
XC352 D6.n42 GND 0.08fF
XC353 D6.t6 GND 0.02fF
XC354 D6.t7 GND 0.02fF
XC355 G1011.n0 GND 2.57fF
XC356 G1011.n1 GND 0.07fF
XC357 G1011.n2 GND 0.01fF
XC358 G1011.n3 GND 0.90fF
XC359 G1011.n4 GND 0.23fF
XC360 G1011.n5 GND 1.05fF
XC361 G1011.n6 GND 0.22fF
XC362 G1011.n7 GND 0.22fF
XC363 G1011.n8 GND 0.27fF
XC364 G1011.n9 GND 0.22fF
XC365 G1011.n10 GND 0.22fF
XC366 G1011.n11 GND 0.22fF
XC367 G1011.n12 GND 0.22fF
XC368 G1011.n13 GND 0.22fF
XC369 G1011.n14 GND 0.22fF
XC370 G1011.n15 GND 0.23fF
XC371 G1011.n16 GND 0.22fF
XC372 G1011.n17 GND 0.22fF
XC373 G1011.n18 GND 0.64fF
XC374 G1011.n19 GND 0.23fF
XC375 G1011.n20 GND 0.22fF
XC376 G1011.n21 GND 0.22fF
XC377 G1011.n22 GND 0.22fF
XC378 G1011.n23 GND 0.22fF
XC379 G1011.n24 GND 0.22fF
XC380 G1011.n25 GND 0.22fF
XC381 G1011.n26 GND 0.22fF
XC382 G1011.n27 GND 0.22fF
XC383 G1011.n28 GND 4.27fF
XC384 G1011.n29 GND 0.19fF
XC385 G1011.n30 GND 0.19fF
XC386 G1011.n31 GND 0.19fF
XC387 G1011.n32 GND 0.19fF
XC388 G1011.n33 GND 0.19fF
XC389 G1011.n34 GND 0.19fF
XC390 G1011.n35 GND 0.19fF
XC391 G1011.n36 GND 0.19fF
XC392 G1011.n37 GND 0.19fF
XC393 G1011.n38 GND 0.60fF
XC394 G1011.n39 GND 0.19fF
XC395 G1011.n40 GND 0.19fF
XC396 G1011.n41 GND 0.19fF
XC397 G1011.n42 GND 0.19fF
XC398 G1011.n43 GND 0.19fF
XC399 G1011.n44 GND 0.19fF
XC400 G1011.n45 GND 0.19fF
XC401 G1011.n46 GND 0.19fF
XC402 G1011.n47 GND 0.19fF
XC403 G1011.n48 GND 0.19fF
XC404 G1011.n49 GND 0.04fF
XC405 G1011.n50 GND 0.01fF
XC406 G1011.n51 GND 0.31fF
XC407 G1011.n52 GND 0.02fF
XC408 G1011.n53 GND 0.02fF
XC409 G1011.n54 GND 0.02fF
XC410 G1011.n55 GND 0.02fF
XC411 G1011.n56 GND 0.02fF
XC412 G1011.n57 GND 0.02fF
XC413 G1011.n58 GND 0.02fF
XC414 G1011.n59 GND 0.02fF
XC415 G1011.n60 GND 0.02fF
XC416 G1011.n61 GND 0.02fF
XC417 G1011.n62 GND 0.02fF
XC418 G1011.n63 GND 0.02fF
XC419 G1011.n64 GND 0.02fF
XC420 G1011.n65 GND 0.02fF
XC421 G1011.n66 GND 0.02fF
XC422 G1011.n67 GND 0.02fF
XC423 G1011.n68 GND 0.02fF
XC424 G1011.n69 GND 0.02fF
XC425 G1011.n70 GND 0.02fF
XC426 G1011.n71 GND 0.02fF
XC427 G1011.n72 GND 0.02fF
XC428 G1011.n73 GND 0.02fF
XC429 G1011.n74 GND 0.02fF
XC430 G1011.n75 GND 0.02fF
XC431 G1011.n76 GND 0.02fF
XC432 G1011.n77 GND 0.02fF
XC433 G1011.n78 GND 0.02fF
XC434 G1011.n79 GND 0.02fF
XC435 G1011.n80 GND 0.02fF
XC436 G1011.n81 GND 0.02fF
XC437 G1011.n82 GND 0.02fF
XC438 G1011.n83 GND 0.02fF
XC439 G1011.n84 GND 0.02fF
XC440 G1011.n85 GND 0.02fF
XC441 G1011.n86 GND 0.02fF
XC442 G1011.n87 GND 0.02fF
XC443 G1011.n88 GND 0.02fF
XC444 G1011.n89 GND 0.02fF
XC445 G1011.n90 GND 0.02fF
XC446 G1011.n91 GND 0.02fF
XC447 G1011.n92 GND 0.02fF
XC448 G1011.n93 GND 0.02fF
XC449 G1011.n94 GND 0.02fF
XC450 G1011.n95 GND 0.02fF
XC451 G1011.n96 GND 0.02fF
XC452 G1011.n97 GND 0.03fF
XC453 G1011.t101 GND 3.51fF
XC454 G1011.n98 GND 1.93fF
XC455 G1011.n99 GND 0.04fF
XC456 G1011.n100 GND 0.04fF
XC457 G1011.n101 GND 1.93fF
XC458 G1011.n102 GND 0.01fF
XC459 G1011.n105 GND 0.02fF
XC460 G1011.n112 GND 0.02fF
XC461 G1011.n113 GND 0.02fF
XC462 G1011.n120 GND 0.02fF
XC463 G1011.n121 GND 0.03fF
XC464 G1011.n122 GND 0.01fF
XC465 G1011.t107 GND 7.53fF
XC466 G1011.n123 GND 0.75fF
XC467 G1011.n124 GND 0.33fF
XC468 G1011.n125 GND 0.03fF
XC469 G1011.n127 GND 0.02fF
XC470 G1011.n132 GND 0.02fF
XC471 G1011.n135 GND 0.02fF
XC472 G1011.n140 GND 0.02fF
XC473 G1011.n143 GND 0.02fF
XC474 G1011.n148 GND 0.02fF
XC475 G1011.n151 GND 0.02fF
XC476 G1011.n156 GND 0.02fF
XC477 G1011.n159 GND 0.02fF
XC478 G1011.n163 GND 1.79fF
XC479 G1011.n164 GND 0.17fF
XC480 G1011.n168 GND 0.01fF
XC481 G1011.n169 GND 0.51fF
XC482 G1011.n170 GND 0.56fF
XC483 G1011.n171 GND 0.09fF
XC484 G1011.n174 GND 0.05fF
XC485 G1011.n175 GND 0.02fF
XC486 G1011.n178 GND 0.02fF
XC487 G1011.n181 GND 0.05fF
XC488 G1011.n182 GND 1.65fF
XC489 G1011.t105 GND 3.26fF
XC490 G1011.n183 GND 1.65fF
XC491 G1011.n184 GND 0.05fF
XC492 G1011.n188 GND 0.03fF
XC493 G1011.n189 GND 0.05fF
XC494 G1011.n192 GND 0.02fF
XC495 G1011.n195 GND 0.02fF
XC496 G1011.n196 GND 0.02fF
XC497 G1011.n197 GND 0.02fF
XC498 G1011.n198 GND 0.12fF
XC499 G1011.n199 GND 0.02fF
XC500 G1011.t109 GND 0.63fF
XC501 G1011.t104 GND 0.63fF
XC502 G1011.n200 GND 0.54fF
XC503 G1011.t106 GND 0.63fF
XC504 G1011.n201 GND 0.28fF
XC505 G1011.t110 GND 0.58fF
XC506 G1011.n204 GND 0.01fF
XC507 G1011.n205 GND 0.01fF
XC508 G1011.t100 GND 0.63fF
XC509 G1011.t102 GND 0.63fF
XC510 G1011.t103 GND 0.63fF
XC511 G1011.t108 GND 0.63fF
XC512 G1011.n206 GND 0.54fF
XC513 G1011.n207 GND 0.27fF
XC514 G1011.n208 GND 0.32fF
XC515 G1011.n209 GND 3.43fF
XC516 G1011.n210 GND 3.48fF
XC517 G1011.t68 GND 0.13fF
XC518 G1011.t78 GND 0.13fF
XC519 G1011.t14 GND 0.13fF
XC520 G1011.t15 GND 0.02fF
XC521 G1011.t41 GND 0.02fF
XC522 G1011.n214 GND 0.06fF
XC523 G1011.n215 GND 0.01fF
XC524 G1011.n216 GND 0.02fF
XC525 G1011.t40 GND 0.13fF
XC526 G1011.t82 GND 0.13fF
XC527 G1011.t22 GND 0.13fF
XC528 G1011.n217 GND 0.10fF
XC529 G1011.n218 GND 0.05fF
XC530 G1011.n219 GND 0.10fF
XC531 G1011.n220 GND 0.10fF
XC532 G1011.n221 GND 0.05fF
XC533 G1011.n222 GND 0.10fF
XC534 G1011.n223 GND 0.10fF
XC535 G1011.n224 GND 0.14fF
XC536 G1011.n225 GND 0.01fF
XC537 G1011.n226 GND 0.02fF
XC538 G1011.t69 GND 0.02fF
XC539 G1011.t79 GND 0.02fF
XC540 G1011.n232 GND 0.06fF
XC541 G1011.n233 GND 0.01fF
XC542 G1011.n234 GND 0.08fF
XC543 G1011.t30 GND 0.13fF
XC544 G1011.n235 GND 0.10fF
XC545 G1011.t86 GND 0.13fF
XC546 G1011.n236 GND 0.14fF
XC547 G1011.n237 GND 0.01fF
XC548 G1011.n238 GND 0.02fF
XC549 G1011.t31 GND 0.02fF
XC550 G1011.t87 GND 0.02fF
XC551 G1011.n244 GND 0.06fF
XC552 G1011.n245 GND 0.01fF
XC553 G1011.n246 GND 0.14fF
XC554 G1011.n247 GND 0.11fF
XC555 G1011.n248 GND 0.05fF
XC556 G1011.t90 GND 0.05fF
XC557 G1011.n249 GND 0.05fF
XC558 G1011.n250 GND 0.05fF
XC559 G1011.n251 GND 0.30fF
XC560 G1011.n252 GND 0.05fF
XC561 G1011.n253 GND 0.19fF
XC562 G1011.n254 GND 0.05fF
XC563 G1011.n255 GND 0.05fF
XC564 G1011.n256 GND 0.30fF
XC565 G1011.n257 GND 0.05fF
XC566 G1011.n258 GND 1.01fF
XC567 G1011.n259 GND 0.05fF
XC568 G1011.n260 GND 0.05fF
XC569 G1011.n261 GND 0.30fF
XC570 G1011.n262 GND 0.05fF
XC571 G1011.n263 GND 0.19fF
XC572 G1011.n264 GND 0.05fF
XC573 G1011.n265 GND 0.05fF
XC574 G1011.n266 GND 0.30fF
XC575 G1011.n267 GND 0.05fF
XC576 G1011.n268 GND 0.19fF
XC577 G1011.n269 GND 0.05fF
XC578 G1011.t91 GND 0.05fF
XC579 G1011.n270 GND 0.32fF
XC580 G1011.n271 GND 0.05fF
XC581 G1011.n272 GND 4.19fF
XC582 G1011.n273 GND 0.05fF
XC583 G1011.n274 GND 0.19fF
XC584 G1011.n275 GND 0.05fF
XC585 G1011.t70 GND 0.13fF
XC586 G1011.n276 GND 0.10fF
XC587 G1011.t34 GND 0.13fF
XC588 G1011.n277 GND 0.10fF
XC589 G1011.n278 GND 0.05fF
XC590 G1011.n279 GND 0.01fF
XC591 G1011.n280 GND 0.02fF
XC592 G1011.t71 GND 0.02fF
XC593 G1011.t35 GND 0.02fF
XC594 G1011.n286 GND 0.06fF
XC595 G1011.n287 GND 0.01fF
XC596 G1011.n288 GND 0.14fF
XC597 G1011.n289 GND 0.11fF
XC598 G1011.n290 GND 0.05fF
XC599 G1011.n291 GND 0.05fF
XC600 G1011.t32 GND 0.13fF
XC601 G1011.n292 GND 0.10fF
XC602 G1011.t56 GND 0.13fF
XC603 G1011.n293 GND 0.10fF
XC604 G1011.n294 GND 0.05fF
XC605 G1011.n295 GND 0.01fF
XC606 G1011.n296 GND 0.02fF
XC607 G1011.t33 GND 0.02fF
XC608 G1011.t57 GND 0.02fF
XC609 G1011.n302 GND 0.06fF
XC610 G1011.n303 GND 0.01fF
XC611 G1011.n304 GND 0.14fF
XC612 G1011.n305 GND 0.11fF
XC613 G1011.n306 GND 0.05fF
XC614 G1011.n307 GND 0.05fF
XC615 G1011.t72 GND 0.13fF
XC616 G1011.n308 GND 0.10fF
XC617 G1011.t36 GND 0.13fF
XC618 G1011.n309 GND 0.10fF
XC619 G1011.n310 GND 0.05fF
XC620 G1011.n311 GND 0.01fF
XC621 G1011.n312 GND 0.02fF
XC622 G1011.t73 GND 0.02fF
XC623 G1011.t37 GND 0.02fF
XC624 G1011.n318 GND 0.06fF
XC625 G1011.n319 GND 0.01fF
XC626 G1011.n320 GND 0.14fF
XC627 G1011.n321 GND 0.11fF
XC628 G1011.n322 GND 0.05fF
XC629 G1011.n323 GND 0.05fF
XC630 G1011.t18 GND 0.13fF
XC631 G1011.n324 GND 0.10fF
XC632 G1011.t10 GND 0.13fF
XC633 G1011.n325 GND 0.10fF
XC634 G1011.n326 GND 0.05fF
XC635 G1011.n327 GND 0.01fF
XC636 G1011.n328 GND 0.02fF
XC637 G1011.t19 GND 0.02fF
XC638 G1011.t11 GND 0.02fF
XC639 G1011.n334 GND 0.06fF
XC640 G1011.n335 GND 0.01fF
XC641 G1011.n336 GND 0.14fF
XC642 G1011.n337 GND 0.11fF
XC643 G1011.n338 GND 0.05fF
XC644 G1011.n339 GND 0.05fF
XC645 G1011.t74 GND 0.13fF
XC646 G1011.n340 GND 0.10fF
XC647 G1011.t64 GND 0.13fF
XC648 G1011.n341 GND 0.10fF
XC649 G1011.n342 GND 0.05fF
XC650 G1011.n343 GND 0.01fF
XC651 G1011.n344 GND 0.02fF
XC652 G1011.t75 GND 0.02fF
XC653 G1011.t65 GND 0.02fF
XC654 G1011.n350 GND 0.06fF
XC655 G1011.n351 GND 0.01fF
XC656 G1011.n352 GND 0.14fF
XC657 G1011.n353 GND 0.11fF
XC658 G1011.n354 GND 0.05fF
XC659 G1011.n355 GND 0.05fF
XC660 G1011.t44 GND 0.13fF
XC661 G1011.n356 GND 0.10fF
XC662 G1011.t12 GND 0.13fF
XC663 G1011.n357 GND 0.10fF
XC664 G1011.n358 GND 0.05fF
XC665 G1011.n359 GND 0.01fF
XC666 G1011.n360 GND 0.02fF
XC667 G1011.t45 GND 0.02fF
XC668 G1011.t13 GND 0.02fF
XC669 G1011.n366 GND 0.06fF
XC670 G1011.n367 GND 0.01fF
XC671 G1011.n368 GND 0.14fF
XC672 G1011.n369 GND 0.11fF
XC673 G1011.n370 GND 0.05fF
XC674 G1011.n371 GND 0.05fF
XC675 G1011.t20 GND 0.13fF
XC676 G1011.n372 GND 0.10fF
XC677 G1011.t48 GND 0.13fF
XC678 G1011.n373 GND 0.10fF
XC679 G1011.n374 GND 0.05fF
XC680 G1011.n375 GND 0.01fF
XC681 G1011.n376 GND 0.02fF
XC682 G1011.t21 GND 0.02fF
XC683 G1011.t49 GND 0.02fF
XC684 G1011.n382 GND 0.06fF
XC685 G1011.n383 GND 0.01fF
XC686 G1011.n384 GND 0.14fF
XC687 G1011.n385 GND 0.11fF
XC688 G1011.n386 GND 0.05fF
XC689 G1011.n387 GND 0.05fF
XC690 G1011.t52 GND 0.13fF
XC691 G1011.n388 GND 0.10fF
XC692 G1011.t28 GND 0.13fF
XC693 G1011.n389 GND 0.10fF
XC694 G1011.n390 GND 0.05fF
XC695 G1011.n391 GND 0.01fF
XC696 G1011.n392 GND 0.02fF
XC697 G1011.t53 GND 0.02fF
XC698 G1011.t29 GND 0.02fF
XC699 G1011.n398 GND 0.06fF
XC700 G1011.n399 GND 0.01fF
XC701 G1011.n400 GND 0.14fF
XC702 G1011.n401 GND 0.11fF
XC703 G1011.n402 GND 0.05fF
XC704 G1011.n403 GND 0.05fF
XC705 G1011.t6 GND 0.13fF
XC706 G1011.n404 GND 0.10fF
XC707 G1011.t58 GND 0.13fF
XC708 G1011.n405 GND 0.10fF
XC709 G1011.n406 GND 0.05fF
XC710 G1011.n407 GND 0.01fF
XC711 G1011.n408 GND 0.02fF
XC712 G1011.t7 GND 0.02fF
XC713 G1011.t59 GND 0.02fF
XC714 G1011.n414 GND 0.06fF
XC715 G1011.n415 GND 0.01fF
XC716 G1011.n416 GND 0.14fF
XC717 G1011.n417 GND 0.11fF
XC718 G1011.n418 GND 0.05fF
XC719 G1011.n419 GND 0.05fF
XC720 G1011.t111 GND 0.13fF
XC721 G1011.n420 GND 0.12fF
XC722 G1011.t98 GND 0.13fF
XC723 G1011.n421 GND 0.12fF
XC724 G1011.t76 GND 0.13fF
XC725 G1011.n422 GND 0.10fF
XC726 G1011.t66 GND 0.13fF
XC727 G1011.n423 GND 0.10fF
XC728 G1011.n424 GND 0.05fF
XC729 G1011.n425 GND 0.01fF
XC730 G1011.n426 GND 0.02fF
XC731 G1011.t77 GND 0.02fF
XC732 G1011.t67 GND 0.02fF
XC733 G1011.n432 GND 0.06fF
XC734 G1011.n433 GND 0.01fF
XC735 G1011.n434 GND 0.14fF
XC736 G1011.n435 GND 0.11fF
XC737 G1011.n436 GND 0.05fF
XC738 G1011.n437 GND 0.05fF
XC739 G1011.t4 GND 0.13fF
XC740 G1011.n438 GND 0.10fF
XC741 G1011.t38 GND 0.13fF
XC742 G1011.t99 GND 0.13fF
XC743 G1011.t112 GND 0.13fF
XC744 G1011.n439 GND 0.12fF
XC745 G1011.n440 GND 0.12fF
XC746 G1011.n441 GND 0.10fF
XC747 G1011.n442 GND 0.05fF
XC748 G1011.n443 GND 0.01fF
XC749 G1011.n444 GND 0.02fF
XC750 G1011.t5 GND 0.02fF
XC751 G1011.t39 GND 0.02fF
XC752 G1011.n450 GND 0.06fF
XC753 G1011.n451 GND 0.01fF
XC754 G1011.n452 GND 0.14fF
XC755 G1011.n453 GND 0.11fF
XC756 G1011.n454 GND 0.05fF
XC757 G1011.n455 GND 0.05fF
XC758 G1011.t80 GND 0.13fF
XC759 G1011.n456 GND 0.10fF
XC760 G1011.t2 GND 0.13fF
XC761 G1011.n457 GND 0.10fF
XC762 G1011.n458 GND 0.05fF
XC763 G1011.n459 GND 0.01fF
XC764 G1011.n460 GND 0.02fF
XC765 G1011.t81 GND 0.02fF
XC766 G1011.t3 GND 0.02fF
XC767 G1011.n466 GND 0.06fF
XC768 G1011.n467 GND 0.01fF
XC769 G1011.n468 GND 0.14fF
XC770 G1011.n469 GND 0.11fF
XC771 G1011.n470 GND 0.05fF
XC772 G1011.n471 GND 0.05fF
XC773 G1011.t8 GND 0.13fF
XC774 G1011.n472 GND 0.10fF
XC775 G1011.t42 GND 0.13fF
XC776 G1011.n473 GND 0.10fF
XC777 G1011.n474 GND 0.05fF
XC778 G1011.n475 GND 0.01fF
XC779 G1011.n476 GND 0.02fF
XC780 G1011.t9 GND 0.02fF
XC781 G1011.t43 GND 0.02fF
XC782 G1011.n482 GND 0.06fF
XC783 G1011.n483 GND 0.01fF
XC784 G1011.n484 GND 0.14fF
XC785 G1011.n485 GND 0.11fF
XC786 G1011.n486 GND 0.05fF
XC787 G1011.n487 GND 0.05fF
XC788 G1011.t54 GND 0.13fF
XC789 G1011.n488 GND 0.10fF
XC790 G1011.t62 GND 0.13fF
XC791 G1011.n489 GND 0.10fF
XC792 G1011.n490 GND 0.05fF
XC793 G1011.n491 GND 0.01fF
XC794 G1011.n492 GND 0.02fF
XC795 G1011.t55 GND 0.02fF
XC796 G1011.t63 GND 0.02fF
XC797 G1011.n498 GND 0.06fF
XC798 G1011.n499 GND 0.01fF
XC799 G1011.n500 GND 0.14fF
XC800 G1011.n501 GND 0.11fF
XC801 G1011.n502 GND 0.05fF
XC802 G1011.n503 GND 0.05fF
XC803 G1011.t0 GND 0.13fF
XC804 G1011.n504 GND 0.10fF
XC805 G1011.t26 GND 0.13fF
XC806 G1011.n505 GND 0.10fF
XC807 G1011.n506 GND 0.05fF
XC808 G1011.n507 GND 0.01fF
XC809 G1011.n508 GND 0.02fF
XC810 G1011.t1 GND 0.02fF
XC811 G1011.t27 GND 0.02fF
XC812 G1011.n514 GND 0.06fF
XC813 G1011.n515 GND 0.01fF
XC814 G1011.n516 GND 0.14fF
XC815 G1011.n517 GND 0.11fF
XC816 G1011.n518 GND 0.05fF
XC817 G1011.n519 GND 0.05fF
XC818 G1011.t50 GND 0.13fF
XC819 G1011.n520 GND 0.10fF
XC820 G1011.t60 GND 0.13fF
XC821 G1011.n521 GND 0.10fF
XC822 G1011.n522 GND 0.05fF
XC823 G1011.n523 GND 0.01fF
XC824 G1011.n524 GND 0.02fF
XC825 G1011.t51 GND 0.02fF
XC826 G1011.t61 GND 0.02fF
XC827 G1011.n530 GND 0.06fF
XC828 G1011.n531 GND 0.01fF
XC829 G1011.n532 GND 0.14fF
XC830 G1011.n533 GND 0.11fF
XC831 G1011.n534 GND 0.05fF
XC832 G1011.n535 GND 0.05fF
XC833 G1011.t84 GND 0.13fF
XC834 G1011.n536 GND 0.10fF
XC835 G1011.t24 GND 0.13fF
XC836 G1011.n537 GND 0.10fF
XC837 G1011.n538 GND 0.05fF
XC838 G1011.n539 GND 0.01fF
XC839 G1011.n540 GND 0.02fF
XC840 G1011.t85 GND 0.02fF
XC841 G1011.t25 GND 0.02fF
XC842 G1011.n546 GND 0.06fF
XC843 G1011.n547 GND 0.01fF
XC844 G1011.n548 GND 0.14fF
XC845 G1011.n549 GND 0.11fF
XC846 G1011.n550 GND 0.05fF
XC847 G1011.n551 GND 0.05fF
XC848 G1011.t16 GND 0.13fF
XC849 G1011.n552 GND 0.10fF
XC850 G1011.t46 GND 0.13fF
XC851 G1011.n553 GND 0.10fF
XC852 G1011.n554 GND 0.05fF
XC853 G1011.n555 GND 0.01fF
XC854 G1011.n556 GND 0.02fF
XC855 G1011.t17 GND 0.02fF
XC856 G1011.t47 GND 0.02fF
XC857 G1011.n562 GND 0.06fF
XC858 G1011.n563 GND 0.01fF
XC859 G1011.n564 GND 0.14fF
XC860 G1011.n565 GND 0.11fF
XC861 G1011.n566 GND 0.05fF
XC862 G1011.n567 GND 0.05fF
XC863 G1011.n568 GND 0.01fF
XC864 G1011.n569 GND 0.02fF
XC865 G1011.t83 GND 0.02fF
XC866 G1011.t23 GND 0.02fF
XC867 G1011.n575 GND 0.06fF
XC868 G1011.n576 GND 0.01fF
XC869 G1011.n577 GND 0.14fF
XC870 G1011.n578 GND 0.11fF
XC871 G1011.n579 GND 0.05fF
XC872 G1011.n580 GND 0.05fF
XC873 G1011.n583 GND 0.01fF
XC874 G1011.n584 GND 0.14fF
XC875 G1011.n585 GND 0.11fF
XC876 G1011.n586 GND 0.05fF
XC877 G1011.n587 GND 1.26fF
.ends


** flattened .save nodes
.end
