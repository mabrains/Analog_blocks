magic
tech sky130A
magscale 1 2
timestamp 1624883981
<< checkpaint >>
rect -1260 -1260 3542 3598
<< pwell >>
rect 1176 1289 1197 1338
<< metal1 >>
rect 0 2331 2282 2338
rect 0 2282 88 2331
rect 0 2230 7 2282
rect 59 2279 88 2282
rect 140 2279 152 2331
rect 204 2279 216 2331
rect 268 2279 280 2331
rect 332 2279 344 2331
rect 396 2279 408 2331
rect 460 2279 472 2331
rect 524 2279 536 2331
rect 588 2279 600 2331
rect 652 2279 664 2331
rect 716 2279 728 2331
rect 780 2279 792 2331
rect 844 2279 856 2331
rect 908 2279 920 2331
rect 972 2279 984 2331
rect 1036 2279 1246 2331
rect 1298 2279 1310 2331
rect 1362 2279 1374 2331
rect 1426 2279 1438 2331
rect 1490 2279 1502 2331
rect 1554 2279 1566 2331
rect 1618 2279 1630 2331
rect 1682 2279 1694 2331
rect 1746 2279 1758 2331
rect 1810 2279 1822 2331
rect 1874 2279 1886 2331
rect 1938 2279 1950 2331
rect 2002 2279 2014 2331
rect 2066 2279 2078 2331
rect 2130 2279 2142 2331
rect 2194 2282 2282 2331
rect 2194 2279 2223 2282
rect 59 2272 2223 2279
rect 59 2230 72 2272
rect 0 2218 72 2230
rect 0 2166 7 2218
rect 59 2166 72 2218
rect 0 2154 72 2166
rect 0 2102 7 2154
rect 59 2102 72 2154
rect 0 2090 72 2102
rect 0 2038 7 2090
rect 59 2038 72 2090
rect 0 2026 72 2038
rect 0 1974 7 2026
rect 59 1974 72 2026
rect 0 1962 72 1974
rect 0 1910 7 1962
rect 59 1910 72 1962
rect 0 1898 72 1910
rect 0 1846 7 1898
rect 59 1846 72 1898
rect 0 1834 72 1846
rect 0 1782 7 1834
rect 59 1782 72 1834
rect 0 1770 72 1782
rect 0 1718 7 1770
rect 59 1718 72 1770
rect 0 1706 72 1718
rect 0 1654 7 1706
rect 59 1654 72 1706
rect 0 1642 72 1654
rect 0 1590 7 1642
rect 59 1590 72 1642
rect 0 1578 72 1590
rect 0 1526 7 1578
rect 59 1526 72 1578
rect 0 1514 72 1526
rect 0 1462 7 1514
rect 59 1462 72 1514
rect 0 1450 72 1462
rect 0 1398 7 1450
rect 59 1398 72 1450
rect 0 1386 72 1398
rect 0 1334 7 1386
rect 59 1334 72 1386
rect 0 1322 72 1334
rect 0 1270 7 1322
rect 59 1270 72 1322
rect 0 1068 72 1270
rect 0 1016 7 1068
rect 59 1016 72 1068
rect 0 1004 72 1016
rect 0 952 7 1004
rect 59 952 72 1004
rect 0 940 72 952
rect 0 888 7 940
rect 59 888 72 940
rect 0 876 72 888
rect 0 824 7 876
rect 59 824 72 876
rect 0 812 72 824
rect 0 760 7 812
rect 59 760 72 812
rect 0 748 72 760
rect 0 696 7 748
rect 59 696 72 748
rect 0 684 72 696
rect 0 632 7 684
rect 59 632 72 684
rect 0 620 72 632
rect 0 568 7 620
rect 59 568 72 620
rect 0 556 72 568
rect 0 504 7 556
rect 59 504 72 556
rect 0 492 72 504
rect 0 440 7 492
rect 59 440 72 492
rect 0 428 72 440
rect 0 376 7 428
rect 59 376 72 428
rect 0 364 72 376
rect 0 312 7 364
rect 59 312 72 364
rect 0 300 72 312
rect 0 248 7 300
rect 59 248 72 300
rect 0 236 72 248
rect 0 184 7 236
rect 59 184 72 236
rect 0 172 72 184
rect 0 120 7 172
rect 59 120 72 172
rect 0 108 72 120
rect 0 56 7 108
rect 59 66 72 108
rect 100 1201 128 2244
rect 156 1229 184 2272
rect 212 1201 240 2244
rect 268 1229 296 2272
rect 324 1201 352 2244
rect 380 1229 408 2272
rect 436 1201 464 2244
rect 492 1229 520 2272
rect 548 1201 576 2244
rect 604 1229 632 2272
rect 660 1201 688 2244
rect 716 1229 744 2272
rect 772 1201 800 2244
rect 828 1229 856 2272
rect 884 1201 912 2244
rect 940 1229 968 2272
rect 996 1201 1024 2244
rect 1052 1229 1080 2272
rect 1108 2237 1174 2244
rect 1108 2185 1115 2237
rect 1167 2185 1174 2237
rect 1108 2173 1174 2185
rect 1108 2121 1115 2173
rect 1167 2121 1174 2173
rect 1108 2109 1174 2121
rect 1108 2057 1115 2109
rect 1167 2057 1174 2109
rect 1108 2045 1174 2057
rect 1108 1993 1115 2045
rect 1167 1993 1174 2045
rect 1108 1981 1174 1993
rect 1108 1929 1115 1981
rect 1167 1929 1174 1981
rect 1108 1917 1174 1929
rect 1108 1865 1115 1917
rect 1167 1865 1174 1917
rect 1108 1853 1174 1865
rect 1108 1801 1115 1853
rect 1167 1801 1174 1853
rect 1108 1789 1174 1801
rect 1108 1737 1115 1789
rect 1167 1737 1174 1789
rect 1108 1725 1174 1737
rect 1108 1673 1115 1725
rect 1167 1673 1174 1725
rect 1108 1661 1174 1673
rect 1108 1609 1115 1661
rect 1167 1609 1174 1661
rect 1108 1597 1174 1609
rect 1108 1545 1115 1597
rect 1167 1545 1174 1597
rect 1108 1533 1174 1545
rect 1108 1481 1115 1533
rect 1167 1481 1174 1533
rect 1108 1469 1174 1481
rect 1108 1417 1115 1469
rect 1167 1417 1174 1469
rect 1108 1405 1174 1417
rect 1108 1353 1115 1405
rect 1167 1353 1174 1405
rect 1108 1341 1174 1353
rect 1108 1289 1115 1341
rect 1167 1289 1174 1341
rect 1108 1277 1174 1289
rect 1108 1225 1115 1277
rect 1167 1225 1174 1277
rect 1202 1229 1230 2272
rect 1108 1201 1174 1225
rect 1258 1201 1286 2244
rect 1314 1229 1342 2272
rect 1370 1201 1398 2244
rect 1426 1229 1454 2272
rect 1482 1201 1510 2244
rect 1538 1229 1566 2272
rect 1594 1201 1622 2244
rect 1650 1229 1678 2272
rect 1706 1201 1734 2244
rect 1762 1229 1790 2272
rect 1818 1201 1846 2244
rect 1874 1229 1902 2272
rect 1930 1201 1958 2244
rect 1986 1229 2014 2272
rect 2042 1201 2070 2244
rect 2098 1229 2126 2272
rect 2154 1201 2182 2244
rect 100 1195 2182 1201
rect 100 1143 152 1195
rect 204 1143 216 1195
rect 268 1143 280 1195
rect 332 1143 344 1195
rect 396 1143 408 1195
rect 460 1143 472 1195
rect 524 1143 536 1195
rect 588 1143 600 1195
rect 652 1143 664 1195
rect 716 1143 728 1195
rect 780 1143 792 1195
rect 844 1143 856 1195
rect 908 1143 920 1195
rect 972 1143 984 1195
rect 1036 1143 1048 1195
rect 1100 1143 1182 1195
rect 1234 1143 1246 1195
rect 1298 1143 1310 1195
rect 1362 1143 1374 1195
rect 1426 1143 1438 1195
rect 1490 1143 1502 1195
rect 1554 1143 1566 1195
rect 1618 1143 1630 1195
rect 1682 1143 1694 1195
rect 1746 1143 1758 1195
rect 1810 1143 1822 1195
rect 1874 1143 1886 1195
rect 1938 1143 1950 1195
rect 2002 1143 2014 1195
rect 2066 1143 2078 1195
rect 2130 1143 2182 1195
rect 100 1137 2182 1143
rect 100 94 128 1137
rect 156 66 184 1109
rect 212 94 240 1137
rect 268 66 296 1109
rect 324 94 352 1137
rect 380 66 408 1109
rect 436 94 464 1137
rect 492 66 520 1109
rect 548 94 576 1137
rect 604 66 632 1109
rect 660 94 688 1137
rect 716 66 744 1109
rect 772 94 800 1137
rect 828 66 856 1109
rect 884 94 912 1137
rect 940 66 968 1109
rect 996 94 1024 1137
rect 1108 1113 1174 1137
rect 1052 66 1080 1109
rect 1108 1061 1115 1113
rect 1167 1061 1174 1113
rect 1108 1049 1174 1061
rect 1108 997 1115 1049
rect 1167 997 1174 1049
rect 1108 985 1174 997
rect 1108 933 1115 985
rect 1167 933 1174 985
rect 1108 921 1174 933
rect 1108 869 1115 921
rect 1167 869 1174 921
rect 1108 857 1174 869
rect 1108 805 1115 857
rect 1167 805 1174 857
rect 1108 793 1174 805
rect 1108 741 1115 793
rect 1167 741 1174 793
rect 1108 729 1174 741
rect 1108 677 1115 729
rect 1167 677 1174 729
rect 1108 665 1174 677
rect 1108 613 1115 665
rect 1167 613 1174 665
rect 1108 601 1174 613
rect 1108 549 1115 601
rect 1167 549 1174 601
rect 1108 537 1174 549
rect 1108 485 1115 537
rect 1167 485 1174 537
rect 1108 473 1174 485
rect 1108 421 1115 473
rect 1167 421 1174 473
rect 1108 409 1174 421
rect 1108 357 1115 409
rect 1167 357 1174 409
rect 1108 345 1174 357
rect 1108 293 1115 345
rect 1167 293 1174 345
rect 1108 281 1174 293
rect 1108 229 1115 281
rect 1167 229 1174 281
rect 1108 217 1174 229
rect 1108 165 1115 217
rect 1167 165 1174 217
rect 1108 153 1174 165
rect 1108 101 1115 153
rect 1167 101 1174 153
rect 1108 94 1174 101
rect 1202 66 1230 1109
rect 1258 94 1286 1137
rect 1314 66 1342 1109
rect 1370 94 1398 1137
rect 1426 66 1454 1109
rect 1482 94 1510 1137
rect 1538 66 1566 1109
rect 1594 94 1622 1137
rect 1650 66 1678 1109
rect 1706 94 1734 1137
rect 1762 66 1790 1109
rect 1818 94 1846 1137
rect 1874 66 1902 1109
rect 1930 94 1958 1137
rect 1986 66 2014 1109
rect 2042 94 2070 1137
rect 2098 66 2126 1109
rect 2154 94 2182 1137
rect 2210 2230 2223 2272
rect 2275 2230 2282 2282
rect 2210 2218 2282 2230
rect 2210 2166 2223 2218
rect 2275 2166 2282 2218
rect 2210 2154 2282 2166
rect 2210 2102 2223 2154
rect 2275 2102 2282 2154
rect 2210 2090 2282 2102
rect 2210 2038 2223 2090
rect 2275 2038 2282 2090
rect 2210 2026 2282 2038
rect 2210 1974 2223 2026
rect 2275 1974 2282 2026
rect 2210 1962 2282 1974
rect 2210 1910 2223 1962
rect 2275 1910 2282 1962
rect 2210 1898 2282 1910
rect 2210 1846 2223 1898
rect 2275 1846 2282 1898
rect 2210 1834 2282 1846
rect 2210 1782 2223 1834
rect 2275 1782 2282 1834
rect 2210 1770 2282 1782
rect 2210 1718 2223 1770
rect 2275 1718 2282 1770
rect 2210 1706 2282 1718
rect 2210 1654 2223 1706
rect 2275 1654 2282 1706
rect 2210 1642 2282 1654
rect 2210 1590 2223 1642
rect 2275 1590 2282 1642
rect 2210 1578 2282 1590
rect 2210 1526 2223 1578
rect 2275 1526 2282 1578
rect 2210 1514 2282 1526
rect 2210 1462 2223 1514
rect 2275 1462 2282 1514
rect 2210 1450 2282 1462
rect 2210 1398 2223 1450
rect 2275 1398 2282 1450
rect 2210 1386 2282 1398
rect 2210 1334 2223 1386
rect 2275 1334 2282 1386
rect 2210 1322 2282 1334
rect 2210 1270 2223 1322
rect 2275 1270 2282 1322
rect 2210 1068 2282 1270
rect 2210 1016 2223 1068
rect 2275 1016 2282 1068
rect 2210 1004 2282 1016
rect 2210 952 2223 1004
rect 2275 952 2282 1004
rect 2210 940 2282 952
rect 2210 888 2223 940
rect 2275 888 2282 940
rect 2210 876 2282 888
rect 2210 824 2223 876
rect 2275 824 2282 876
rect 2210 812 2282 824
rect 2210 760 2223 812
rect 2275 760 2282 812
rect 2210 748 2282 760
rect 2210 696 2223 748
rect 2275 696 2282 748
rect 2210 684 2282 696
rect 2210 632 2223 684
rect 2275 632 2282 684
rect 2210 620 2282 632
rect 2210 568 2223 620
rect 2275 568 2282 620
rect 2210 556 2282 568
rect 2210 504 2223 556
rect 2275 504 2282 556
rect 2210 492 2282 504
rect 2210 440 2223 492
rect 2275 440 2282 492
rect 2210 428 2282 440
rect 2210 376 2223 428
rect 2275 376 2282 428
rect 2210 364 2282 376
rect 2210 312 2223 364
rect 2275 312 2282 364
rect 2210 300 2282 312
rect 2210 248 2223 300
rect 2275 248 2282 300
rect 2210 236 2282 248
rect 2210 184 2223 236
rect 2275 184 2282 236
rect 2210 172 2282 184
rect 2210 120 2223 172
rect 2275 120 2282 172
rect 2210 108 2282 120
rect 2210 66 2223 108
rect 59 59 2223 66
rect 59 56 88 59
rect 0 7 88 56
rect 140 7 152 59
rect 204 7 216 59
rect 268 7 280 59
rect 332 7 344 59
rect 396 7 408 59
rect 460 7 472 59
rect 524 7 536 59
rect 588 7 600 59
rect 652 7 664 59
rect 716 7 728 59
rect 780 7 792 59
rect 844 7 856 59
rect 908 7 920 59
rect 972 7 984 59
rect 1036 7 1246 59
rect 1298 7 1310 59
rect 1362 7 1374 59
rect 1426 7 1438 59
rect 1490 7 1502 59
rect 1554 7 1566 59
rect 1618 7 1630 59
rect 1682 7 1694 59
rect 1746 7 1758 59
rect 1810 7 1822 59
rect 1874 7 1886 59
rect 1938 7 1950 59
rect 2002 7 2014 59
rect 2066 7 2078 59
rect 2130 7 2142 59
rect 2194 56 2223 59
rect 2275 56 2282 108
rect 2194 7 2282 56
rect 0 0 2282 7
<< via1 >>
rect 7 2230 59 2282
rect 88 2279 140 2331
rect 152 2279 204 2331
rect 216 2279 268 2331
rect 280 2279 332 2331
rect 344 2279 396 2331
rect 408 2279 460 2331
rect 472 2279 524 2331
rect 536 2279 588 2331
rect 600 2279 652 2331
rect 664 2279 716 2331
rect 728 2279 780 2331
rect 792 2279 844 2331
rect 856 2279 908 2331
rect 920 2279 972 2331
rect 984 2279 1036 2331
rect 1246 2279 1298 2331
rect 1310 2279 1362 2331
rect 1374 2279 1426 2331
rect 1438 2279 1490 2331
rect 1502 2279 1554 2331
rect 1566 2279 1618 2331
rect 1630 2279 1682 2331
rect 1694 2279 1746 2331
rect 1758 2279 1810 2331
rect 1822 2279 1874 2331
rect 1886 2279 1938 2331
rect 1950 2279 2002 2331
rect 2014 2279 2066 2331
rect 2078 2279 2130 2331
rect 2142 2279 2194 2331
rect 7 2166 59 2218
rect 7 2102 59 2154
rect 7 2038 59 2090
rect 7 1974 59 2026
rect 7 1910 59 1962
rect 7 1846 59 1898
rect 7 1782 59 1834
rect 7 1718 59 1770
rect 7 1654 59 1706
rect 7 1590 59 1642
rect 7 1526 59 1578
rect 7 1462 59 1514
rect 7 1398 59 1450
rect 7 1334 59 1386
rect 7 1270 59 1322
rect 7 1016 59 1068
rect 7 952 59 1004
rect 7 888 59 940
rect 7 824 59 876
rect 7 760 59 812
rect 7 696 59 748
rect 7 632 59 684
rect 7 568 59 620
rect 7 504 59 556
rect 7 440 59 492
rect 7 376 59 428
rect 7 312 59 364
rect 7 248 59 300
rect 7 184 59 236
rect 7 120 59 172
rect 7 56 59 108
rect 1115 2185 1167 2237
rect 1115 2121 1167 2173
rect 1115 2057 1167 2109
rect 1115 1993 1167 2045
rect 1115 1929 1167 1981
rect 1115 1865 1167 1917
rect 1115 1801 1167 1853
rect 1115 1737 1167 1789
rect 1115 1673 1167 1725
rect 1115 1609 1167 1661
rect 1115 1545 1167 1597
rect 1115 1481 1167 1533
rect 1115 1417 1167 1469
rect 1115 1353 1167 1405
rect 1115 1289 1167 1341
rect 1115 1225 1167 1277
rect 152 1143 204 1195
rect 216 1143 268 1195
rect 280 1143 332 1195
rect 344 1143 396 1195
rect 408 1143 460 1195
rect 472 1143 524 1195
rect 536 1143 588 1195
rect 600 1143 652 1195
rect 664 1143 716 1195
rect 728 1143 780 1195
rect 792 1143 844 1195
rect 856 1143 908 1195
rect 920 1143 972 1195
rect 984 1143 1036 1195
rect 1048 1143 1100 1195
rect 1182 1143 1234 1195
rect 1246 1143 1298 1195
rect 1310 1143 1362 1195
rect 1374 1143 1426 1195
rect 1438 1143 1490 1195
rect 1502 1143 1554 1195
rect 1566 1143 1618 1195
rect 1630 1143 1682 1195
rect 1694 1143 1746 1195
rect 1758 1143 1810 1195
rect 1822 1143 1874 1195
rect 1886 1143 1938 1195
rect 1950 1143 2002 1195
rect 2014 1143 2066 1195
rect 2078 1143 2130 1195
rect 1115 1061 1167 1113
rect 1115 997 1167 1049
rect 1115 933 1167 985
rect 1115 869 1167 921
rect 1115 805 1167 857
rect 1115 741 1167 793
rect 1115 677 1167 729
rect 1115 613 1167 665
rect 1115 549 1167 601
rect 1115 485 1167 537
rect 1115 421 1167 473
rect 1115 357 1167 409
rect 1115 293 1167 345
rect 1115 229 1167 281
rect 1115 165 1167 217
rect 1115 101 1167 153
rect 2223 2230 2275 2282
rect 2223 2166 2275 2218
rect 2223 2102 2275 2154
rect 2223 2038 2275 2090
rect 2223 1974 2275 2026
rect 2223 1910 2275 1962
rect 2223 1846 2275 1898
rect 2223 1782 2275 1834
rect 2223 1718 2275 1770
rect 2223 1654 2275 1706
rect 2223 1590 2275 1642
rect 2223 1526 2275 1578
rect 2223 1462 2275 1514
rect 2223 1398 2275 1450
rect 2223 1334 2275 1386
rect 2223 1270 2275 1322
rect 2223 1016 2275 1068
rect 2223 952 2275 1004
rect 2223 888 2275 940
rect 2223 824 2275 876
rect 2223 760 2275 812
rect 2223 696 2275 748
rect 2223 632 2275 684
rect 2223 568 2275 620
rect 2223 504 2275 556
rect 2223 440 2275 492
rect 2223 376 2275 428
rect 2223 312 2275 364
rect 2223 248 2275 300
rect 2223 184 2275 236
rect 2223 120 2275 172
rect 88 7 140 59
rect 152 7 204 59
rect 216 7 268 59
rect 280 7 332 59
rect 344 7 396 59
rect 408 7 460 59
rect 472 7 524 59
rect 536 7 588 59
rect 600 7 652 59
rect 664 7 716 59
rect 728 7 780 59
rect 792 7 844 59
rect 856 7 908 59
rect 920 7 972 59
rect 984 7 1036 59
rect 1246 7 1298 59
rect 1310 7 1362 59
rect 1374 7 1426 59
rect 1438 7 1490 59
rect 1502 7 1554 59
rect 1566 7 1618 59
rect 1630 7 1682 59
rect 1694 7 1746 59
rect 1758 7 1810 59
rect 1822 7 1874 59
rect 1886 7 1938 59
rect 1950 7 2002 59
rect 2014 7 2066 59
rect 2078 7 2130 59
rect 2142 7 2194 59
rect 2223 56 2275 108
<< metal2 >>
rect 0 2333 1086 2338
rect 0 2282 61 2333
rect 117 2331 141 2333
rect 197 2331 221 2333
rect 277 2331 301 2333
rect 357 2331 381 2333
rect 437 2331 461 2333
rect 517 2331 541 2333
rect 597 2331 621 2333
rect 677 2331 701 2333
rect 757 2331 781 2333
rect 837 2331 861 2333
rect 917 2331 941 2333
rect 997 2331 1021 2333
rect 0 2249 7 2282
rect 59 2277 61 2282
rect 140 2279 141 2331
rect 204 2279 216 2331
rect 277 2279 280 2331
rect 460 2279 461 2331
rect 524 2279 536 2331
rect 597 2279 600 2331
rect 780 2279 781 2331
rect 844 2279 856 2331
rect 917 2279 920 2331
rect 117 2277 141 2279
rect 197 2277 221 2279
rect 277 2277 301 2279
rect 357 2277 381 2279
rect 437 2277 461 2279
rect 517 2277 541 2279
rect 597 2277 621 2279
rect 677 2277 701 2279
rect 757 2277 781 2279
rect 837 2277 861 2279
rect 917 2277 941 2279
rect 997 2277 1021 2279
rect 1077 2277 1086 2333
rect 59 2272 1086 2277
rect 59 2249 66 2272
rect 0 2193 5 2249
rect 61 2193 66 2249
rect 1114 2244 1168 2338
rect 1196 2333 2282 2338
rect 1196 2277 1205 2333
rect 1261 2331 1285 2333
rect 1341 2331 1365 2333
rect 1421 2331 1445 2333
rect 1501 2331 1525 2333
rect 1581 2331 1605 2333
rect 1661 2331 1685 2333
rect 1741 2331 1765 2333
rect 1821 2331 1845 2333
rect 1901 2331 1925 2333
rect 1981 2331 2005 2333
rect 2061 2331 2085 2333
rect 2141 2331 2165 2333
rect 1362 2279 1365 2331
rect 1426 2279 1438 2331
rect 1501 2279 1502 2331
rect 1682 2279 1685 2331
rect 1746 2279 1758 2331
rect 1821 2279 1822 2331
rect 2002 2279 2005 2331
rect 2066 2279 2078 2331
rect 2141 2279 2142 2331
rect 2221 2282 2282 2333
rect 1261 2277 1285 2279
rect 1341 2277 1365 2279
rect 1421 2277 1445 2279
rect 1501 2277 1525 2279
rect 1581 2277 1605 2279
rect 1661 2277 1685 2279
rect 1741 2277 1765 2279
rect 1821 2277 1845 2279
rect 1901 2277 1925 2279
rect 1981 2277 2005 2279
rect 2061 2277 2085 2279
rect 2141 2277 2165 2279
rect 2221 2277 2223 2282
rect 1196 2272 2223 2277
rect 2216 2249 2223 2272
rect 2275 2249 2282 2282
rect 94 2237 2188 2244
rect 94 2216 1115 2237
rect 0 2169 7 2193
rect 59 2188 66 2193
rect 59 2169 1085 2188
rect 0 2113 5 2169
rect 61 2160 1085 2169
rect 1113 2185 1115 2216
rect 1167 2216 2188 2237
rect 1167 2185 1169 2216
rect 2216 2193 2221 2249
rect 2277 2193 2282 2249
rect 2216 2188 2223 2193
rect 1113 2173 1169 2185
rect 61 2113 66 2160
rect 1113 2157 1115 2173
rect 1167 2157 1169 2173
rect 1197 2169 2223 2188
rect 2275 2169 2282 2193
rect 1197 2160 2221 2169
rect 0 2102 7 2113
rect 59 2102 66 2113
rect 94 2104 1113 2132
rect 0 2090 66 2102
rect 0 2089 7 2090
rect 59 2089 66 2090
rect 0 2033 5 2089
rect 61 2076 66 2089
rect 1169 2104 2188 2132
rect 2216 2113 2221 2160
rect 2277 2113 2282 2169
rect 1113 2077 1115 2101
rect 1167 2077 1169 2101
rect 61 2048 1085 2076
rect 2216 2102 2223 2113
rect 2275 2102 2282 2113
rect 2216 2090 2282 2102
rect 2216 2089 2223 2090
rect 2275 2089 2282 2090
rect 2216 2076 2221 2089
rect 61 2033 66 2048
rect 0 2026 66 2033
rect 0 2009 7 2026
rect 59 2009 66 2026
rect 1197 2048 2221 2076
rect 1113 2020 1115 2021
rect 0 1953 5 2009
rect 61 1964 66 2009
rect 94 1997 1115 2020
rect 1167 2020 1169 2021
rect 2216 2033 2221 2048
rect 2277 2033 2282 2089
rect 2216 2026 2282 2033
rect 1167 1997 2188 2020
rect 94 1992 1113 1997
rect 1169 1992 2188 1997
rect 2216 2009 2223 2026
rect 2275 2009 2282 2026
rect 61 1953 1085 1964
rect 0 1929 7 1953
rect 59 1936 1085 1953
rect 2216 1964 2221 2009
rect 59 1929 66 1936
rect 0 1873 5 1929
rect 61 1873 66 1929
rect 1113 1929 1115 1941
rect 1167 1929 1169 1941
rect 1197 1953 2221 1964
rect 2277 1953 2282 2009
rect 1197 1936 2223 1953
rect 1113 1917 1169 1929
rect 94 1880 1113 1908
rect 0 1849 7 1873
rect 59 1852 66 1873
rect 2216 1929 2223 1936
rect 2275 1929 2282 1953
rect 1169 1880 2188 1908
rect 1113 1853 1169 1861
rect 59 1849 1085 1852
rect 0 1793 5 1849
rect 61 1824 1085 1849
rect 1113 1837 1115 1853
rect 1167 1837 1169 1853
rect 2216 1873 2221 1929
rect 2277 1873 2282 1929
rect 2216 1852 2223 1873
rect 61 1793 66 1824
rect 1197 1849 2223 1852
rect 2275 1849 2282 1873
rect 1197 1824 2221 1849
rect 0 1782 7 1793
rect 59 1782 66 1793
rect 0 1770 66 1782
rect 0 1769 7 1770
rect 59 1769 66 1770
rect 0 1713 5 1769
rect 61 1740 66 1769
rect 94 1781 1113 1796
rect 1169 1781 2188 1796
rect 94 1768 1115 1781
rect 1113 1757 1115 1768
rect 1167 1768 2188 1781
rect 2216 1793 2221 1824
rect 2277 1793 2282 1849
rect 2216 1782 2223 1793
rect 2275 1782 2282 1793
rect 2216 1770 2282 1782
rect 2216 1769 2223 1770
rect 2275 1769 2282 1770
rect 1167 1757 1169 1768
rect 61 1713 1085 1740
rect 0 1712 1085 1713
rect 2216 1740 2221 1769
rect 0 1706 66 1712
rect 0 1689 7 1706
rect 59 1689 66 1706
rect 0 1633 5 1689
rect 61 1633 66 1689
rect 1197 1713 2221 1740
rect 2277 1713 2282 1769
rect 1197 1712 2282 1713
rect 1113 1684 1115 1701
rect 94 1677 1115 1684
rect 1167 1684 1169 1701
rect 2216 1706 2282 1712
rect 2216 1689 2223 1706
rect 2275 1689 2282 1706
rect 1167 1677 2188 1684
rect 94 1656 1113 1677
rect 0 1609 7 1633
rect 59 1628 66 1633
rect 59 1609 1085 1628
rect 0 1553 5 1609
rect 61 1600 1085 1609
rect 1169 1656 2188 1677
rect 2216 1633 2221 1689
rect 2277 1633 2282 1689
rect 2216 1628 2223 1633
rect 1113 1609 1115 1621
rect 1167 1609 1169 1621
rect 61 1553 66 1600
rect 1113 1597 1169 1609
rect 1197 1609 2223 1628
rect 2275 1609 2282 1633
rect 1197 1600 2221 1609
rect 0 1529 7 1553
rect 59 1529 66 1553
rect 94 1544 1113 1572
rect 0 1473 5 1529
rect 61 1516 66 1529
rect 1169 1544 2188 1572
rect 2216 1553 2221 1600
rect 2277 1553 2282 1609
rect 1113 1533 1169 1541
rect 1113 1517 1115 1533
rect 1167 1517 1169 1533
rect 61 1488 1085 1516
rect 61 1473 66 1488
rect 0 1462 7 1473
rect 59 1462 66 1473
rect 0 1450 66 1462
rect 2216 1529 2223 1553
rect 2275 1529 2282 1553
rect 2216 1516 2221 1529
rect 1197 1488 2221 1516
rect 1113 1460 1115 1461
rect 0 1449 7 1450
rect 59 1449 66 1450
rect 0 1393 5 1449
rect 61 1404 66 1449
rect 94 1437 1115 1460
rect 1167 1460 1169 1461
rect 2216 1473 2221 1488
rect 2277 1473 2282 1529
rect 2216 1462 2223 1473
rect 2275 1462 2282 1473
rect 1167 1437 2188 1460
rect 94 1432 1113 1437
rect 1169 1432 2188 1437
rect 2216 1450 2282 1462
rect 2216 1449 2223 1450
rect 2275 1449 2282 1450
rect 61 1393 1085 1404
rect 0 1386 1085 1393
rect 0 1369 7 1386
rect 59 1376 1085 1386
rect 2216 1404 2221 1449
rect 59 1369 66 1376
rect 0 1313 5 1369
rect 61 1313 66 1369
rect 1113 1357 1115 1381
rect 1167 1357 1169 1381
rect 1197 1393 2221 1404
rect 2277 1393 2282 1449
rect 1197 1386 2282 1393
rect 1197 1376 2223 1386
rect 94 1320 1113 1348
rect 2216 1369 2223 1376
rect 2275 1369 2282 1386
rect 0 1289 7 1313
rect 59 1292 66 1313
rect 1169 1320 2188 1348
rect 59 1289 1085 1292
rect 0 1233 5 1289
rect 61 1233 1085 1289
rect 0 1225 1085 1233
rect 1113 1289 1115 1301
rect 1167 1289 1169 1301
rect 2216 1313 2221 1369
rect 2277 1313 2282 1369
rect 2216 1292 2223 1313
rect 1113 1277 1169 1289
rect 1197 1289 2223 1292
rect 2275 1289 2282 1313
rect 1197 1233 2221 1289
rect 2277 1233 2282 1289
rect 1197 1225 2282 1233
rect 0 1224 66 1225
rect 2216 1224 2282 1225
rect 1113 1197 1169 1221
rect 74 1196 153 1197
rect 0 1195 153 1196
rect 209 1195 233 1197
rect 289 1195 313 1197
rect 369 1195 393 1197
rect 449 1195 473 1197
rect 529 1195 553 1197
rect 609 1195 633 1197
rect 689 1195 713 1197
rect 769 1195 793 1197
rect 849 1195 873 1197
rect 929 1195 953 1197
rect 1009 1195 1033 1197
rect 1089 1195 1113 1197
rect 0 1143 152 1195
rect 209 1143 216 1195
rect 460 1143 472 1195
rect 529 1143 536 1195
rect 780 1143 792 1195
rect 849 1143 856 1195
rect 1100 1143 1113 1195
rect 0 1142 153 1143
rect 74 1141 153 1142
rect 209 1141 233 1143
rect 289 1141 313 1143
rect 369 1141 393 1143
rect 449 1141 473 1143
rect 529 1141 553 1143
rect 609 1141 633 1143
rect 689 1141 713 1143
rect 769 1141 793 1143
rect 849 1141 873 1143
rect 929 1141 953 1143
rect 1009 1141 1033 1143
rect 1089 1141 1113 1143
rect 1169 1195 1193 1197
rect 1249 1195 1273 1197
rect 1329 1195 1353 1197
rect 1409 1195 1433 1197
rect 1489 1195 1513 1197
rect 1569 1195 1593 1197
rect 1649 1195 1673 1197
rect 1729 1195 1753 1197
rect 1809 1195 1833 1197
rect 1889 1195 1913 1197
rect 1969 1195 1993 1197
rect 2049 1195 2073 1197
rect 2129 1196 2208 1197
rect 2129 1195 2282 1196
rect 1169 1143 1182 1195
rect 1426 1143 1433 1195
rect 1490 1143 1502 1195
rect 1746 1143 1753 1195
rect 1810 1143 1822 1195
rect 2066 1143 2073 1195
rect 2130 1143 2282 1195
rect 1169 1141 1193 1143
rect 1249 1141 1273 1143
rect 1329 1141 1353 1143
rect 1409 1141 1433 1143
rect 1489 1141 1513 1143
rect 1569 1141 1593 1143
rect 1649 1141 1673 1143
rect 1729 1141 1753 1143
rect 1809 1141 1833 1143
rect 1889 1141 1913 1143
rect 1969 1141 1993 1143
rect 2049 1141 2073 1143
rect 2129 1142 2282 1143
rect 2129 1141 2208 1142
rect 1113 1117 1169 1141
rect 0 1113 66 1114
rect 2216 1113 2282 1114
rect 0 1105 1085 1113
rect 0 1049 5 1105
rect 61 1049 1085 1105
rect 0 1025 7 1049
rect 59 1046 1085 1049
rect 1113 1049 1169 1061
rect 59 1025 66 1046
rect 0 969 5 1025
rect 61 969 66 1025
rect 1113 1037 1115 1049
rect 1167 1037 1169 1049
rect 1197 1105 2282 1113
rect 1197 1049 2221 1105
rect 2277 1049 2282 1105
rect 1197 1046 2223 1049
rect 94 990 1113 1018
rect 2216 1025 2223 1046
rect 2275 1025 2282 1049
rect 0 952 7 969
rect 59 962 66 969
rect 1169 990 2188 1018
rect 59 952 1085 962
rect 0 945 1085 952
rect 0 889 5 945
rect 61 934 1085 945
rect 1113 957 1115 981
rect 1167 957 1169 981
rect 2216 969 2221 1025
rect 2277 969 2282 1025
rect 2216 962 2223 969
rect 61 889 66 934
rect 1197 952 2223 962
rect 2275 952 2282 969
rect 1197 945 2282 952
rect 1197 934 2221 945
rect 0 888 7 889
rect 59 888 66 889
rect 0 876 66 888
rect 94 901 1113 906
rect 1169 901 2188 906
rect 94 878 1115 901
rect 0 865 7 876
rect 59 865 66 876
rect 0 809 5 865
rect 61 850 66 865
rect 1113 877 1115 878
rect 1167 878 2188 901
rect 2216 889 2221 934
rect 2277 889 2282 945
rect 2216 888 2223 889
rect 2275 888 2282 889
rect 1167 877 1169 878
rect 61 822 1085 850
rect 61 809 66 822
rect 0 785 7 809
rect 59 785 66 809
rect 2216 876 2282 888
rect 2216 865 2223 876
rect 2275 865 2282 876
rect 2216 850 2221 865
rect 1197 822 2221 850
rect 1113 805 1115 821
rect 1167 805 1169 821
rect 1113 797 1169 805
rect 0 729 5 785
rect 61 738 66 785
rect 94 766 1113 794
rect 2216 809 2221 822
rect 2277 809 2282 865
rect 1169 766 2188 794
rect 2216 785 2223 809
rect 2275 785 2282 809
rect 61 729 1085 738
rect 0 705 7 729
rect 59 710 1085 729
rect 1113 729 1169 741
rect 2216 738 2221 785
rect 1113 717 1115 729
rect 1167 717 1169 729
rect 59 705 66 710
rect 0 649 5 705
rect 61 649 66 705
rect 94 661 1113 682
rect 1197 729 2221 738
rect 2277 729 2282 785
rect 1197 710 2223 729
rect 2216 705 2223 710
rect 2275 705 2282 729
rect 1169 661 2188 682
rect 94 654 1115 661
rect 0 632 7 649
rect 59 632 66 649
rect 0 626 66 632
rect 1113 637 1115 654
rect 1167 654 2188 661
rect 1167 637 1169 654
rect 0 625 1085 626
rect 0 569 5 625
rect 61 598 1085 625
rect 2216 649 2221 705
rect 2277 649 2282 705
rect 2216 632 2223 649
rect 2275 632 2282 649
rect 2216 626 2282 632
rect 61 569 66 598
rect 1197 625 2282 626
rect 1197 598 2221 625
rect 1113 570 1115 581
rect 0 568 7 569
rect 59 568 66 569
rect 0 556 66 568
rect 0 545 7 556
rect 59 545 66 556
rect 0 489 5 545
rect 61 514 66 545
rect 94 557 1115 570
rect 1167 570 1169 581
rect 1167 557 2188 570
rect 94 542 1113 557
rect 1169 542 2188 557
rect 2216 569 2221 598
rect 2277 569 2282 625
rect 2216 568 2223 569
rect 2275 568 2282 569
rect 2216 556 2282 568
rect 2216 545 2223 556
rect 2275 545 2282 556
rect 61 489 1085 514
rect 0 465 7 489
rect 59 486 1085 489
rect 2216 514 2221 545
rect 59 465 66 486
rect 0 409 5 465
rect 61 409 66 465
rect 1113 485 1115 501
rect 1167 485 1169 501
rect 1197 489 2221 514
rect 2277 489 2282 545
rect 1197 486 2223 489
rect 1113 477 1169 485
rect 94 430 1113 458
rect 0 385 7 409
rect 59 402 66 409
rect 2216 465 2223 486
rect 2275 465 2282 489
rect 1169 430 2188 458
rect 1113 409 1169 421
rect 59 385 1085 402
rect 0 329 5 385
rect 61 374 1085 385
rect 1113 397 1115 409
rect 1167 397 1169 409
rect 2216 409 2221 465
rect 2277 409 2282 465
rect 2216 402 2223 409
rect 61 329 66 374
rect 1197 385 2223 402
rect 2275 385 2282 409
rect 1197 374 2221 385
rect 0 312 7 329
rect 59 312 66 329
rect 94 341 1113 346
rect 1169 341 2188 346
rect 94 318 1115 341
rect 0 305 66 312
rect 0 249 5 305
rect 61 290 66 305
rect 1113 317 1115 318
rect 1167 318 2188 341
rect 2216 329 2221 374
rect 2277 329 2282 385
rect 1167 317 1169 318
rect 61 262 1085 290
rect 2216 312 2223 329
rect 2275 312 2282 329
rect 2216 305 2282 312
rect 2216 290 2221 305
rect 61 249 66 262
rect 0 248 7 249
rect 59 248 66 249
rect 0 236 66 248
rect 0 225 7 236
rect 59 225 66 236
rect 1197 262 2221 290
rect 1113 237 1115 261
rect 1167 237 1169 261
rect 0 169 5 225
rect 61 178 66 225
rect 94 206 1113 234
rect 2216 249 2221 262
rect 2277 249 2282 305
rect 2216 248 2223 249
rect 2275 248 2282 249
rect 2216 236 2282 248
rect 1169 206 2188 234
rect 2216 225 2223 236
rect 2275 225 2282 236
rect 61 169 1085 178
rect 0 145 7 169
rect 59 150 1085 169
rect 1113 165 1115 181
rect 1167 165 1169 181
rect 2216 178 2221 225
rect 1113 153 1169 165
rect 59 145 66 150
rect 0 89 5 145
rect 61 89 66 145
rect 1113 122 1115 153
rect 94 101 1115 122
rect 1167 122 1169 153
rect 1197 169 2221 178
rect 2277 169 2282 225
rect 1197 150 2223 169
rect 2216 145 2223 150
rect 2275 145 2282 169
rect 1167 101 2188 122
rect 94 94 2188 101
rect 0 56 7 89
rect 59 66 66 89
rect 59 61 1086 66
rect 59 56 61 61
rect 117 59 141 61
rect 197 59 221 61
rect 277 59 301 61
rect 357 59 381 61
rect 437 59 461 61
rect 517 59 541 61
rect 597 59 621 61
rect 677 59 701 61
rect 757 59 781 61
rect 837 59 861 61
rect 917 59 941 61
rect 997 59 1021 61
rect 0 5 61 56
rect 140 7 141 59
rect 204 7 216 59
rect 277 7 280 59
rect 460 7 461 59
rect 524 7 536 59
rect 597 7 600 59
rect 780 7 781 59
rect 844 7 856 59
rect 917 7 920 59
rect 117 5 141 7
rect 197 5 221 7
rect 277 5 301 7
rect 357 5 381 7
rect 437 5 461 7
rect 517 5 541 7
rect 597 5 621 7
rect 677 5 701 7
rect 757 5 781 7
rect 837 5 861 7
rect 917 5 941 7
rect 997 5 1021 7
rect 1077 5 1086 61
rect 0 0 1086 5
rect 1114 0 1168 94
rect 2216 89 2221 145
rect 2277 89 2282 145
rect 2216 66 2223 89
rect 1196 61 2223 66
rect 1196 5 1205 61
rect 1261 59 1285 61
rect 1341 59 1365 61
rect 1421 59 1445 61
rect 1501 59 1525 61
rect 1581 59 1605 61
rect 1661 59 1685 61
rect 1741 59 1765 61
rect 1821 59 1845 61
rect 1901 59 1925 61
rect 1981 59 2005 61
rect 2061 59 2085 61
rect 2141 59 2165 61
rect 1362 7 1365 59
rect 1426 7 1438 59
rect 1501 7 1502 59
rect 1682 7 1685 59
rect 1746 7 1758 59
rect 1821 7 1822 59
rect 2002 7 2005 59
rect 2066 7 2078 59
rect 2141 7 2142 59
rect 2221 56 2223 61
rect 2275 56 2282 89
rect 1261 5 1285 7
rect 1341 5 1365 7
rect 1421 5 1445 7
rect 1501 5 1525 7
rect 1581 5 1605 7
rect 1661 5 1685 7
rect 1741 5 1765 7
rect 1821 5 1845 7
rect 1901 5 1925 7
rect 1981 5 2005 7
rect 2061 5 2085 7
rect 2141 5 2165 7
rect 2221 5 2282 56
rect 1196 0 2282 5
<< via2 >>
rect 61 2331 117 2333
rect 141 2331 197 2333
rect 221 2331 277 2333
rect 301 2331 357 2333
rect 381 2331 437 2333
rect 461 2331 517 2333
rect 541 2331 597 2333
rect 621 2331 677 2333
rect 701 2331 757 2333
rect 781 2331 837 2333
rect 861 2331 917 2333
rect 941 2331 997 2333
rect 1021 2331 1077 2333
rect 61 2279 88 2331
rect 88 2279 117 2331
rect 141 2279 152 2331
rect 152 2279 197 2331
rect 221 2279 268 2331
rect 268 2279 277 2331
rect 301 2279 332 2331
rect 332 2279 344 2331
rect 344 2279 357 2331
rect 381 2279 396 2331
rect 396 2279 408 2331
rect 408 2279 437 2331
rect 461 2279 472 2331
rect 472 2279 517 2331
rect 541 2279 588 2331
rect 588 2279 597 2331
rect 621 2279 652 2331
rect 652 2279 664 2331
rect 664 2279 677 2331
rect 701 2279 716 2331
rect 716 2279 728 2331
rect 728 2279 757 2331
rect 781 2279 792 2331
rect 792 2279 837 2331
rect 861 2279 908 2331
rect 908 2279 917 2331
rect 941 2279 972 2331
rect 972 2279 984 2331
rect 984 2279 997 2331
rect 1021 2279 1036 2331
rect 1036 2279 1077 2331
rect 61 2277 117 2279
rect 141 2277 197 2279
rect 221 2277 277 2279
rect 301 2277 357 2279
rect 381 2277 437 2279
rect 461 2277 517 2279
rect 541 2277 597 2279
rect 621 2277 677 2279
rect 701 2277 757 2279
rect 781 2277 837 2279
rect 861 2277 917 2279
rect 941 2277 997 2279
rect 1021 2277 1077 2279
rect 5 2230 7 2249
rect 7 2230 59 2249
rect 59 2230 61 2249
rect 5 2218 61 2230
rect 5 2193 7 2218
rect 7 2193 59 2218
rect 59 2193 61 2218
rect 1205 2331 1261 2333
rect 1285 2331 1341 2333
rect 1365 2331 1421 2333
rect 1445 2331 1501 2333
rect 1525 2331 1581 2333
rect 1605 2331 1661 2333
rect 1685 2331 1741 2333
rect 1765 2331 1821 2333
rect 1845 2331 1901 2333
rect 1925 2331 1981 2333
rect 2005 2331 2061 2333
rect 2085 2331 2141 2333
rect 2165 2331 2221 2333
rect 1205 2279 1246 2331
rect 1246 2279 1261 2331
rect 1285 2279 1298 2331
rect 1298 2279 1310 2331
rect 1310 2279 1341 2331
rect 1365 2279 1374 2331
rect 1374 2279 1421 2331
rect 1445 2279 1490 2331
rect 1490 2279 1501 2331
rect 1525 2279 1554 2331
rect 1554 2279 1566 2331
rect 1566 2279 1581 2331
rect 1605 2279 1618 2331
rect 1618 2279 1630 2331
rect 1630 2279 1661 2331
rect 1685 2279 1694 2331
rect 1694 2279 1741 2331
rect 1765 2279 1810 2331
rect 1810 2279 1821 2331
rect 1845 2279 1874 2331
rect 1874 2279 1886 2331
rect 1886 2279 1901 2331
rect 1925 2279 1938 2331
rect 1938 2279 1950 2331
rect 1950 2279 1981 2331
rect 2005 2279 2014 2331
rect 2014 2279 2061 2331
rect 2085 2279 2130 2331
rect 2130 2279 2141 2331
rect 2165 2279 2194 2331
rect 2194 2279 2221 2331
rect 1205 2277 1261 2279
rect 1285 2277 1341 2279
rect 1365 2277 1421 2279
rect 1445 2277 1501 2279
rect 1525 2277 1581 2279
rect 1605 2277 1661 2279
rect 1685 2277 1741 2279
rect 1765 2277 1821 2279
rect 1845 2277 1901 2279
rect 1925 2277 1981 2279
rect 2005 2277 2061 2279
rect 2085 2277 2141 2279
rect 2165 2277 2221 2279
rect 5 2166 7 2169
rect 7 2166 59 2169
rect 59 2166 61 2169
rect 5 2154 61 2166
rect 2221 2230 2223 2249
rect 2223 2230 2275 2249
rect 2275 2230 2277 2249
rect 2221 2218 2277 2230
rect 2221 2193 2223 2218
rect 2223 2193 2275 2218
rect 2275 2193 2277 2218
rect 5 2113 7 2154
rect 7 2113 59 2154
rect 59 2113 61 2154
rect 2221 2166 2223 2169
rect 2223 2166 2275 2169
rect 2275 2166 2277 2169
rect 1113 2121 1115 2157
rect 1115 2121 1167 2157
rect 1167 2121 1169 2157
rect 1113 2109 1169 2121
rect 5 2038 7 2089
rect 7 2038 59 2089
rect 59 2038 61 2089
rect 1113 2101 1115 2109
rect 1115 2101 1167 2109
rect 1167 2101 1169 2109
rect 2221 2154 2277 2166
rect 2221 2113 2223 2154
rect 2223 2113 2275 2154
rect 2275 2113 2277 2154
rect 1113 2057 1115 2077
rect 1115 2057 1167 2077
rect 1167 2057 1169 2077
rect 5 2033 61 2038
rect 1113 2045 1169 2057
rect 1113 2021 1115 2045
rect 1115 2021 1167 2045
rect 1167 2021 1169 2045
rect 5 1974 7 2009
rect 7 1974 59 2009
rect 59 1974 61 2009
rect 5 1962 61 1974
rect 2221 2038 2223 2089
rect 2223 2038 2275 2089
rect 2275 2038 2277 2089
rect 2221 2033 2277 2038
rect 1113 1993 1115 1997
rect 1115 1993 1167 1997
rect 1167 1993 1169 1997
rect 1113 1981 1169 1993
rect 5 1953 7 1962
rect 7 1953 59 1962
rect 59 1953 61 1962
rect 1113 1941 1115 1981
rect 1115 1941 1167 1981
rect 1167 1941 1169 1981
rect 2221 1974 2223 2009
rect 2223 1974 2275 2009
rect 2275 1974 2277 2009
rect 5 1910 7 1929
rect 7 1910 59 1929
rect 59 1910 61 1929
rect 5 1898 61 1910
rect 5 1873 7 1898
rect 7 1873 59 1898
rect 59 1873 61 1898
rect 2221 1962 2277 1974
rect 2221 1953 2223 1962
rect 2223 1953 2275 1962
rect 2275 1953 2277 1962
rect 1113 1865 1115 1917
rect 1115 1865 1167 1917
rect 1167 1865 1169 1917
rect 1113 1861 1169 1865
rect 5 1846 7 1849
rect 7 1846 59 1849
rect 59 1846 61 1849
rect 5 1834 61 1846
rect 5 1793 7 1834
rect 7 1793 59 1834
rect 59 1793 61 1834
rect 2221 1910 2223 1929
rect 2223 1910 2275 1929
rect 2275 1910 2277 1929
rect 2221 1898 2277 1910
rect 2221 1873 2223 1898
rect 2223 1873 2275 1898
rect 2275 1873 2277 1898
rect 1113 1801 1115 1837
rect 1115 1801 1167 1837
rect 1167 1801 1169 1837
rect 2221 1846 2223 1849
rect 2223 1846 2275 1849
rect 2275 1846 2277 1849
rect 2221 1834 2277 1846
rect 5 1718 7 1769
rect 7 1718 59 1769
rect 59 1718 61 1769
rect 1113 1789 1169 1801
rect 1113 1781 1115 1789
rect 1115 1781 1167 1789
rect 1167 1781 1169 1789
rect 2221 1793 2223 1834
rect 2223 1793 2275 1834
rect 2275 1793 2277 1834
rect 5 1713 61 1718
rect 1113 1737 1115 1757
rect 1115 1737 1167 1757
rect 1167 1737 1169 1757
rect 1113 1725 1169 1737
rect 5 1654 7 1689
rect 7 1654 59 1689
rect 59 1654 61 1689
rect 5 1642 61 1654
rect 5 1633 7 1642
rect 7 1633 59 1642
rect 59 1633 61 1642
rect 1113 1701 1115 1725
rect 1115 1701 1167 1725
rect 1167 1701 1169 1725
rect 2221 1718 2223 1769
rect 2223 1718 2275 1769
rect 2275 1718 2277 1769
rect 2221 1713 2277 1718
rect 1113 1673 1115 1677
rect 1115 1673 1167 1677
rect 1167 1673 1169 1677
rect 1113 1661 1169 1673
rect 5 1590 7 1609
rect 7 1590 59 1609
rect 59 1590 61 1609
rect 1113 1621 1115 1661
rect 1115 1621 1167 1661
rect 1167 1621 1169 1661
rect 2221 1654 2223 1689
rect 2223 1654 2275 1689
rect 2275 1654 2277 1689
rect 2221 1642 2277 1654
rect 2221 1633 2223 1642
rect 2223 1633 2275 1642
rect 2275 1633 2277 1642
rect 5 1578 61 1590
rect 5 1553 7 1578
rect 7 1553 59 1578
rect 59 1553 61 1578
rect 1113 1545 1115 1597
rect 1115 1545 1167 1597
rect 1167 1545 1169 1597
rect 5 1526 7 1529
rect 7 1526 59 1529
rect 59 1526 61 1529
rect 5 1514 61 1526
rect 1113 1541 1169 1545
rect 2221 1590 2223 1609
rect 2223 1590 2275 1609
rect 2275 1590 2277 1609
rect 2221 1578 2277 1590
rect 2221 1553 2223 1578
rect 2223 1553 2275 1578
rect 2275 1553 2277 1578
rect 5 1473 7 1514
rect 7 1473 59 1514
rect 59 1473 61 1514
rect 1113 1481 1115 1517
rect 1115 1481 1167 1517
rect 1167 1481 1169 1517
rect 2221 1526 2223 1529
rect 2223 1526 2275 1529
rect 2275 1526 2277 1529
rect 2221 1514 2277 1526
rect 1113 1469 1169 1481
rect 1113 1461 1115 1469
rect 1115 1461 1167 1469
rect 1167 1461 1169 1469
rect 5 1398 7 1449
rect 7 1398 59 1449
rect 59 1398 61 1449
rect 2221 1473 2223 1514
rect 2223 1473 2275 1514
rect 2275 1473 2277 1514
rect 1113 1417 1115 1437
rect 1115 1417 1167 1437
rect 1167 1417 1169 1437
rect 1113 1405 1169 1417
rect 5 1393 61 1398
rect 1113 1381 1115 1405
rect 1115 1381 1167 1405
rect 1167 1381 1169 1405
rect 5 1334 7 1369
rect 7 1334 59 1369
rect 59 1334 61 1369
rect 5 1322 61 1334
rect 5 1313 7 1322
rect 7 1313 59 1322
rect 59 1313 61 1322
rect 2221 1398 2223 1449
rect 2223 1398 2275 1449
rect 2275 1398 2277 1449
rect 2221 1393 2277 1398
rect 1113 1353 1115 1357
rect 1115 1353 1167 1357
rect 1167 1353 1169 1357
rect 1113 1341 1169 1353
rect 1113 1301 1115 1341
rect 1115 1301 1167 1341
rect 1167 1301 1169 1341
rect 5 1270 7 1289
rect 7 1270 59 1289
rect 59 1270 61 1289
rect 5 1233 61 1270
rect 2221 1334 2223 1369
rect 2223 1334 2275 1369
rect 2275 1334 2277 1369
rect 2221 1322 2277 1334
rect 2221 1313 2223 1322
rect 2223 1313 2275 1322
rect 2275 1313 2277 1322
rect 1113 1225 1115 1277
rect 1115 1225 1167 1277
rect 1167 1225 1169 1277
rect 2221 1270 2223 1289
rect 2223 1270 2275 1289
rect 2275 1270 2277 1289
rect 2221 1233 2277 1270
rect 1113 1221 1169 1225
rect 153 1195 209 1197
rect 233 1195 289 1197
rect 313 1195 369 1197
rect 393 1195 449 1197
rect 473 1195 529 1197
rect 553 1195 609 1197
rect 633 1195 689 1197
rect 713 1195 769 1197
rect 793 1195 849 1197
rect 873 1195 929 1197
rect 953 1195 1009 1197
rect 1033 1195 1089 1197
rect 153 1143 204 1195
rect 204 1143 209 1195
rect 233 1143 268 1195
rect 268 1143 280 1195
rect 280 1143 289 1195
rect 313 1143 332 1195
rect 332 1143 344 1195
rect 344 1143 369 1195
rect 393 1143 396 1195
rect 396 1143 408 1195
rect 408 1143 449 1195
rect 473 1143 524 1195
rect 524 1143 529 1195
rect 553 1143 588 1195
rect 588 1143 600 1195
rect 600 1143 609 1195
rect 633 1143 652 1195
rect 652 1143 664 1195
rect 664 1143 689 1195
rect 713 1143 716 1195
rect 716 1143 728 1195
rect 728 1143 769 1195
rect 793 1143 844 1195
rect 844 1143 849 1195
rect 873 1143 908 1195
rect 908 1143 920 1195
rect 920 1143 929 1195
rect 953 1143 972 1195
rect 972 1143 984 1195
rect 984 1143 1009 1195
rect 1033 1143 1036 1195
rect 1036 1143 1048 1195
rect 1048 1143 1089 1195
rect 153 1141 209 1143
rect 233 1141 289 1143
rect 313 1141 369 1143
rect 393 1141 449 1143
rect 473 1141 529 1143
rect 553 1141 609 1143
rect 633 1141 689 1143
rect 713 1141 769 1143
rect 793 1141 849 1143
rect 873 1141 929 1143
rect 953 1141 1009 1143
rect 1033 1141 1089 1143
rect 1113 1141 1169 1197
rect 1193 1195 1249 1197
rect 1273 1195 1329 1197
rect 1353 1195 1409 1197
rect 1433 1195 1489 1197
rect 1513 1195 1569 1197
rect 1593 1195 1649 1197
rect 1673 1195 1729 1197
rect 1753 1195 1809 1197
rect 1833 1195 1889 1197
rect 1913 1195 1969 1197
rect 1993 1195 2049 1197
rect 2073 1195 2129 1197
rect 1193 1143 1234 1195
rect 1234 1143 1246 1195
rect 1246 1143 1249 1195
rect 1273 1143 1298 1195
rect 1298 1143 1310 1195
rect 1310 1143 1329 1195
rect 1353 1143 1362 1195
rect 1362 1143 1374 1195
rect 1374 1143 1409 1195
rect 1433 1143 1438 1195
rect 1438 1143 1489 1195
rect 1513 1143 1554 1195
rect 1554 1143 1566 1195
rect 1566 1143 1569 1195
rect 1593 1143 1618 1195
rect 1618 1143 1630 1195
rect 1630 1143 1649 1195
rect 1673 1143 1682 1195
rect 1682 1143 1694 1195
rect 1694 1143 1729 1195
rect 1753 1143 1758 1195
rect 1758 1143 1809 1195
rect 1833 1143 1874 1195
rect 1874 1143 1886 1195
rect 1886 1143 1889 1195
rect 1913 1143 1938 1195
rect 1938 1143 1950 1195
rect 1950 1143 1969 1195
rect 1993 1143 2002 1195
rect 2002 1143 2014 1195
rect 2014 1143 2049 1195
rect 2073 1143 2078 1195
rect 2078 1143 2129 1195
rect 1193 1141 1249 1143
rect 1273 1141 1329 1143
rect 1353 1141 1409 1143
rect 1433 1141 1489 1143
rect 1513 1141 1569 1143
rect 1593 1141 1649 1143
rect 1673 1141 1729 1143
rect 1753 1141 1809 1143
rect 1833 1141 1889 1143
rect 1913 1141 1969 1143
rect 1993 1141 2049 1143
rect 2073 1141 2129 1143
rect 1113 1113 1169 1117
rect 5 1068 61 1105
rect 5 1049 7 1068
rect 7 1049 59 1068
rect 59 1049 61 1068
rect 1113 1061 1115 1113
rect 1115 1061 1167 1113
rect 1167 1061 1169 1113
rect 5 1016 7 1025
rect 7 1016 59 1025
rect 59 1016 61 1025
rect 5 1004 61 1016
rect 5 969 7 1004
rect 7 969 59 1004
rect 59 969 61 1004
rect 2221 1068 2277 1105
rect 2221 1049 2223 1068
rect 2223 1049 2275 1068
rect 2275 1049 2277 1068
rect 1113 997 1115 1037
rect 1115 997 1167 1037
rect 1167 997 1169 1037
rect 1113 985 1169 997
rect 1113 981 1115 985
rect 1115 981 1167 985
rect 1167 981 1169 985
rect 5 940 61 945
rect 5 889 7 940
rect 7 889 59 940
rect 59 889 61 940
rect 2221 1016 2223 1025
rect 2223 1016 2275 1025
rect 2275 1016 2277 1025
rect 2221 1004 2277 1016
rect 2221 969 2223 1004
rect 2223 969 2275 1004
rect 2275 969 2277 1004
rect 1113 933 1115 957
rect 1115 933 1167 957
rect 1167 933 1169 957
rect 2221 940 2277 945
rect 1113 921 1169 933
rect 1113 901 1115 921
rect 1115 901 1167 921
rect 1167 901 1169 921
rect 5 824 7 865
rect 7 824 59 865
rect 59 824 61 865
rect 2221 889 2223 940
rect 2223 889 2275 940
rect 2275 889 2277 940
rect 1113 869 1115 877
rect 1115 869 1167 877
rect 1167 869 1169 877
rect 1113 857 1169 869
rect 5 812 61 824
rect 5 809 7 812
rect 7 809 59 812
rect 59 809 61 812
rect 1113 821 1115 857
rect 1115 821 1167 857
rect 1167 821 1169 857
rect 2221 824 2223 865
rect 2223 824 2275 865
rect 2275 824 2277 865
rect 5 760 7 785
rect 7 760 59 785
rect 59 760 61 785
rect 5 748 61 760
rect 5 729 7 748
rect 7 729 59 748
rect 59 729 61 748
rect 1113 793 1169 797
rect 2221 812 2277 824
rect 2221 809 2223 812
rect 2223 809 2275 812
rect 2275 809 2277 812
rect 1113 741 1115 793
rect 1115 741 1167 793
rect 1167 741 1169 793
rect 2221 760 2223 785
rect 2223 760 2275 785
rect 2275 760 2277 785
rect 2221 748 2277 760
rect 5 696 7 705
rect 7 696 59 705
rect 59 696 61 705
rect 5 684 61 696
rect 5 649 7 684
rect 7 649 59 684
rect 59 649 61 684
rect 1113 677 1115 717
rect 1115 677 1167 717
rect 1167 677 1169 717
rect 2221 729 2223 748
rect 2223 729 2275 748
rect 2275 729 2277 748
rect 1113 665 1169 677
rect 1113 661 1115 665
rect 1115 661 1167 665
rect 1167 661 1169 665
rect 5 620 61 625
rect 5 569 7 620
rect 7 569 59 620
rect 59 569 61 620
rect 1113 613 1115 637
rect 1115 613 1167 637
rect 1167 613 1169 637
rect 2221 696 2223 705
rect 2223 696 2275 705
rect 2275 696 2277 705
rect 2221 684 2277 696
rect 2221 649 2223 684
rect 2223 649 2275 684
rect 2275 649 2277 684
rect 1113 601 1169 613
rect 1113 581 1115 601
rect 1115 581 1167 601
rect 1167 581 1169 601
rect 2221 620 2277 625
rect 5 504 7 545
rect 7 504 59 545
rect 59 504 61 545
rect 1113 549 1115 557
rect 1115 549 1167 557
rect 1167 549 1169 557
rect 1113 537 1169 549
rect 2221 569 2223 620
rect 2223 569 2275 620
rect 2275 569 2277 620
rect 5 492 61 504
rect 5 489 7 492
rect 7 489 59 492
rect 59 489 61 492
rect 1113 501 1115 537
rect 1115 501 1167 537
rect 1167 501 1169 537
rect 5 440 7 465
rect 7 440 59 465
rect 59 440 61 465
rect 5 428 61 440
rect 5 409 7 428
rect 7 409 59 428
rect 59 409 61 428
rect 2221 504 2223 545
rect 2223 504 2275 545
rect 2275 504 2277 545
rect 2221 492 2277 504
rect 2221 489 2223 492
rect 2223 489 2275 492
rect 2275 489 2277 492
rect 1113 473 1169 477
rect 1113 421 1115 473
rect 1115 421 1167 473
rect 1167 421 1169 473
rect 5 376 7 385
rect 7 376 59 385
rect 59 376 61 385
rect 5 364 61 376
rect 2221 440 2223 465
rect 2223 440 2275 465
rect 2275 440 2277 465
rect 2221 428 2277 440
rect 2221 409 2223 428
rect 2223 409 2275 428
rect 2275 409 2277 428
rect 5 329 7 364
rect 7 329 59 364
rect 59 329 61 364
rect 1113 357 1115 397
rect 1115 357 1167 397
rect 1167 357 1169 397
rect 2221 376 2223 385
rect 2223 376 2275 385
rect 2275 376 2277 385
rect 1113 345 1169 357
rect 1113 341 1115 345
rect 1115 341 1167 345
rect 1167 341 1169 345
rect 5 300 61 305
rect 5 249 7 300
rect 7 249 59 300
rect 59 249 61 300
rect 2221 364 2277 376
rect 2221 329 2223 364
rect 2223 329 2275 364
rect 2275 329 2277 364
rect 1113 293 1115 317
rect 1115 293 1167 317
rect 1167 293 1169 317
rect 1113 281 1169 293
rect 2221 300 2277 305
rect 1113 261 1115 281
rect 1115 261 1167 281
rect 1167 261 1169 281
rect 5 184 7 225
rect 7 184 59 225
rect 59 184 61 225
rect 5 172 61 184
rect 1113 229 1115 237
rect 1115 229 1167 237
rect 1167 229 1169 237
rect 2221 249 2223 300
rect 2223 249 2275 300
rect 2275 249 2277 300
rect 1113 217 1169 229
rect 1113 181 1115 217
rect 1115 181 1167 217
rect 1167 181 1169 217
rect 5 169 7 172
rect 7 169 59 172
rect 59 169 61 172
rect 2221 184 2223 225
rect 2223 184 2275 225
rect 2275 184 2277 225
rect 5 120 7 145
rect 7 120 59 145
rect 59 120 61 145
rect 5 108 61 120
rect 5 89 7 108
rect 7 89 59 108
rect 59 89 61 108
rect 2221 172 2277 184
rect 2221 169 2223 172
rect 2223 169 2275 172
rect 2275 169 2277 172
rect 61 59 117 61
rect 141 59 197 61
rect 221 59 277 61
rect 301 59 357 61
rect 381 59 437 61
rect 461 59 517 61
rect 541 59 597 61
rect 621 59 677 61
rect 701 59 757 61
rect 781 59 837 61
rect 861 59 917 61
rect 941 59 997 61
rect 1021 59 1077 61
rect 61 7 88 59
rect 88 7 117 59
rect 141 7 152 59
rect 152 7 197 59
rect 221 7 268 59
rect 268 7 277 59
rect 301 7 332 59
rect 332 7 344 59
rect 344 7 357 59
rect 381 7 396 59
rect 396 7 408 59
rect 408 7 437 59
rect 461 7 472 59
rect 472 7 517 59
rect 541 7 588 59
rect 588 7 597 59
rect 621 7 652 59
rect 652 7 664 59
rect 664 7 677 59
rect 701 7 716 59
rect 716 7 728 59
rect 728 7 757 59
rect 781 7 792 59
rect 792 7 837 59
rect 861 7 908 59
rect 908 7 917 59
rect 941 7 972 59
rect 972 7 984 59
rect 984 7 997 59
rect 1021 7 1036 59
rect 1036 7 1077 59
rect 61 5 117 7
rect 141 5 197 7
rect 221 5 277 7
rect 301 5 357 7
rect 381 5 437 7
rect 461 5 517 7
rect 541 5 597 7
rect 621 5 677 7
rect 701 5 757 7
rect 781 5 837 7
rect 861 5 917 7
rect 941 5 997 7
rect 1021 5 1077 7
rect 2221 120 2223 145
rect 2223 120 2275 145
rect 2275 120 2277 145
rect 2221 108 2277 120
rect 2221 89 2223 108
rect 2223 89 2275 108
rect 2275 89 2277 108
rect 1205 59 1261 61
rect 1285 59 1341 61
rect 1365 59 1421 61
rect 1445 59 1501 61
rect 1525 59 1581 61
rect 1605 59 1661 61
rect 1685 59 1741 61
rect 1765 59 1821 61
rect 1845 59 1901 61
rect 1925 59 1981 61
rect 2005 59 2061 61
rect 2085 59 2141 61
rect 2165 59 2221 61
rect 1205 7 1246 59
rect 1246 7 1261 59
rect 1285 7 1298 59
rect 1298 7 1310 59
rect 1310 7 1341 59
rect 1365 7 1374 59
rect 1374 7 1421 59
rect 1445 7 1490 59
rect 1490 7 1501 59
rect 1525 7 1554 59
rect 1554 7 1566 59
rect 1566 7 1581 59
rect 1605 7 1618 59
rect 1618 7 1630 59
rect 1630 7 1661 59
rect 1685 7 1694 59
rect 1694 7 1741 59
rect 1765 7 1810 59
rect 1810 7 1821 59
rect 1845 7 1874 59
rect 1874 7 1886 59
rect 1886 7 1901 59
rect 1925 7 1938 59
rect 1938 7 1950 59
rect 1950 7 1981 59
rect 2005 7 2014 59
rect 2014 7 2061 59
rect 2085 7 2130 59
rect 2130 7 2141 59
rect 2165 7 2194 59
rect 2194 7 2221 59
rect 1205 5 1261 7
rect 1285 5 1341 7
rect 1365 5 1421 7
rect 1445 5 1501 7
rect 1525 5 1581 7
rect 1605 5 1661 7
rect 1685 5 1741 7
rect 1765 5 1821 7
rect 1845 5 1901 7
rect 1925 5 1981 7
rect 2005 5 2061 7
rect 2085 5 2141 7
rect 2165 5 2221 7
<< metal3 >>
rect 0 2337 2282 2338
rect 0 2333 85 2337
rect 149 2333 165 2337
rect 229 2333 245 2337
rect 309 2333 325 2337
rect 389 2333 405 2337
rect 469 2333 485 2337
rect 549 2333 565 2337
rect 629 2333 645 2337
rect 709 2333 725 2337
rect 789 2333 805 2337
rect 869 2333 885 2337
rect 949 2333 965 2337
rect 1029 2333 1045 2337
rect 1109 2333 1229 2337
rect 1293 2333 1309 2337
rect 1373 2333 1389 2337
rect 1453 2333 1469 2337
rect 1533 2333 1549 2337
rect 1613 2333 1629 2337
rect 1693 2333 1709 2337
rect 1773 2333 1789 2337
rect 1853 2333 1869 2337
rect 1933 2333 1949 2337
rect 2013 2333 2029 2337
rect 2093 2333 2109 2337
rect 2173 2333 2282 2337
rect 0 2277 61 2333
rect 1109 2277 1205 2333
rect 2221 2277 2282 2333
rect 0 2273 85 2277
rect 149 2273 165 2277
rect 229 2273 245 2277
rect 309 2273 325 2277
rect 389 2273 405 2277
rect 469 2273 485 2277
rect 549 2273 565 2277
rect 629 2273 645 2277
rect 709 2273 725 2277
rect 789 2273 805 2277
rect 869 2273 885 2277
rect 949 2273 965 2277
rect 1029 2273 1045 2277
rect 1109 2273 1229 2277
rect 1293 2273 1309 2277
rect 1373 2273 1389 2277
rect 1453 2273 1469 2277
rect 1533 2273 1549 2277
rect 1613 2273 1629 2277
rect 1693 2273 1709 2277
rect 1773 2273 1789 2277
rect 1853 2273 1869 2277
rect 1933 2273 1949 2277
rect 2013 2273 2029 2277
rect 2093 2273 2109 2277
rect 2173 2273 2282 2277
rect 0 2272 2282 2273
rect 0 2249 66 2272
rect 0 2225 5 2249
rect 61 2225 66 2249
rect 0 2161 1 2225
rect 65 2161 66 2225
rect 0 2145 5 2161
rect 61 2145 66 2161
rect 0 2081 1 2145
rect 65 2081 66 2145
rect 0 2065 5 2081
rect 61 2065 66 2081
rect 0 2001 1 2065
rect 65 2001 66 2065
rect 0 1985 5 2001
rect 61 1985 66 2001
rect 0 1921 1 1985
rect 65 1921 66 1985
rect 0 1905 5 1921
rect 61 1905 66 1921
rect 0 1841 1 1905
rect 65 1841 66 1905
rect 0 1825 5 1841
rect 61 1825 66 1841
rect 0 1761 1 1825
rect 65 1761 66 1825
rect 0 1745 5 1761
rect 61 1745 66 1761
rect 0 1681 1 1745
rect 65 1681 66 1745
rect 0 1665 5 1681
rect 61 1665 66 1681
rect 0 1601 1 1665
rect 65 1601 66 1665
rect 0 1585 5 1601
rect 61 1585 66 1601
rect 0 1521 1 1585
rect 65 1521 66 1585
rect 0 1505 5 1521
rect 61 1505 66 1521
rect 0 1441 1 1505
rect 65 1441 66 1505
rect 0 1425 5 1441
rect 61 1425 66 1441
rect 0 1361 1 1425
rect 65 1361 66 1425
rect 0 1345 5 1361
rect 61 1345 66 1361
rect 0 1281 1 1345
rect 65 1281 66 1345
rect 0 1265 5 1281
rect 61 1265 66 1281
rect 0 1201 1 1265
rect 65 1201 66 1265
rect 0 1105 66 1201
rect 0 1081 5 1105
rect 61 1081 66 1105
rect 0 1017 1 1081
rect 65 1017 66 1081
rect 0 1001 5 1017
rect 61 1001 66 1017
rect 0 937 1 1001
rect 65 937 66 1001
rect 0 921 5 937
rect 61 921 66 937
rect 0 857 1 921
rect 65 857 66 921
rect 0 841 5 857
rect 61 841 66 857
rect 0 777 1 841
rect 65 777 66 841
rect 0 761 5 777
rect 61 761 66 777
rect 0 697 1 761
rect 65 697 66 761
rect 0 681 5 697
rect 61 681 66 697
rect 0 617 1 681
rect 65 617 66 681
rect 0 601 5 617
rect 61 601 66 617
rect 0 537 1 601
rect 65 537 66 601
rect 0 521 5 537
rect 61 521 66 537
rect 0 457 1 521
rect 65 457 66 521
rect 0 441 5 457
rect 61 441 66 457
rect 0 377 1 441
rect 65 377 66 441
rect 0 361 5 377
rect 61 361 66 377
rect 0 297 1 361
rect 65 297 66 361
rect 0 281 5 297
rect 61 281 66 297
rect 0 217 1 281
rect 65 217 66 281
rect 0 201 5 217
rect 61 201 66 217
rect 0 137 1 201
rect 65 137 66 201
rect 0 121 5 137
rect 61 121 66 137
rect 126 1202 186 2212
rect 246 1262 306 2272
rect 366 1202 426 2212
rect 486 1262 546 2272
rect 606 1202 666 2212
rect 726 1262 786 2272
rect 846 1202 906 2212
rect 966 1262 1048 2272
rect 1108 2161 1174 2212
rect 1108 2097 1109 2161
rect 1173 2097 1174 2161
rect 1108 2081 1174 2097
rect 1108 2017 1109 2081
rect 1173 2017 1174 2081
rect 1108 2001 1174 2017
rect 1108 1937 1109 2001
rect 1173 1937 1174 2001
rect 1108 1921 1174 1937
rect 1108 1857 1109 1921
rect 1173 1857 1174 1921
rect 1108 1841 1174 1857
rect 1108 1777 1109 1841
rect 1173 1777 1174 1841
rect 1108 1761 1174 1777
rect 1108 1697 1109 1761
rect 1173 1697 1174 1761
rect 1108 1681 1174 1697
rect 1108 1617 1109 1681
rect 1173 1617 1174 1681
rect 1108 1601 1174 1617
rect 1108 1537 1109 1601
rect 1173 1537 1174 1601
rect 1108 1521 1174 1537
rect 1108 1457 1109 1521
rect 1173 1457 1174 1521
rect 1108 1441 1174 1457
rect 1108 1377 1109 1441
rect 1173 1377 1174 1441
rect 1108 1361 1174 1377
rect 1108 1297 1109 1361
rect 1173 1297 1174 1361
rect 1108 1281 1174 1297
rect 1108 1217 1109 1281
rect 1173 1217 1174 1281
rect 1234 1262 1316 2272
rect 1108 1202 1174 1217
rect 1376 1202 1436 2212
rect 1496 1262 1556 2272
rect 1616 1202 1676 2212
rect 1736 1262 1796 2272
rect 1856 1202 1916 2212
rect 1976 1262 2036 2272
rect 2216 2249 2282 2272
rect 2216 2225 2221 2249
rect 2277 2225 2282 2249
rect 2096 1202 2156 2212
rect 126 1201 2156 1202
rect 126 1137 149 1201
rect 213 1137 229 1201
rect 293 1137 309 1201
rect 373 1137 389 1201
rect 453 1137 469 1201
rect 533 1137 549 1201
rect 613 1137 629 1201
rect 693 1137 709 1201
rect 773 1137 789 1201
rect 853 1137 869 1201
rect 933 1137 949 1201
rect 1013 1137 1029 1201
rect 1093 1137 1109 1201
rect 1173 1137 1189 1201
rect 1253 1137 1269 1201
rect 1333 1137 1349 1201
rect 1413 1137 1429 1201
rect 1493 1137 1509 1201
rect 1573 1137 1589 1201
rect 1653 1137 1669 1201
rect 1733 1137 1749 1201
rect 1813 1137 1829 1201
rect 1893 1137 1909 1201
rect 1973 1137 1989 1201
rect 2053 1137 2069 1201
rect 2133 1137 2156 1201
rect 126 1136 2156 1137
rect 126 126 186 1136
rect 0 57 1 121
rect 65 66 66 121
rect 246 66 306 1076
rect 366 126 426 1136
rect 486 66 546 1076
rect 606 126 666 1136
rect 726 66 786 1076
rect 846 126 906 1136
rect 1108 1121 1174 1136
rect 966 66 1048 1076
rect 1108 1057 1109 1121
rect 1173 1057 1174 1121
rect 1108 1041 1174 1057
rect 1108 977 1109 1041
rect 1173 977 1174 1041
rect 1108 961 1174 977
rect 1108 897 1109 961
rect 1173 897 1174 961
rect 1108 881 1174 897
rect 1108 817 1109 881
rect 1173 817 1174 881
rect 1108 801 1174 817
rect 1108 737 1109 801
rect 1173 737 1174 801
rect 1108 721 1174 737
rect 1108 657 1109 721
rect 1173 657 1174 721
rect 1108 641 1174 657
rect 1108 577 1109 641
rect 1173 577 1174 641
rect 1108 561 1174 577
rect 1108 497 1109 561
rect 1173 497 1174 561
rect 1108 481 1174 497
rect 1108 417 1109 481
rect 1173 417 1174 481
rect 1108 401 1174 417
rect 1108 337 1109 401
rect 1173 337 1174 401
rect 1108 321 1174 337
rect 1108 257 1109 321
rect 1173 257 1174 321
rect 1108 241 1174 257
rect 1108 177 1109 241
rect 1173 177 1174 241
rect 1108 126 1174 177
rect 1234 66 1316 1076
rect 1376 126 1436 1136
rect 1496 66 1556 1076
rect 1616 126 1676 1136
rect 1736 66 1796 1076
rect 1856 126 1916 1136
rect 1976 66 2036 1076
rect 2096 126 2156 1136
rect 2216 2161 2217 2225
rect 2281 2161 2282 2225
rect 2216 2145 2221 2161
rect 2277 2145 2282 2161
rect 2216 2081 2217 2145
rect 2281 2081 2282 2145
rect 2216 2065 2221 2081
rect 2277 2065 2282 2081
rect 2216 2001 2217 2065
rect 2281 2001 2282 2065
rect 2216 1985 2221 2001
rect 2277 1985 2282 2001
rect 2216 1921 2217 1985
rect 2281 1921 2282 1985
rect 2216 1905 2221 1921
rect 2277 1905 2282 1921
rect 2216 1841 2217 1905
rect 2281 1841 2282 1905
rect 2216 1825 2221 1841
rect 2277 1825 2282 1841
rect 2216 1761 2217 1825
rect 2281 1761 2282 1825
rect 2216 1745 2221 1761
rect 2277 1745 2282 1761
rect 2216 1681 2217 1745
rect 2281 1681 2282 1745
rect 2216 1665 2221 1681
rect 2277 1665 2282 1681
rect 2216 1601 2217 1665
rect 2281 1601 2282 1665
rect 2216 1585 2221 1601
rect 2277 1585 2282 1601
rect 2216 1521 2217 1585
rect 2281 1521 2282 1585
rect 2216 1505 2221 1521
rect 2277 1505 2282 1521
rect 2216 1441 2217 1505
rect 2281 1441 2282 1505
rect 2216 1425 2221 1441
rect 2277 1425 2282 1441
rect 2216 1361 2217 1425
rect 2281 1361 2282 1425
rect 2216 1345 2221 1361
rect 2277 1345 2282 1361
rect 2216 1281 2217 1345
rect 2281 1281 2282 1345
rect 2216 1265 2221 1281
rect 2277 1265 2282 1281
rect 2216 1201 2217 1265
rect 2281 1201 2282 1265
rect 2216 1105 2282 1201
rect 2216 1081 2221 1105
rect 2277 1081 2282 1105
rect 2216 1017 2217 1081
rect 2281 1017 2282 1081
rect 2216 1001 2221 1017
rect 2277 1001 2282 1017
rect 2216 937 2217 1001
rect 2281 937 2282 1001
rect 2216 921 2221 937
rect 2277 921 2282 937
rect 2216 857 2217 921
rect 2281 857 2282 921
rect 2216 841 2221 857
rect 2277 841 2282 857
rect 2216 777 2217 841
rect 2281 777 2282 841
rect 2216 761 2221 777
rect 2277 761 2282 777
rect 2216 697 2217 761
rect 2281 697 2282 761
rect 2216 681 2221 697
rect 2277 681 2282 697
rect 2216 617 2217 681
rect 2281 617 2282 681
rect 2216 601 2221 617
rect 2277 601 2282 617
rect 2216 537 2217 601
rect 2281 537 2282 601
rect 2216 521 2221 537
rect 2277 521 2282 537
rect 2216 457 2217 521
rect 2281 457 2282 521
rect 2216 441 2221 457
rect 2277 441 2282 457
rect 2216 377 2217 441
rect 2281 377 2282 441
rect 2216 361 2221 377
rect 2277 361 2282 377
rect 2216 297 2217 361
rect 2281 297 2282 361
rect 2216 281 2221 297
rect 2277 281 2282 297
rect 2216 217 2217 281
rect 2281 217 2282 281
rect 2216 201 2221 217
rect 2277 201 2282 217
rect 2216 137 2217 201
rect 2281 137 2282 201
rect 2216 121 2221 137
rect 2277 121 2282 137
rect 2216 66 2217 121
rect 65 65 2217 66
rect 65 61 85 65
rect 149 61 165 65
rect 229 61 245 65
rect 309 61 325 65
rect 389 61 405 65
rect 469 61 485 65
rect 549 61 565 65
rect 629 61 645 65
rect 709 61 725 65
rect 789 61 805 65
rect 869 61 885 65
rect 949 61 965 65
rect 1029 61 1045 65
rect 1109 61 1229 65
rect 1293 61 1309 65
rect 1373 61 1389 65
rect 1453 61 1469 65
rect 1533 61 1549 65
rect 1613 61 1629 65
rect 1693 61 1709 65
rect 1773 61 1789 65
rect 1853 61 1869 65
rect 1933 61 1949 65
rect 2013 61 2029 65
rect 2093 61 2109 65
rect 2173 61 2217 65
rect 0 5 61 57
rect 1109 5 1205 61
rect 2281 57 2282 121
rect 2221 5 2282 57
rect 0 1 85 5
rect 149 1 165 5
rect 229 1 245 5
rect 309 1 325 5
rect 389 1 405 5
rect 469 1 485 5
rect 549 1 565 5
rect 629 1 645 5
rect 709 1 725 5
rect 789 1 805 5
rect 869 1 885 5
rect 949 1 965 5
rect 1029 1 1045 5
rect 1109 1 1229 5
rect 1293 1 1309 5
rect 1373 1 1389 5
rect 1453 1 1469 5
rect 1533 1 1549 5
rect 1613 1 1629 5
rect 1693 1 1709 5
rect 1773 1 1789 5
rect 1853 1 1869 5
rect 1933 1 1949 5
rect 2013 1 2029 5
rect 2093 1 2109 5
rect 2173 1 2282 5
rect 0 0 2282 1
<< via3 >>
rect 85 2333 149 2337
rect 165 2333 229 2337
rect 245 2333 309 2337
rect 325 2333 389 2337
rect 405 2333 469 2337
rect 485 2333 549 2337
rect 565 2333 629 2337
rect 645 2333 709 2337
rect 725 2333 789 2337
rect 805 2333 869 2337
rect 885 2333 949 2337
rect 965 2333 1029 2337
rect 1045 2333 1109 2337
rect 1229 2333 1293 2337
rect 1309 2333 1373 2337
rect 1389 2333 1453 2337
rect 1469 2333 1533 2337
rect 1549 2333 1613 2337
rect 1629 2333 1693 2337
rect 1709 2333 1773 2337
rect 1789 2333 1853 2337
rect 1869 2333 1933 2337
rect 1949 2333 2013 2337
rect 2029 2333 2093 2337
rect 2109 2333 2173 2337
rect 85 2277 117 2333
rect 117 2277 141 2333
rect 141 2277 149 2333
rect 165 2277 197 2333
rect 197 2277 221 2333
rect 221 2277 229 2333
rect 245 2277 277 2333
rect 277 2277 301 2333
rect 301 2277 309 2333
rect 325 2277 357 2333
rect 357 2277 381 2333
rect 381 2277 389 2333
rect 405 2277 437 2333
rect 437 2277 461 2333
rect 461 2277 469 2333
rect 485 2277 517 2333
rect 517 2277 541 2333
rect 541 2277 549 2333
rect 565 2277 597 2333
rect 597 2277 621 2333
rect 621 2277 629 2333
rect 645 2277 677 2333
rect 677 2277 701 2333
rect 701 2277 709 2333
rect 725 2277 757 2333
rect 757 2277 781 2333
rect 781 2277 789 2333
rect 805 2277 837 2333
rect 837 2277 861 2333
rect 861 2277 869 2333
rect 885 2277 917 2333
rect 917 2277 941 2333
rect 941 2277 949 2333
rect 965 2277 997 2333
rect 997 2277 1021 2333
rect 1021 2277 1029 2333
rect 1045 2277 1077 2333
rect 1077 2277 1109 2333
rect 1229 2277 1261 2333
rect 1261 2277 1285 2333
rect 1285 2277 1293 2333
rect 1309 2277 1341 2333
rect 1341 2277 1365 2333
rect 1365 2277 1373 2333
rect 1389 2277 1421 2333
rect 1421 2277 1445 2333
rect 1445 2277 1453 2333
rect 1469 2277 1501 2333
rect 1501 2277 1525 2333
rect 1525 2277 1533 2333
rect 1549 2277 1581 2333
rect 1581 2277 1605 2333
rect 1605 2277 1613 2333
rect 1629 2277 1661 2333
rect 1661 2277 1685 2333
rect 1685 2277 1693 2333
rect 1709 2277 1741 2333
rect 1741 2277 1765 2333
rect 1765 2277 1773 2333
rect 1789 2277 1821 2333
rect 1821 2277 1845 2333
rect 1845 2277 1853 2333
rect 1869 2277 1901 2333
rect 1901 2277 1925 2333
rect 1925 2277 1933 2333
rect 1949 2277 1981 2333
rect 1981 2277 2005 2333
rect 2005 2277 2013 2333
rect 2029 2277 2061 2333
rect 2061 2277 2085 2333
rect 2085 2277 2093 2333
rect 2109 2277 2141 2333
rect 2141 2277 2165 2333
rect 2165 2277 2173 2333
rect 85 2273 149 2277
rect 165 2273 229 2277
rect 245 2273 309 2277
rect 325 2273 389 2277
rect 405 2273 469 2277
rect 485 2273 549 2277
rect 565 2273 629 2277
rect 645 2273 709 2277
rect 725 2273 789 2277
rect 805 2273 869 2277
rect 885 2273 949 2277
rect 965 2273 1029 2277
rect 1045 2273 1109 2277
rect 1229 2273 1293 2277
rect 1309 2273 1373 2277
rect 1389 2273 1453 2277
rect 1469 2273 1533 2277
rect 1549 2273 1613 2277
rect 1629 2273 1693 2277
rect 1709 2273 1773 2277
rect 1789 2273 1853 2277
rect 1869 2273 1933 2277
rect 1949 2273 2013 2277
rect 2029 2273 2093 2277
rect 2109 2273 2173 2277
rect 1 2193 5 2225
rect 5 2193 61 2225
rect 61 2193 65 2225
rect 1 2169 65 2193
rect 1 2161 5 2169
rect 5 2161 61 2169
rect 61 2161 65 2169
rect 1 2113 5 2145
rect 5 2113 61 2145
rect 61 2113 65 2145
rect 1 2089 65 2113
rect 1 2081 5 2089
rect 5 2081 61 2089
rect 61 2081 65 2089
rect 1 2033 5 2065
rect 5 2033 61 2065
rect 61 2033 65 2065
rect 1 2009 65 2033
rect 1 2001 5 2009
rect 5 2001 61 2009
rect 61 2001 65 2009
rect 1 1953 5 1985
rect 5 1953 61 1985
rect 61 1953 65 1985
rect 1 1929 65 1953
rect 1 1921 5 1929
rect 5 1921 61 1929
rect 61 1921 65 1929
rect 1 1873 5 1905
rect 5 1873 61 1905
rect 61 1873 65 1905
rect 1 1849 65 1873
rect 1 1841 5 1849
rect 5 1841 61 1849
rect 61 1841 65 1849
rect 1 1793 5 1825
rect 5 1793 61 1825
rect 61 1793 65 1825
rect 1 1769 65 1793
rect 1 1761 5 1769
rect 5 1761 61 1769
rect 61 1761 65 1769
rect 1 1713 5 1745
rect 5 1713 61 1745
rect 61 1713 65 1745
rect 1 1689 65 1713
rect 1 1681 5 1689
rect 5 1681 61 1689
rect 61 1681 65 1689
rect 1 1633 5 1665
rect 5 1633 61 1665
rect 61 1633 65 1665
rect 1 1609 65 1633
rect 1 1601 5 1609
rect 5 1601 61 1609
rect 61 1601 65 1609
rect 1 1553 5 1585
rect 5 1553 61 1585
rect 61 1553 65 1585
rect 1 1529 65 1553
rect 1 1521 5 1529
rect 5 1521 61 1529
rect 61 1521 65 1529
rect 1 1473 5 1505
rect 5 1473 61 1505
rect 61 1473 65 1505
rect 1 1449 65 1473
rect 1 1441 5 1449
rect 5 1441 61 1449
rect 61 1441 65 1449
rect 1 1393 5 1425
rect 5 1393 61 1425
rect 61 1393 65 1425
rect 1 1369 65 1393
rect 1 1361 5 1369
rect 5 1361 61 1369
rect 61 1361 65 1369
rect 1 1313 5 1345
rect 5 1313 61 1345
rect 61 1313 65 1345
rect 1 1289 65 1313
rect 1 1281 5 1289
rect 5 1281 61 1289
rect 61 1281 65 1289
rect 1 1233 5 1265
rect 5 1233 61 1265
rect 61 1233 65 1265
rect 1 1201 65 1233
rect 1 1049 5 1081
rect 5 1049 61 1081
rect 61 1049 65 1081
rect 1 1025 65 1049
rect 1 1017 5 1025
rect 5 1017 61 1025
rect 61 1017 65 1025
rect 1 969 5 1001
rect 5 969 61 1001
rect 61 969 65 1001
rect 1 945 65 969
rect 1 937 5 945
rect 5 937 61 945
rect 61 937 65 945
rect 1 889 5 921
rect 5 889 61 921
rect 61 889 65 921
rect 1 865 65 889
rect 1 857 5 865
rect 5 857 61 865
rect 61 857 65 865
rect 1 809 5 841
rect 5 809 61 841
rect 61 809 65 841
rect 1 785 65 809
rect 1 777 5 785
rect 5 777 61 785
rect 61 777 65 785
rect 1 729 5 761
rect 5 729 61 761
rect 61 729 65 761
rect 1 705 65 729
rect 1 697 5 705
rect 5 697 61 705
rect 61 697 65 705
rect 1 649 5 681
rect 5 649 61 681
rect 61 649 65 681
rect 1 625 65 649
rect 1 617 5 625
rect 5 617 61 625
rect 61 617 65 625
rect 1 569 5 601
rect 5 569 61 601
rect 61 569 65 601
rect 1 545 65 569
rect 1 537 5 545
rect 5 537 61 545
rect 61 537 65 545
rect 1 489 5 521
rect 5 489 61 521
rect 61 489 65 521
rect 1 465 65 489
rect 1 457 5 465
rect 5 457 61 465
rect 61 457 65 465
rect 1 409 5 441
rect 5 409 61 441
rect 61 409 65 441
rect 1 385 65 409
rect 1 377 5 385
rect 5 377 61 385
rect 61 377 65 385
rect 1 329 5 361
rect 5 329 61 361
rect 61 329 65 361
rect 1 305 65 329
rect 1 297 5 305
rect 5 297 61 305
rect 61 297 65 305
rect 1 249 5 281
rect 5 249 61 281
rect 61 249 65 281
rect 1 225 65 249
rect 1 217 5 225
rect 5 217 61 225
rect 61 217 65 225
rect 1 169 5 201
rect 5 169 61 201
rect 61 169 65 201
rect 1 145 65 169
rect 1 137 5 145
rect 5 137 61 145
rect 61 137 65 145
rect 1109 2157 1173 2161
rect 1109 2101 1113 2157
rect 1113 2101 1169 2157
rect 1169 2101 1173 2157
rect 1109 2097 1173 2101
rect 1109 2077 1173 2081
rect 1109 2021 1113 2077
rect 1113 2021 1169 2077
rect 1169 2021 1173 2077
rect 1109 2017 1173 2021
rect 1109 1997 1173 2001
rect 1109 1941 1113 1997
rect 1113 1941 1169 1997
rect 1169 1941 1173 1997
rect 1109 1937 1173 1941
rect 1109 1917 1173 1921
rect 1109 1861 1113 1917
rect 1113 1861 1169 1917
rect 1169 1861 1173 1917
rect 1109 1857 1173 1861
rect 1109 1837 1173 1841
rect 1109 1781 1113 1837
rect 1113 1781 1169 1837
rect 1169 1781 1173 1837
rect 1109 1777 1173 1781
rect 1109 1757 1173 1761
rect 1109 1701 1113 1757
rect 1113 1701 1169 1757
rect 1169 1701 1173 1757
rect 1109 1697 1173 1701
rect 1109 1677 1173 1681
rect 1109 1621 1113 1677
rect 1113 1621 1169 1677
rect 1169 1621 1173 1677
rect 1109 1617 1173 1621
rect 1109 1597 1173 1601
rect 1109 1541 1113 1597
rect 1113 1541 1169 1597
rect 1169 1541 1173 1597
rect 1109 1537 1173 1541
rect 1109 1517 1173 1521
rect 1109 1461 1113 1517
rect 1113 1461 1169 1517
rect 1169 1461 1173 1517
rect 1109 1457 1173 1461
rect 1109 1437 1173 1441
rect 1109 1381 1113 1437
rect 1113 1381 1169 1437
rect 1169 1381 1173 1437
rect 1109 1377 1173 1381
rect 1109 1357 1173 1361
rect 1109 1301 1113 1357
rect 1113 1301 1169 1357
rect 1169 1301 1173 1357
rect 1109 1297 1173 1301
rect 1109 1277 1173 1281
rect 1109 1221 1113 1277
rect 1113 1221 1169 1277
rect 1169 1221 1173 1277
rect 1109 1217 1173 1221
rect 149 1197 213 1201
rect 149 1141 153 1197
rect 153 1141 209 1197
rect 209 1141 213 1197
rect 149 1137 213 1141
rect 229 1197 293 1201
rect 229 1141 233 1197
rect 233 1141 289 1197
rect 289 1141 293 1197
rect 229 1137 293 1141
rect 309 1197 373 1201
rect 309 1141 313 1197
rect 313 1141 369 1197
rect 369 1141 373 1197
rect 309 1137 373 1141
rect 389 1197 453 1201
rect 389 1141 393 1197
rect 393 1141 449 1197
rect 449 1141 453 1197
rect 389 1137 453 1141
rect 469 1197 533 1201
rect 469 1141 473 1197
rect 473 1141 529 1197
rect 529 1141 533 1197
rect 469 1137 533 1141
rect 549 1197 613 1201
rect 549 1141 553 1197
rect 553 1141 609 1197
rect 609 1141 613 1197
rect 549 1137 613 1141
rect 629 1197 693 1201
rect 629 1141 633 1197
rect 633 1141 689 1197
rect 689 1141 693 1197
rect 629 1137 693 1141
rect 709 1197 773 1201
rect 709 1141 713 1197
rect 713 1141 769 1197
rect 769 1141 773 1197
rect 709 1137 773 1141
rect 789 1197 853 1201
rect 789 1141 793 1197
rect 793 1141 849 1197
rect 849 1141 853 1197
rect 789 1137 853 1141
rect 869 1197 933 1201
rect 869 1141 873 1197
rect 873 1141 929 1197
rect 929 1141 933 1197
rect 869 1137 933 1141
rect 949 1197 1013 1201
rect 949 1141 953 1197
rect 953 1141 1009 1197
rect 1009 1141 1013 1197
rect 949 1137 1013 1141
rect 1029 1197 1093 1201
rect 1029 1141 1033 1197
rect 1033 1141 1089 1197
rect 1089 1141 1093 1197
rect 1029 1137 1093 1141
rect 1109 1197 1173 1201
rect 1109 1141 1113 1197
rect 1113 1141 1169 1197
rect 1169 1141 1173 1197
rect 1109 1137 1173 1141
rect 1189 1197 1253 1201
rect 1189 1141 1193 1197
rect 1193 1141 1249 1197
rect 1249 1141 1253 1197
rect 1189 1137 1253 1141
rect 1269 1197 1333 1201
rect 1269 1141 1273 1197
rect 1273 1141 1329 1197
rect 1329 1141 1333 1197
rect 1269 1137 1333 1141
rect 1349 1197 1413 1201
rect 1349 1141 1353 1197
rect 1353 1141 1409 1197
rect 1409 1141 1413 1197
rect 1349 1137 1413 1141
rect 1429 1197 1493 1201
rect 1429 1141 1433 1197
rect 1433 1141 1489 1197
rect 1489 1141 1493 1197
rect 1429 1137 1493 1141
rect 1509 1197 1573 1201
rect 1509 1141 1513 1197
rect 1513 1141 1569 1197
rect 1569 1141 1573 1197
rect 1509 1137 1573 1141
rect 1589 1197 1653 1201
rect 1589 1141 1593 1197
rect 1593 1141 1649 1197
rect 1649 1141 1653 1197
rect 1589 1137 1653 1141
rect 1669 1197 1733 1201
rect 1669 1141 1673 1197
rect 1673 1141 1729 1197
rect 1729 1141 1733 1197
rect 1669 1137 1733 1141
rect 1749 1197 1813 1201
rect 1749 1141 1753 1197
rect 1753 1141 1809 1197
rect 1809 1141 1813 1197
rect 1749 1137 1813 1141
rect 1829 1197 1893 1201
rect 1829 1141 1833 1197
rect 1833 1141 1889 1197
rect 1889 1141 1893 1197
rect 1829 1137 1893 1141
rect 1909 1197 1973 1201
rect 1909 1141 1913 1197
rect 1913 1141 1969 1197
rect 1969 1141 1973 1197
rect 1909 1137 1973 1141
rect 1989 1197 2053 1201
rect 1989 1141 1993 1197
rect 1993 1141 2049 1197
rect 2049 1141 2053 1197
rect 1989 1137 2053 1141
rect 2069 1197 2133 1201
rect 2069 1141 2073 1197
rect 2073 1141 2129 1197
rect 2129 1141 2133 1197
rect 2069 1137 2133 1141
rect 1 89 5 121
rect 5 89 61 121
rect 61 89 65 121
rect 1 61 65 89
rect 1109 1117 1173 1121
rect 1109 1061 1113 1117
rect 1113 1061 1169 1117
rect 1169 1061 1173 1117
rect 1109 1057 1173 1061
rect 1109 1037 1173 1041
rect 1109 981 1113 1037
rect 1113 981 1169 1037
rect 1169 981 1173 1037
rect 1109 977 1173 981
rect 1109 957 1173 961
rect 1109 901 1113 957
rect 1113 901 1169 957
rect 1169 901 1173 957
rect 1109 897 1173 901
rect 1109 877 1173 881
rect 1109 821 1113 877
rect 1113 821 1169 877
rect 1169 821 1173 877
rect 1109 817 1173 821
rect 1109 797 1173 801
rect 1109 741 1113 797
rect 1113 741 1169 797
rect 1169 741 1173 797
rect 1109 737 1173 741
rect 1109 717 1173 721
rect 1109 661 1113 717
rect 1113 661 1169 717
rect 1169 661 1173 717
rect 1109 657 1173 661
rect 1109 637 1173 641
rect 1109 581 1113 637
rect 1113 581 1169 637
rect 1169 581 1173 637
rect 1109 577 1173 581
rect 1109 557 1173 561
rect 1109 501 1113 557
rect 1113 501 1169 557
rect 1169 501 1173 557
rect 1109 497 1173 501
rect 1109 477 1173 481
rect 1109 421 1113 477
rect 1113 421 1169 477
rect 1169 421 1173 477
rect 1109 417 1173 421
rect 1109 397 1173 401
rect 1109 341 1113 397
rect 1113 341 1169 397
rect 1169 341 1173 397
rect 1109 337 1173 341
rect 1109 317 1173 321
rect 1109 261 1113 317
rect 1113 261 1169 317
rect 1169 261 1173 317
rect 1109 257 1173 261
rect 1109 237 1173 241
rect 1109 181 1113 237
rect 1113 181 1169 237
rect 1169 181 1173 237
rect 1109 177 1173 181
rect 2217 2193 2221 2225
rect 2221 2193 2277 2225
rect 2277 2193 2281 2225
rect 2217 2169 2281 2193
rect 2217 2161 2221 2169
rect 2221 2161 2277 2169
rect 2277 2161 2281 2169
rect 2217 2113 2221 2145
rect 2221 2113 2277 2145
rect 2277 2113 2281 2145
rect 2217 2089 2281 2113
rect 2217 2081 2221 2089
rect 2221 2081 2277 2089
rect 2277 2081 2281 2089
rect 2217 2033 2221 2065
rect 2221 2033 2277 2065
rect 2277 2033 2281 2065
rect 2217 2009 2281 2033
rect 2217 2001 2221 2009
rect 2221 2001 2277 2009
rect 2277 2001 2281 2009
rect 2217 1953 2221 1985
rect 2221 1953 2277 1985
rect 2277 1953 2281 1985
rect 2217 1929 2281 1953
rect 2217 1921 2221 1929
rect 2221 1921 2277 1929
rect 2277 1921 2281 1929
rect 2217 1873 2221 1905
rect 2221 1873 2277 1905
rect 2277 1873 2281 1905
rect 2217 1849 2281 1873
rect 2217 1841 2221 1849
rect 2221 1841 2277 1849
rect 2277 1841 2281 1849
rect 2217 1793 2221 1825
rect 2221 1793 2277 1825
rect 2277 1793 2281 1825
rect 2217 1769 2281 1793
rect 2217 1761 2221 1769
rect 2221 1761 2277 1769
rect 2277 1761 2281 1769
rect 2217 1713 2221 1745
rect 2221 1713 2277 1745
rect 2277 1713 2281 1745
rect 2217 1689 2281 1713
rect 2217 1681 2221 1689
rect 2221 1681 2277 1689
rect 2277 1681 2281 1689
rect 2217 1633 2221 1665
rect 2221 1633 2277 1665
rect 2277 1633 2281 1665
rect 2217 1609 2281 1633
rect 2217 1601 2221 1609
rect 2221 1601 2277 1609
rect 2277 1601 2281 1609
rect 2217 1553 2221 1585
rect 2221 1553 2277 1585
rect 2277 1553 2281 1585
rect 2217 1529 2281 1553
rect 2217 1521 2221 1529
rect 2221 1521 2277 1529
rect 2277 1521 2281 1529
rect 2217 1473 2221 1505
rect 2221 1473 2277 1505
rect 2277 1473 2281 1505
rect 2217 1449 2281 1473
rect 2217 1441 2221 1449
rect 2221 1441 2277 1449
rect 2277 1441 2281 1449
rect 2217 1393 2221 1425
rect 2221 1393 2277 1425
rect 2277 1393 2281 1425
rect 2217 1369 2281 1393
rect 2217 1361 2221 1369
rect 2221 1361 2277 1369
rect 2277 1361 2281 1369
rect 2217 1313 2221 1345
rect 2221 1313 2277 1345
rect 2277 1313 2281 1345
rect 2217 1289 2281 1313
rect 2217 1281 2221 1289
rect 2221 1281 2277 1289
rect 2277 1281 2281 1289
rect 2217 1233 2221 1265
rect 2221 1233 2277 1265
rect 2277 1233 2281 1265
rect 2217 1201 2281 1233
rect 2217 1049 2221 1081
rect 2221 1049 2277 1081
rect 2277 1049 2281 1081
rect 2217 1025 2281 1049
rect 2217 1017 2221 1025
rect 2221 1017 2277 1025
rect 2277 1017 2281 1025
rect 2217 969 2221 1001
rect 2221 969 2277 1001
rect 2277 969 2281 1001
rect 2217 945 2281 969
rect 2217 937 2221 945
rect 2221 937 2277 945
rect 2277 937 2281 945
rect 2217 889 2221 921
rect 2221 889 2277 921
rect 2277 889 2281 921
rect 2217 865 2281 889
rect 2217 857 2221 865
rect 2221 857 2277 865
rect 2277 857 2281 865
rect 2217 809 2221 841
rect 2221 809 2277 841
rect 2277 809 2281 841
rect 2217 785 2281 809
rect 2217 777 2221 785
rect 2221 777 2277 785
rect 2277 777 2281 785
rect 2217 729 2221 761
rect 2221 729 2277 761
rect 2277 729 2281 761
rect 2217 705 2281 729
rect 2217 697 2221 705
rect 2221 697 2277 705
rect 2277 697 2281 705
rect 2217 649 2221 681
rect 2221 649 2277 681
rect 2277 649 2281 681
rect 2217 625 2281 649
rect 2217 617 2221 625
rect 2221 617 2277 625
rect 2277 617 2281 625
rect 2217 569 2221 601
rect 2221 569 2277 601
rect 2277 569 2281 601
rect 2217 545 2281 569
rect 2217 537 2221 545
rect 2221 537 2277 545
rect 2277 537 2281 545
rect 2217 489 2221 521
rect 2221 489 2277 521
rect 2277 489 2281 521
rect 2217 465 2281 489
rect 2217 457 2221 465
rect 2221 457 2277 465
rect 2277 457 2281 465
rect 2217 409 2221 441
rect 2221 409 2277 441
rect 2277 409 2281 441
rect 2217 385 2281 409
rect 2217 377 2221 385
rect 2221 377 2277 385
rect 2277 377 2281 385
rect 2217 329 2221 361
rect 2221 329 2277 361
rect 2277 329 2281 361
rect 2217 305 2281 329
rect 2217 297 2221 305
rect 2221 297 2277 305
rect 2277 297 2281 305
rect 2217 249 2221 281
rect 2221 249 2277 281
rect 2277 249 2281 281
rect 2217 225 2281 249
rect 2217 217 2221 225
rect 2221 217 2277 225
rect 2277 217 2281 225
rect 2217 169 2221 201
rect 2221 169 2277 201
rect 2277 169 2281 201
rect 2217 145 2281 169
rect 2217 137 2221 145
rect 2221 137 2277 145
rect 2277 137 2281 145
rect 2217 89 2221 121
rect 2221 89 2277 121
rect 2277 89 2281 121
rect 85 61 149 65
rect 165 61 229 65
rect 245 61 309 65
rect 325 61 389 65
rect 405 61 469 65
rect 485 61 549 65
rect 565 61 629 65
rect 645 61 709 65
rect 725 61 789 65
rect 805 61 869 65
rect 885 61 949 65
rect 965 61 1029 65
rect 1045 61 1109 65
rect 1229 61 1293 65
rect 1309 61 1373 65
rect 1389 61 1453 65
rect 1469 61 1533 65
rect 1549 61 1613 65
rect 1629 61 1693 65
rect 1709 61 1773 65
rect 1789 61 1853 65
rect 1869 61 1933 65
rect 1949 61 2013 65
rect 2029 61 2093 65
rect 2109 61 2173 65
rect 2217 61 2281 89
rect 1 57 61 61
rect 61 57 65 61
rect 85 5 117 61
rect 117 5 141 61
rect 141 5 149 61
rect 165 5 197 61
rect 197 5 221 61
rect 221 5 229 61
rect 245 5 277 61
rect 277 5 301 61
rect 301 5 309 61
rect 325 5 357 61
rect 357 5 381 61
rect 381 5 389 61
rect 405 5 437 61
rect 437 5 461 61
rect 461 5 469 61
rect 485 5 517 61
rect 517 5 541 61
rect 541 5 549 61
rect 565 5 597 61
rect 597 5 621 61
rect 621 5 629 61
rect 645 5 677 61
rect 677 5 701 61
rect 701 5 709 61
rect 725 5 757 61
rect 757 5 781 61
rect 781 5 789 61
rect 805 5 837 61
rect 837 5 861 61
rect 861 5 869 61
rect 885 5 917 61
rect 917 5 941 61
rect 941 5 949 61
rect 965 5 997 61
rect 997 5 1021 61
rect 1021 5 1029 61
rect 1045 5 1077 61
rect 1077 5 1109 61
rect 1229 5 1261 61
rect 1261 5 1285 61
rect 1285 5 1293 61
rect 1309 5 1341 61
rect 1341 5 1365 61
rect 1365 5 1373 61
rect 1389 5 1421 61
rect 1421 5 1445 61
rect 1445 5 1453 61
rect 1469 5 1501 61
rect 1501 5 1525 61
rect 1525 5 1533 61
rect 1549 5 1581 61
rect 1581 5 1605 61
rect 1605 5 1613 61
rect 1629 5 1661 61
rect 1661 5 1685 61
rect 1685 5 1693 61
rect 1709 5 1741 61
rect 1741 5 1765 61
rect 1765 5 1773 61
rect 1789 5 1821 61
rect 1821 5 1845 61
rect 1845 5 1853 61
rect 1869 5 1901 61
rect 1901 5 1925 61
rect 1925 5 1933 61
rect 1949 5 1981 61
rect 1981 5 2005 61
rect 2005 5 2013 61
rect 2029 5 2061 61
rect 2061 5 2085 61
rect 2085 5 2093 61
rect 2109 5 2141 61
rect 2141 5 2165 61
rect 2165 5 2173 61
rect 2217 57 2221 61
rect 2221 57 2281 61
rect 85 1 149 5
rect 165 1 229 5
rect 245 1 309 5
rect 325 1 389 5
rect 405 1 469 5
rect 485 1 549 5
rect 565 1 629 5
rect 645 1 709 5
rect 725 1 789 5
rect 805 1 869 5
rect 885 1 949 5
rect 965 1 1029 5
rect 1045 1 1109 5
rect 1229 1 1293 5
rect 1309 1 1373 5
rect 1389 1 1453 5
rect 1469 1 1533 5
rect 1549 1 1613 5
rect 1629 1 1693 5
rect 1709 1 1773 5
rect 1789 1 1853 5
rect 1869 1 1933 5
rect 1949 1 2013 5
rect 2029 1 2093 5
rect 2109 1 2173 5
<< metal4 >>
rect 0 2337 2282 2338
rect 0 2273 85 2337
rect 149 2273 165 2337
rect 229 2273 245 2337
rect 309 2273 325 2337
rect 389 2273 405 2337
rect 469 2273 485 2337
rect 549 2273 565 2337
rect 629 2273 645 2337
rect 709 2273 725 2337
rect 789 2273 805 2337
rect 869 2273 885 2337
rect 949 2273 965 2337
rect 1029 2273 1045 2337
rect 1109 2273 1229 2337
rect 1293 2273 1309 2337
rect 1373 2273 1389 2337
rect 1453 2273 1469 2337
rect 1533 2273 1549 2337
rect 1613 2273 1629 2337
rect 1693 2273 1709 2337
rect 1773 2273 1789 2337
rect 1853 2273 1869 2337
rect 1933 2273 1949 2337
rect 2013 2273 2029 2337
rect 2093 2273 2109 2337
rect 2173 2273 2282 2337
rect 0 2272 2282 2273
rect 0 2225 66 2272
rect 0 2161 1 2225
rect 65 2161 66 2225
rect 2216 2225 2282 2272
rect 0 2145 66 2161
rect 126 2161 2156 2212
rect 126 2152 1109 2161
rect 0 2081 1 2145
rect 65 2092 66 2145
rect 1108 2097 1109 2152
rect 1173 2152 2156 2161
rect 2216 2161 2217 2225
rect 2281 2161 2282 2225
rect 1173 2097 1174 2152
rect 65 2081 1048 2092
rect 0 2065 1048 2081
rect 0 2001 1 2065
rect 65 2032 1048 2065
rect 1108 2081 1174 2097
rect 2216 2145 2282 2161
rect 2216 2092 2217 2145
rect 65 2001 66 2032
rect 0 1985 66 2001
rect 0 1921 1 1985
rect 65 1921 66 1985
rect 1108 2017 1109 2081
rect 1173 2017 1174 2081
rect 1234 2081 2217 2092
rect 2281 2081 2282 2145
rect 1234 2065 2282 2081
rect 1234 2032 2217 2065
rect 1108 2001 1174 2017
rect 1108 1972 1109 2001
rect 0 1905 66 1921
rect 126 1937 1109 1972
rect 1173 1972 1174 2001
rect 2216 2001 2217 2032
rect 2281 2001 2282 2065
rect 2216 1985 2282 2001
rect 1173 1937 2156 1972
rect 126 1921 2156 1937
rect 126 1912 1109 1921
rect 0 1841 1 1905
rect 65 1852 66 1905
rect 1108 1857 1109 1912
rect 1173 1912 2156 1921
rect 2216 1921 2217 1985
rect 2281 1921 2282 1985
rect 1173 1857 1174 1912
rect 65 1841 1048 1852
rect 0 1825 1048 1841
rect 0 1761 1 1825
rect 65 1792 1048 1825
rect 1108 1841 1174 1857
rect 2216 1905 2282 1921
rect 2216 1852 2217 1905
rect 65 1761 66 1792
rect 0 1745 66 1761
rect 0 1681 1 1745
rect 65 1681 66 1745
rect 1108 1777 1109 1841
rect 1173 1777 1174 1841
rect 1234 1841 2217 1852
rect 2281 1841 2282 1905
rect 1234 1825 2282 1841
rect 1234 1792 2217 1825
rect 1108 1761 1174 1777
rect 1108 1732 1109 1761
rect 0 1665 66 1681
rect 126 1697 1109 1732
rect 1173 1732 1174 1761
rect 2216 1761 2217 1792
rect 2281 1761 2282 1825
rect 2216 1745 2282 1761
rect 1173 1697 2156 1732
rect 126 1681 2156 1697
rect 126 1672 1109 1681
rect 0 1601 1 1665
rect 65 1612 66 1665
rect 1108 1617 1109 1672
rect 1173 1672 2156 1681
rect 2216 1681 2217 1745
rect 2281 1681 2282 1745
rect 1173 1617 1174 1672
rect 65 1601 1048 1612
rect 0 1585 1048 1601
rect 0 1521 1 1585
rect 65 1532 1048 1585
rect 1108 1601 1174 1617
rect 2216 1665 2282 1681
rect 2216 1612 2217 1665
rect 1108 1537 1109 1601
rect 1173 1537 1174 1601
rect 65 1521 66 1532
rect 0 1505 66 1521
rect 0 1441 1 1505
rect 65 1441 66 1505
rect 1108 1521 1174 1537
rect 1234 1601 2217 1612
rect 2281 1601 2282 1665
rect 1234 1585 2282 1601
rect 1234 1532 2217 1585
rect 1108 1472 1109 1521
rect 0 1425 66 1441
rect 0 1361 1 1425
rect 65 1361 66 1425
rect 126 1457 1109 1472
rect 1173 1472 1174 1521
rect 2216 1521 2217 1532
rect 2281 1521 2282 1585
rect 2216 1505 2282 1521
rect 1173 1457 2156 1472
rect 126 1441 2156 1457
rect 126 1412 1109 1441
rect 0 1352 66 1361
rect 1108 1377 1109 1412
rect 1173 1412 2156 1441
rect 2216 1441 2217 1505
rect 2281 1441 2282 1505
rect 2216 1425 2282 1441
rect 1173 1377 1174 1412
rect 1108 1361 1174 1377
rect 0 1345 1048 1352
rect 0 1281 1 1345
rect 65 1281 1048 1345
rect 0 1265 1048 1281
rect 0 1201 1 1265
rect 65 1262 1048 1265
rect 1108 1297 1109 1361
rect 1173 1297 1174 1361
rect 2216 1361 2217 1425
rect 2281 1361 2282 1425
rect 2216 1352 2282 1361
rect 1108 1281 1174 1297
rect 65 1201 66 1262
rect 1108 1217 1109 1281
rect 1173 1217 1174 1281
rect 1234 1345 2282 1352
rect 1234 1281 2217 1345
rect 2281 1281 2282 1345
rect 1234 1265 2282 1281
rect 1234 1262 2217 1265
rect 1108 1202 1174 1217
rect 0 1081 66 1201
rect 126 1201 2156 1202
rect 126 1137 149 1201
rect 213 1137 229 1201
rect 293 1137 309 1201
rect 373 1137 389 1201
rect 453 1137 469 1201
rect 533 1137 549 1201
rect 613 1137 629 1201
rect 693 1137 709 1201
rect 773 1137 789 1201
rect 853 1137 869 1201
rect 933 1137 949 1201
rect 1013 1137 1029 1201
rect 1093 1137 1109 1201
rect 1173 1137 1189 1201
rect 1253 1137 1269 1201
rect 1333 1137 1349 1201
rect 1413 1137 1429 1201
rect 1493 1137 1509 1201
rect 1573 1137 1589 1201
rect 1653 1137 1669 1201
rect 1733 1137 1749 1201
rect 1813 1137 1829 1201
rect 1893 1137 1909 1201
rect 1973 1137 1989 1201
rect 2053 1137 2069 1201
rect 2133 1137 2156 1201
rect 126 1136 2156 1137
rect 2216 1201 2217 1262
rect 2281 1201 2282 1265
rect 0 1017 1 1081
rect 65 1076 66 1081
rect 1108 1121 1174 1136
rect 65 1017 1048 1076
rect 0 1001 1048 1017
rect 0 937 1 1001
rect 65 986 1048 1001
rect 1108 1057 1109 1121
rect 1173 1057 1174 1121
rect 2216 1081 2282 1201
rect 2216 1076 2217 1081
rect 1108 1041 1174 1057
rect 65 937 66 986
rect 0 921 66 937
rect 1108 977 1109 1041
rect 1173 977 1174 1041
rect 1234 1017 2217 1076
rect 2281 1017 2282 1081
rect 1234 1001 2282 1017
rect 1234 986 2217 1001
rect 1108 961 1174 977
rect 1108 926 1109 961
rect 0 857 1 921
rect 65 857 66 921
rect 126 897 1109 926
rect 1173 926 1174 961
rect 2216 937 2217 986
rect 2281 937 2282 1001
rect 1173 897 2156 926
rect 126 881 2156 897
rect 126 866 1109 881
rect 0 841 66 857
rect 0 777 1 841
rect 65 806 66 841
rect 1108 817 1109 866
rect 1173 866 2156 881
rect 2216 921 2282 937
rect 1173 817 1174 866
rect 65 777 1048 806
rect 0 761 1048 777
rect 0 697 1 761
rect 65 726 1048 761
rect 1108 801 1174 817
rect 2216 857 2217 921
rect 2281 857 2282 921
rect 2216 841 2282 857
rect 2216 806 2217 841
rect 1108 737 1109 801
rect 1173 737 1174 801
rect 65 697 66 726
rect 0 681 66 697
rect 0 617 1 681
rect 65 617 66 681
rect 1108 721 1174 737
rect 1234 777 2217 806
rect 2281 777 2282 841
rect 1234 761 2282 777
rect 1234 726 2217 761
rect 1108 666 1109 721
rect 0 601 66 617
rect 126 657 1109 666
rect 1173 666 1174 721
rect 2216 697 2217 726
rect 2281 697 2282 761
rect 2216 681 2282 697
rect 1173 657 2156 666
rect 126 641 2156 657
rect 126 606 1109 641
rect 0 537 1 601
rect 65 546 66 601
rect 1108 577 1109 606
rect 1173 606 2156 641
rect 2216 617 2217 681
rect 2281 617 2282 681
rect 1173 577 1174 606
rect 1108 561 1174 577
rect 65 537 1048 546
rect 0 521 1048 537
rect 0 457 1 521
rect 65 486 1048 521
rect 1108 497 1109 561
rect 1173 497 1174 561
rect 2216 601 2282 617
rect 2216 546 2217 601
rect 65 457 66 486
rect 0 441 66 457
rect 0 377 1 441
rect 65 377 66 441
rect 1108 481 1174 497
rect 1234 537 2217 546
rect 2281 537 2282 601
rect 1234 521 2282 537
rect 1234 486 2217 521
rect 1108 426 1109 481
rect 0 361 66 377
rect 126 417 1109 426
rect 1173 426 1174 481
rect 2216 457 2217 486
rect 2281 457 2282 521
rect 2216 441 2282 457
rect 1173 417 2156 426
rect 126 401 2156 417
rect 126 366 1109 401
rect 0 297 1 361
rect 65 306 66 361
rect 1108 337 1109 366
rect 1173 366 2156 401
rect 2216 377 2217 441
rect 2281 377 2282 441
rect 1173 337 1174 366
rect 1108 321 1174 337
rect 65 297 1048 306
rect 0 281 1048 297
rect 0 217 1 281
rect 65 246 1048 281
rect 1108 257 1109 321
rect 1173 257 1174 321
rect 2216 361 2282 377
rect 2216 306 2217 361
rect 65 217 66 246
rect 0 201 66 217
rect 0 137 1 201
rect 65 137 66 201
rect 1108 241 1174 257
rect 1234 297 2217 306
rect 2281 297 2282 361
rect 1234 281 2282 297
rect 1234 246 2217 281
rect 1108 186 1109 241
rect 0 121 66 137
rect 126 177 1109 186
rect 1173 186 1174 241
rect 2216 217 2217 246
rect 2281 217 2282 281
rect 2216 201 2282 217
rect 1173 177 2156 186
rect 126 126 2156 177
rect 2216 137 2217 201
rect 2281 137 2282 201
rect 0 57 1 121
rect 65 66 66 121
rect 2216 121 2282 137
rect 2216 66 2217 121
rect 65 65 2217 66
rect 65 57 85 65
rect 0 1 85 57
rect 149 1 165 65
rect 229 1 245 65
rect 309 1 325 65
rect 389 1 405 65
rect 469 1 485 65
rect 549 1 565 65
rect 629 1 645 65
rect 709 1 725 65
rect 789 1 805 65
rect 869 1 885 65
rect 949 1 965 65
rect 1029 1 1045 65
rect 1109 1 1229 65
rect 1293 1 1309 65
rect 1373 1 1389 65
rect 1453 1 1469 65
rect 1533 1 1549 65
rect 1613 1 1629 65
rect 1693 1 1709 65
rect 1773 1 1789 65
rect 1853 1 1869 65
rect 1933 1 1949 65
rect 2013 1 2029 65
rect 2093 1 2109 65
rect 2173 57 2217 65
rect 2281 57 2282 121
rect 2173 1 2282 57
rect 0 0 2282 1
<< metal5 >>
rect 0 1889 2282 2338
rect 0 1429 421 1889
rect 881 1429 1401 1889
rect 1861 1429 2282 1889
rect 0 909 2282 1429
rect 0 449 421 909
rect 881 449 1401 909
rect 1861 449 2282 909
rect 0 0 2282 449
<< labels >>
flabel metal2 s 1019 2162 1049 2186 0 FreeSans 200 0 0 0 C0
port 1 nsew
flabel metal2 s 1121 2079 1163 2115 0 FreeSans 200 0 0 0 C1
port 2 nsew
flabel metal5 s 1107 536 1194 631 0 FreeSans 200 0 0 0 MET5
port 3 nsew
flabel pwell s 1176 1289 1197 1338 0 FreeSans 2000 0 0 0 SUB
port 4 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 1164156
string GDS_START 1116270
<< end >>
