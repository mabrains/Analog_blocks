* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__pfet_01v8__toxe_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8__vth0_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8__voff_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8__nfactor_slope_spectre = 0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__pfet_01v8__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt  sky130_fd_pr__pfet_01v8 d g s b
+ 
.param  l = 1 w = 1 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1 
msky130_fd_pr__pfet_01v8 d g s b sky130_fd_pr__pfet_01v8__model l = {l} w = {w} nf = {nf} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd} 
.model sky130_fd_pr__pfet_01v8__model.0 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0498303+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43448553
+ k2 = 0.021784346
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 160312.5
+ ua = -5.9240701e-10
+ ub = 9.3030446e-19
+ uc = -6.6549964e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0104306
+ a0 = 1.171369
+ keta = 0.0051290095
+ a1 = 0.0
+ a2 = 0.9995
+ ags = 0.2846738
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.28370745+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.3961358+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0015228006
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029632464
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 9.3760948e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.6464006
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1181082000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.4485
+ kt2 = -0.0075706
+ at = 90900.0
+ ute = -0.33954
+ ua1 = 1.6104e-9
+ ub1 = -5.609e-19
+ uc1 = -1.0858e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.1 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0498303+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43448553
+ k2 = 0.021784346
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 160312.5
+ ua = -5.9240701e-10
+ ub = 9.3030446e-19
+ uc = -6.6549964e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0104306
+ a0 = 1.171369
+ keta = 0.0051290095
+ a1 = 0.0
+ a2 = 0.9995
+ ags = 0.2846738
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.28370745+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.3961358+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0015228006
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0029632464
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 9.3760948e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.6464006
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1181082000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.4485
+ kt2 = -0.0075706
+ at = 90900.0
+ ute = -0.33954
+ ua1 = 1.6104e-9
+ ub1 = -5.609e-19
+ uc1 = -1.0858e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.2 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.05406354699422+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.38817786648298e-8
+ k1 = 0.438111540819447 lk1 = -2.90216224539694e-8
+ k2 = 0.020847100130831 lk2 = 7.50146569218161e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 267287.24109375 lvsat = -0.856197265458503
+ ua = -6.30146567603303e-10 lua = 3.02057342594953e-16
+ ub = 9.25585349996893e-19 lub = 3.77704964625017e-26
+ uc = -7.3185202562779e-11 luc = 5.31066778477869e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.010066360390325 lu0 = 2.91527658386293e-9
+ a0 = 1.230540170007 la0 = -4.73590246033636e-7
+ keta = 0.0213585060556696 lketa = -1.29896557155999e-07 pketa = 1.0097419586829e-28
+ a1 = 0.0
+ a2 = 1.199186183375 la2 = -1.59823489552254e-06 wa2 = 1.6940658945086e-21
+ ags = 0.24265758492742 lags = 3.36286567111506e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.298175649858108+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.15799608654931e-7
+ nfactor = {1.25726101594877+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.11151669197867e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.430980526189767 lpclm = 3.46164114923705e-06 wpclm = -1.52201232709757e-22 ppclm = 3.40787911055477e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00577216450866307 lpdiblc2 = -2.24818305606042e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.01371115566944e-08 lpscbe2 = -6.09097492910795e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.25291554260215 lbeta0 = 1.11530823389021e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 8.43618292846325e-11 lagidl = 1.25163743014221e-16
+ bgidl = 1362332994.7765 lbgidl = -1450.6845681755
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.431675573243395 lkt1 = -1.34658219637922e-7
+ kt2 = 0.00969919300712574 lkt2 = -1.38222812194302e-07 pkt2 = -1.0097419586829e-28
+ at = 87878.4127328975 lat = 0.0241839777220882
+ ute = -0.47361144551513 lute = 1.07307205282715e-6
+ ua1 = 1.22619747730703e-09 lua1 = 3.07505440956101e-15
+ ub1 = -3.0097092736856e-19 lub1 = -2.08040289627965e-24
+ uc1 = -8.842508796601e-11 luc1 = -1.61314534558543e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.3 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.055275022924+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.87322048235757e-8
+ k1 = 0.424351018216625 lk1 = 2.60718359881974e-8
+ k2 = 0.024934107594989 lk2 = -8.86182096331409e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 53437.5
+ ua = -2.33552580158625e-10 lua = -1.28579909253889e-15
+ ub = 7.69195707129755e-19 lub = 6.63912870467874e-25
+ uc = -8.0640895799503e-11 luc = 8.29572828975356e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0123850632554 lu0 = -6.36819059423241e-9
+ a0 = 1.1425925232195 la0 = -1.21471350318178e-7
+ keta = -0.005531984945704 lketa = -2.22342109475967e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.117939716445715 lags = 8.35623612841368e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.276398142045985+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.86082819697777e-8
+ nfactor = {1.5717742327426+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.47710253034928e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.15964838675 leta0 = -3.18890874427738e-7
+ etab = -0.139629721319197 letab = 2.78778813026474e-7
+ dsub = 0.86055995 ldsub = -1.20336179029335e-6
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.464241322871765 lpclm = -1.2258811017163e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -1.9453378406665e-05 lpdiblc2 = 7.06261097247162e-10
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800440951.502645 lpscbe1 = -1.76545208253947
+ pscbe2 = 8.29037304530805e-09 lpscbe2 = 1.30287299130047e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.9206340066811 lbeta0 = 8.47971588955986e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.31276341430735e-10 lagidl = -6.2669437444031e-17
+ bgidl = 918242083.1476 lbgidl = 327.33686971321
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.466354778793985 lkt1 = 4.18806003875746e-9
+ kt2 = -0.0057096990819635 lkt2 = -7.6529722443776e-8
+ at = 106881.333549731 lat = -0.0518986434486551
+ ute = -0.176067522322505 lute = -1.1821437140863e-7
+ ua1 = 2.34105191043975e-09 lua1 = -1.38852507456877e-15
+ ub1 = -1.02898979966153e-18 lub1 = 8.34390287342497e-25
+ uc1 = -2.41157429708828e-10 luc1 = 4.50184982244457e-16 puc1 = -7.52316384526264e-37
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.4 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0498109691552+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.77836999732568e-8
+ k1 = 0.35649664992175 lk1 = 1.62033872934792e-7
+ k2 = 0.052734565514376 lk2 = -6.45665159115012e-08 wk2 = 5.29395592033938e-23 pk2 = 5.04870979341448e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 35558.5059375 lvsat = 0.0358247304098353
+ ua = -7.5086450953842e-10 lua = -2.49244108346923e-16
+ ub = 1.01442260279428e-18 lub = 1.72543647137309e-25
+ uc = -4.2898643670165e-11 luc = 7.33188681166072e-18
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0096799593629 lu0 = -9.4788465640171e-10
+ a0 = 1.25970100231 la0 = -3.56125474451623e-7
+ keta = -0.006915534800507 lketa = -1.94619464463827e-8
+ a1 = 0.0
+ a2 = 0.6996267 la2 = 2.011212935289e-7
+ ags = 0.41242641448365 lags = 2.45550897921723e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.2631120370841+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.986475016185e-9
+ nfactor = {1.3371515750889+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.22410908653493e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.4908273035 leta0 = 9.84488731823965e-07 weta0 = -1.91905902112302e-22 peta0 = -2.16147888030557e-28
+ etab = 7.4649203674932 letab = -1.49587091500798e-05 wetab = -1.00585162486448e-21 petab = -1.95479732313767e-27
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.18780596974631 lpclm = 4.31314529252497e-7
+ pdiblc1 = 0.40816306053883 lpdiblc1 = -3.63939237826515e-8
+ pdiblc2 = 0.00023567653097224 lpdiblc2 = 1.95048878537641e-10
+ pdiblcb = -0.0493458950609527 lpdiblcb = 4.8782673348168e-8
+ drout = 0.40383213350502 ldrout = 3.12918707635586e-7
+ pscbe1 = 799118096.99471 lpscbe1 = 0.885195149208812
+ pscbe2 = 8.9456890419886e-09 lpscbe2 = -1.02052966762473e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -4.4813805135721e-05 lalpha0 = 8.97951005793136e-11 walpha0 = -1.59706862414257e-26 palpha0 = -4.37929009805622e-32
+ alpha1 = 2.003733e-10 lalpha1 = -2.011212935289e-16
+ beta0 = -13.670975394132 lbeta0 = 4.37286041690793e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 804510852.3414 lbgidl = 555.223890010209
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.45639520260806 lkt1 = -1.57682714309942e-8
+ kt2 = -0.040433002663921 lkt2 = -6.95349318758958e-9
+ at = 71096.512835428 lat = 0.0198045827156774
+ ute = -0.16633222632958 lute = -1.37721305254422e-7
+ ua1 = 1.4213951221082e-09 lua1 = 4.5422158088517e-16
+ ub1 = -2.32019645259997e-20 lub1 = -1.18093998891712e-24
+ uc1 = -2.1485789154501e-11 luc1 = 1.00216669016128e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.5 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.047063872301+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.50263482064995e-8
+ k1 = 0.56078790140908 lk1 = -4.301999779434e-8
+ k2 = -0.035753754167148 lk2 = 2.4252130667394e-08 wk2 = -2.64697796016969e-23 pk2 = 1.26217744835362e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 59266.2926766 lvsat = 0.0120284425028382
+ ua = -6.690174615183e-10 lua = -3.31396691397302e-16
+ ub = 1.01232240728044e-18 lub = 1.74651682681002e-25
+ uc = -5.8251570637308e-11 luc = 2.27421262551721e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.010390362905 lu0 = -1.66094013492437e-9
+ a0 = 0.8997619234 la0 = 5.15725703994801e-9
+ keta = -0.04253162444915 lketa = 1.62870980649187e-8
+ a1 = 0.0
+ a2 = 1.0007466 la2 = -1.011226870578e-7
+ ags = 0.47384338151394 lags = 1.83904661353508e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.26366137734554+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.53786596482088e-9
+ nfactor = {1.6179752970192+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.05388717692274e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = -14.9317815030846 letab = 7.52159960858082e-6
+ dsub = 0.22035862074374 ldsub = 3.97893605250237e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.61188613603502 lpclm = 5.65127170303116e-9
+ pdiblc1 = 0.707442757014598 lpdiblc1 = -3.36790831365364e-7
+ pdiblc2 = 0.00043
+ pdiblcb = 0.225184990121906 lpdiblcb = -2.26773035629078e-07 wpdiblcb = -4.96308367531817e-24 ppdiblcb = 6.7053176943786e-29
+ drout = 0.42905069298996 ldrout = 2.87606007268088e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 8.7234119240386e-09 lpscbe2 = 2.12901581755065e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 8.9627910271442e-05 lalpha0 = -4.51484857514643e-11
+ alpha1 = -1.007466e-10 lalpha1 = 1.011226870578e-16
+ beta0 = 50.5387402081872 lbeta0 = -2.07208063015834e-05 pbeta0 = -2.58493941422821e-26
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1701651032.0586 lbgidl = -345.265313997875
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.43547823230078 lkt1 = -3.67633247884312e-8
+ kt2 = -0.03947483089291 lkt2 = -7.91524181382177e-9
+ at = 106773.04766704 lat = -0.0160051326204611
+ ute = -0.23633461306978 lute = -6.74575996045206e-8
+ ua1 = 3.3034787359484e-09 lua1 = -1.4348878510855e-15
+ ub1 = -2.8245204414334e-18 lub1 = 1.63083580986457e-24
+ uc1 = -4.7590230527604e-11 luc1 = 3.62235561543616e-17 wuc1 = 2.46519032881566e-32 puc1 = -1.17549435082229e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.6 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.9916153578692+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -2.90489831377424e-9
+ k1 = 0.12097473666744 lk1 = 1.78528407120461e-7
+ k2 = 0.13042219941516 lk2 = -5.94561809584828e-08 pk2 = 1.26217744835362e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 53286.5139988 lvsat = 0.0150406543555425
+ ua = -5.633691056756e-10 lua = -3.84615254631013e-16
+ ub = 9.095841041608e-19 lub = 2.26404356326368e-25
+ uc = -2.6502209151207e-11 luc = 6.74892514569395e-18
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.01013907332112 lu0 = -1.53435727896774e-9
+ a0 = 1.16838856412924 la0 = -1.30158846574514e-7
+ keta = 0.062618329972472 lketa = -3.66804039257482e-08 wketa = 2.64697796016969e-23 pketa = -1.26217744835362e-29
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.38868016400772 lags = 6.18386234509771e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.19808734652972+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -3.04939373001245e-8
+ nfactor = {1.3353523605304+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 1.8290537143554e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.985613787305066 leta0 = -2.49657019920543e-7
+ etab = 0.0049827448348032 letab = -2.54145631636992e-09 wetab = -8.27180612553028e-25 petab = -8.38164711797325e-31
+ dsub = 0.1803345523228 ldsub = 5.9950804582909e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.47136627312296 lpclm = 7.6435763807312e-8
+ pdiblc1 = -0.350328483720116 lpdiblc1 = 1.96043449043656e-07 wpdiblc1 = -1.05879118406788e-22 ppdiblc1 = 2.52435489670724e-29
+ pdiblc2 = -0.009375225574176 lpdiblc2 = 4.9392156941564e-09 wpdiblc2 = 1.65436122510606e-24 ppdiblc2 = 2.95822839457879e-30
+ pdiblcb = -0.3772398 lpdiblcb = 7.66882111734e-08 ppdiblcb = -1.0097419586829e-28
+ drout = 1.53912143474972 ldrout = -2.71573257690781e-7
+ pscbe1 = 800003592.85928 lpscbe1 = -0.00180984178371091
+ pscbe2 = 9.41458269657e-09 lpscbe2 = -1.35263945004496e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -8.05815789449e-09 lalpha0 = 4.10953335066513e-15 walpha0 = -2.16936748935778e-30 palpha0 = 1.59867231711831e-36
+ alpha1 = 2.014932e-10 lalpha1 = -5.11254741156e-17
+ beta0 = 3.1239804714936 lbeta0 = 3.16357286486052e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 461943346.4792 lbgidl = 279.216357582093
+ cgidl = 537.508136688744 lcgidl = -0.000119640686218631
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.45726682992 lkt1 = -2.57876891439086e-8
+ kt2 = 0.012581039504 lkt2 = -3.41375015764684e-08 pkt2 = 2.52435489670724e-29
+ at = 62820.816 lat = 0.006135056893872
+ ute = -0.377608257 lute = 3.706596873381e-9
+ ua1 = 7.801034662e-10 lua1 = -1.63780456329325e-16
+ ub1 = 4.3356282096e-19 lub1 = -1.03682461506437e-26
+ uc1 = 1.045095422e-11 luc1 = 6.98629603789674e-18
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.7 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.823745841514286+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -4.54989343070559e-8
+ k1 = 0.305901478718572 lk1 = 1.31606390079601e-7
+ k2 = 0.0785605101573427 lk2 = -4.62971589580291e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 185876.616708571 lvsat = -0.0186018301753159
+ ua = -1.56158896686571e-09 lua = -1.31333934591662e-16
+ ub = 1.34942793818e-18 lub = 1.14801460789174e-25
+ uc = -5.79026830087713e-14 luc = 3.91319325986106e-20
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00567692584828571 lu0 = -4.02163214243079e-10
+ a0 = 0.980575535395571 la0 = -8.25044833548346e-8
+ keta = -0.235670100842443 lketa = 3.90052144902125e-8
+ a1 = 0.0
+ a2 = 0.874270679313286 la2 = -1.88449222741979e-8
+ ags = 4.14427143508 lags = -5.31773173581553e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0964041543790002+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -5.62943186941032e-8
+ nfactor = {0.75577407357143+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 3.299635089205e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.442285423697377 leta0 = 1.1264813058474e-07 weta0 = 1.65436122510606e-22 peta0 = -5.04870979341448e-29
+ etab = 0.131953317290431 letab = -3.47580805772538e-08 wetab = -7.94093388050907e-23 petab = 3.15544362088405e-30
+ dsub = 0.767247788263 ldsub = -8.89684515119057e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.13020133376457 lpclm = -9.0732432634466e-8
+ pdiblc1 = 1.04097151158557 lpdiblc1 = -1.56975272665242e-7
+ pdiblc2 = 0.0256223919961886 lpdiblc2 = -3.94083480482491e-9
+ pdiblcb = -0.075
+ drout = -0.79349313840957 ldrout = 3.20288035800646e-7
+ pscbe1 = 799987168.359714 lpscbe1 = 0.00235759576469263
+ pscbe2 = 8.04351632122143e-09 lpscbe2 = 2.12620839611823e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.92362781946071e-08 lalpha0 = -5.35329580152975e-15
+ alpha1 = -2.62475714285714e-10 lalpha1 = 6.65987504128571e-17
+ beta0 = 33.93082679872 lbeta0 = -4.65314067428562e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.58634322552858e-11 lagidl = 8.66157374356958e-18
+ bgidl = 3038480410.20429 lbgidl = -374.536121208064
+ cgidl = -548.243345316942 lcgidl = 0.000155850294565118 wcgidl = 2.16840434497101e-19 pcgidl = -5.16987882845642e-26
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.5589
+ kt2 = -0.12196
+ at = 215613.1 lat = -0.0326333877023
+ ute = -0.5283597 lute = 4.19572127601e-8
+ ua1 = 1.3462e-10
+ ub1 = 3.927e-19
+ uc1 = 3.7985e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.8 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.768589483199999+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -5.56329774892145e-8
+ k1 = -0.341733350206669 lk1 = 2.50598280102522e-7
+ k2 = 0.391488894107334 lk2 = -1.03792429726313e-7
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 235927.59462 lvsat = -0.0277978464999165
+ ua = -9.78084494193332e-10 lua = -2.38542961869176e-16
+ ub = 6.55962328626665e-19 lub = 2.42213977629237e-25
+ uc = 2.78157227447333e-13 luc = -2.26133629292209e-20
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00626552286666666 lu0 = -5.10307910221268e-10
+ a0 = -0.887083380342002 la0 = 2.60646092210377e-7
+ keta = -0.0965098958122733 lketa = 1.34368925394044e-8
+ a1 = 0.0
+ a2 = -0.395622701731002 la2 = 2.14476398305212e-7
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.265663331828667+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -2.51958222437436e-8
+ nfactor = {-0.706147247333334+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 5.98566698974295e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.674395175969667 leta0 = 1.55294351698985e-7
+ etab = -0.260717309417333 letab = 3.73884716796439e-08 petab = -5.04870979341448e-29
+ dsub = 0.400990212300667 ldsub = -2.16748483076184e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.22551412948367 lpclm = -2.91977538530323e-7
+ pdiblc1 = 1.04292508576367 lpdiblc1 = -1.57334208709706e-7
+ pdiblc2 = 0.0233579651270267 lpdiblc2 = -3.52478486287319e-09 wpdiblc2 = 2.64697796016969e-23
+ pdiblcb = -0.443529158579553 lpdiblcb = 6.77109678932971e-8
+ drout = 0.692138700041332 ldrout = 4.73284412265458e-8
+ pscbe1 = 872184766.462333 lpscbe1 = -13.2627236964239
+ pscbe2 = 1.020073986908e-08 lpscbe2 = -1.83732314506877e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 14.8988522472 lbeta0 = -1.1563388940112e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.79651991404333e-10 lagidl = -1.22451395945624e-17
+ bgidl = 765071891.163333 lbgidl = 43.1640462208874
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = 0.112913210000001 lkt1 = -1.2343425651293e-7
+ kt2 = -0.12196
+ at = 38000.0
+ ute = -0.3
+ ua1 = 1.3462e-10
+ ub1 = 3.927e-19
+ uc1 = 3.7985e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.9 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.06314409338213+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = 9.36017216978696e-8
+ k1 = 0.444350182392039 wk1 = -6.93527698187977e-8
+ k2 = 0.0178871871725287 wk2 = 2.73987109091685e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 160312.5
+ ua = -6.8337407612387e-10 wua = 6.39537790816786e-16
+ ub = 9.25039483898675e-19 wub = 3.70150575149886e-26
+ uc = -7.49057583753778e-11 wuc = 5.87448458332351e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.01020196685651 wu0 = 1.60738981397932e-9
+ a0 = 1.1897275623139 wa0 = -1.29068627637358e-7
+ keta = 0.0302574562880444 wketa = -1.76663841434654e-7
+ a1 = 0.0
+ a2 = 1.22518058161453 wa2 = -1.58663202789754e-6
+ ags = 0.359147361700281 wags = -5.23581326226342e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.302788080551888+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = 1.34145079428299e-7
+ nfactor = {0.83484118121044+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor = 3.94614376162484e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.566314698625682 wpclm = 3.99214303892371e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00999213432141191 wpdiblc2 = -4.94161199728854e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.01282218825559e-08 wpscbe2 = -5.28777845969291e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 0.358552501150871 wbeta0 = 3.01454253428577e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 272285627.87766 wbgidl = 6389.23127781209
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.479805285058396 wkt1 = 2.20089684104728e-7
+ kt2 = 0.100495825740763 wkt2 = -7.59753679266766e-7
+ at = 93163.69449 wat = -0.0159147506334585
+ ute = -0.779269923657029 wute = 3.09149141458192e-6
+ ua1 = 7.3269798691391e-10 wua1 = 6.17062449480527e-15
+ ub1 = -7.91678035807245e-20 wub1 = -3.3867855454828e-24
+ uc1 = -6.63211962253626e-10 wuc1 = 3.89930240657708e-15
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.10 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.06314409338213+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = 9.3601721697873e-8
+ k1 = 0.444350182392038 wk1 = -6.93527698187977e-8
+ k2 = 0.0178871871725287 wk2 = 2.73987109091686e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 160312.5
+ ua = -6.8337407612387e-10 wua = 6.3953779081679e-16
+ ub = 9.25039483898675e-19 wub = 3.70150575149857e-26
+ uc = -7.49057583753778e-11 wuc = 5.87448458332353e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.01020196685651 wu0 = 1.60738981397932e-9
+ a0 = 1.1897275623139 wa0 = -1.29068627637358e-7
+ keta = 0.0302574562880444 wketa = -1.76663841434654e-7
+ a1 = 0.0
+ a2 = 1.22518058161453 wa2 = -1.58663202789754e-6
+ ags = 0.359147361700281 wags = -5.23581326226341e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.302788080551888+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = 1.34145079428296e-7
+ nfactor = {0.834841181210439+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor = 3.94614376162485e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.566314698625682 wpclm = 3.99214303892371e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00999213432141191 wpdiblc2 = -4.94161199728854e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.01282218825559e-08 wpscbe2 = -5.28777845969296e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 0.358552501150864 wbeta0 = 3.01454253428577e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 272285627.87766 wbgidl = 6389.23127781208
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.479805285058396 wkt1 = 2.20089684104726e-7
+ kt2 = 0.100495825740763 wkt2 = -7.59753679266766e-7
+ at = 93163.69449 wat = -0.0159147506334585
+ ute = -0.779269923657029 wute = 3.09149141458192e-6
+ ua1 = 7.3269798691391e-10 wua1 = 6.17062449480527e-15
+ ub1 = -7.91678035807233e-20 wub1 = -3.3867855454828e-24
+ uc1 = -6.63211962253626e-10 wuc1 = 3.89930240657708e-15
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.11 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.06335251172813+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.66812479366851e-09 wvth0 = 6.5305436769891e-08 pvth0 = 2.26475909455482e-13
+ k1 = 0.417748010567478 lk1 = 2.12916680503905e-07 wk1 = 1.43164418789115e-07 pk1 = -1.70093083552838e-12
+ k2 = 0.0269405997198028 lk2 = -7.24610967672312e-08 wk2 = -4.28399357209938e-08 pk2 = 5.62171373909167e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 275661.253709246 lvsat = -0.923220626571569 wvsat = -0.0588729279351927 pvsat = 4.71203196121522e-7
+ ua = -4.20510795511145e-10 lua = -2.10388751352833e-15 wua = -1.47383008238857e-15 pua = 1.69148321879135e-20
+ ub = 6.67240447557752e-19 lub = 2.06335465453005e-24 wub = 1.816276320814e-24 pub = -1.4240732088688e-29
+ uc = -9.31136720706297e-11 luc = 1.4573127970384e-16 wuc = 1.40105753724712e-16 puc = -6.51190983400975e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0107251683542974 lu0 = -4.18756509349062e-09 wu0 = -4.63170472352818e-09 pu0 = 4.99360468399685e-14
+ a0 = 1.3569273789059 la0 = -1.33822268965135e-06 wa0 = -8.88556703110967e-07 pa0 = 6.07873977277466e-12
+ keta = 0.0732581702080277 lketa = -3.4416623302493e-07 wketa = -3.64877070025924e-07 pketa = 1.50640842871249e-12
+ a1 = 0.0
+ a2 = 1.65075796300686 la2 = -3.40620773150333e-06 wa2 = -3.1747447801351e-06 pa2 = 1.27108304428047e-11
+ ags = 0.426359865346333 lags = -5.37950933444531e-07 wags = -1.29150642747056e-06 pags = 6.14626747435668e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.346056350025297+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 3.46307676237215e-07 wvoff = 3.36622016213953e-07 pvoff = -1.62057134069027e-12
+ nfactor = {0.284490795780847+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.40485754142555e-06 wnfactor = 6.83899507906969e-06 pnfactor = -2.31536095535267e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.55057608604438 lpclm = 7.87776534710884e-06 wpclm = 7.87124067497892e-06 ppclm = -3.1047261759917e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0197120134227004 lpdiblc2 = -7.77953171189932e-08 wpdiblc2 = -9.80031626683832e-08 ppdiblc2 = 3.88877716994365e-13
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.37808850517652e-08 lpscbe2 = -2.92349407452849e-14 wpscbe2 = -2.5617302509252e-14 ppscbe2 = 1.6271208250975e-19
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -3.73706636083686 lbeta0 = 3.27802398411136e-05 wbeta0 = 4.91425938513549e-05 pbeta0 = -1.52048264498019e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 4.50284505267915e-11 lagidl = 4.3997760457985e-16 wagidl = 2.7653065255392e-16 pagidl = -2.21327750935734e-21
+ bgidl = 769023572.773279 lbgidl = -3975.75788191325 wbgidl = 4171.22166501484 pbgidl = 0.0177523567322626
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.488169860817833 lkt1 = 6.69478310368075e-08 wkt1 = 3.97179258479388e-07 pkt1 = -1.41737767037846e-12
+ kt2 = 0.158957377229222 lkt2 = -4.67910648879379e-07 wkt2 = -1.04934954446856e-06 pkt2 = 2.31784798297911e-12
+ at = 93422.3916636896 lat = -0.00207054310606614 wat = -0.0389765679911629 pat = 1.84580628625831e-7
+ ute = -1.35347560345259 lute = 4.59578894816713e-06 wute = 6.18582530758937e-06 pute = -2.47662222924822e-11
+ ua1 = -5.89938272296149e-11 lua1 = 6.33648989869039e-15 wua1 = 9.03545033057439e-15 pua1 = -2.29293010809979e-20
+ ub1 = 4.04631367150108e-19 lub1 = -3.872199388151e-24 wub1 = -4.96068909177793e-24 pub1 = 1.25971037522993e-29
+ uc1 = -1.2022990983295e-09 luc1 = 4.31470950088599e-15 wuc1 = 7.83101570920264e-15 puc1 = -3.14683835067632e-20
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.12 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0749937278555+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.82764459629791e-08 wvth0 = 1.3863101809275e-07 pvth0 = -6.71001402310366e-14
+ k1 = 0.516059375208804 lk1 = -1.80695774385606e-07 wk1 = -6.44749386006914e-07 pk1 = 1.45366566588903e-12
+ k2 = -0.00611712770355521 lk2 = 5.98932174226719e-08 wk2 = 2.18303604492662e-07 pk2 = -4.83377635781072e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 36689.4747690071 lvsat = 0.0335585708401731 wvsat = 0.117745855870385 pvsat = -2.35931257020734e-7
+ ua = -1.29357249485663e-09 lua = 1.39161842317726e-15 wua = 7.45239814093409e-15 pua = -1.88234023153348e-20
+ ub = 1.41835709246261e-18 lub = -9.43915843524823e-25 wub = -4.56388510644073e-24 pub = 1.13037307629389e-29
+ uc = -6.20613235831544e-11 luc = 2.14059673370353e-17 wuc = -1.30622422772042e-16 puc = 4.32732350868903e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0087793886415943 lu0 = 3.60281735298934e-09 wu0 = 2.53494509076221e-08 pu0 = -7.0100495338604e-14
+ a0 = 1.10904077867381 la0 = -3.45750928044309e-07 wa0 = 2.35883265220201e-07 pa0 = 1.57678236504821e-12
+ keta = -0.00906547104953757 lketa = -1.45643538418543e-08 wketa = 2.48419344826442e-08 pketa = -5.39224103656099e-14
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.101674165059227 lags = 1.57615633921322e-06 wags = 1.54398050409933e-06 pags = -5.20626512463842e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.285589615559577+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.04215016054573e-07 wvoff = 6.4620031355402e-08 pvoff = -5.31548017846579e-13
+ nfactor = {1.07056739948853+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.25761670263318e-06 wnfactor = 3.52370065936947e-06 pnfactor = -9.88005588065708e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.15964839156303 leta0 = -3.18890893697823e-07 weta0 = -3.38376779056965e-14 peta0 = 1.35477027705489e-19
+ etab = -0.139629721293998 letab = 2.78778812925584e-07 wetab = -1.771607525665e-16 petab = 7.09303336296386e-22
+ dsub = 0.86055995 ldsub = -1.20336179029335e-6
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.02576092559086 lpclm = -2.43720016549656e-06 wpclm = -3.94772549588753e-06 ppclm = 1.62727231242646e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000473902657424833 lpdiblc2 = -7.71058190404067e-10 wpdiblc2 = -3.46850616037412e-09 ppdiblc2 = 1.03861930895843e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 772447464.564305 lpscbe1 = 110.312995357559 wpscbe1 = 196.806311961584 ppscbe1 = -0.000787959925808886
+ pscbe2 = 5.30884827750386e-09 lpscbe2 = 4.6848324650386e-15 wpscbe2 = 2.0961407732668e-14 ppscbe2 = -2.37766367832636e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 0.942988286908729 lbeta0 = 1.40425506061312e-05 wbeta0 = 2.09341363484798e-05 pbeta0 = -3.91091323146611e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.09943098946417e-10 lagidl = -2.202966154812e-16 wagidl = -5.5306130510784e-16 pagidl = 1.10818718806765e-21
+ bgidl = -867722965.588937 lbgidl = 2577.33824636332 wbgidl = 12556.1061867119 pbgidl = -0.0158184821284452
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.481232740769185 lkt1 = 3.9173454573072e-08 wkt1 = 1.04598502940819e-07 pkt1 = -2.45962444263741e-13
+ kt2 = 0.125981455220248 lkt2 = -3.35883861726626e-07 wkt2 = -9.25845731661438e-07 pkt2 = 1.82337169201743e-12
+ at = 101232.224651025 lat = -0.0333390291619506 wat = 0.0397156771027678 pat = -1.30482109900827e-7
+ ute = -0.326488745051784 lute = 4.84007772621514e-07 wute = 1.0575262078393e-06 pute = -4.23388195294257e-12
+ ua1 = 1.02449598397185e-09 lua1 = 1.99848598641932e-15 wua1 = 9.25595717854076e-15 pua1 = -2.38121516249269e-20
+ ub1 = -3.5158941581117e-19 lub1 = -8.44493284123087e-25 wub1 = -4.76241747091393e-24 pub1 = 1.18032771208826e-29
+ uc1 = 9.60217797845031e-11 luc1 = -8.83420643408035e-16 wuc1 = -2.37051557159247e-15 puc1 = 9.37582393268843e-21
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.13 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.06828927846333+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.48425194690553e-08 wvth0 = 1.29910500761461e-07 pvth0 = -4.96265518772558e-14
+ k1 = 0.326566465937276 lk1 = 1.98997421187763e-07 wk1 = 2.10422129236375e-07 pk1 = -2.59869719863941e-13
+ k2 = 0.061150688798939 lk2 = -7.48935263413203e-08 wk2 = -5.9168984138961e-08 pk2 = 7.26033466555361e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -73722.0355817526 lvsat = 0.254793757709832 wvsat = 0.76828943793039 pvsat = -1.53944690033257e-6
+ ua = -5.95014570620854e-10 lua = -8.10514202546046e-18 wua = -1.09569242893409e-15 pua = -1.69531115350113e-21
+ ub = 9.0356074292101e-19 lub = 8.75985903312195e-26 wub = 7.79406789404933e-25 pub = 5.9720046260036e-31
+ uc = -5.36704484158479e-11 luc = 4.59289386542234e-18 wuc = 7.57304429361613e-17 puc = 1.92563042048074e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0103933458297272 lu0 = 3.68878074540344e-10 wu0 = -5.01541518742586e-09 pu0 = -9.25741110337503e-15
+ a0 = 0.076704027381334 la0 = 1.72277628763321e-06 wa0 = 8.31698002504109e-06 pa0 = -1.4615577888798e-11
+ keta = -0.0716996616387246 lketa = 1.10937840769989e-07 wketa = 4.55460411372289e-07 pketa = -9.16766862919129e-13
+ a1 = 0.0
+ a2 = 0.44716615982987 la2 = 7.06984809065615e-07 wa2 = 1.77490671084147e-06 pa2 = -3.55643914843452e-12
+ ags = 2.35210280502763 lags = -3.34055755038984e-06 wags = -1.36367633536602e-05 pags = 2.52118923077016e-11
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.236166299421282+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 5.18388653883806e-09 wvoff = -1.8944018171743e-07 pvoff = -2.24791849255107e-14
+ nfactor = {1.45533858469696+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.8663798138194e-07 wnfactor = -8.30905757970197e-07 pnfactor = -1.15458730022181e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.490827313126059 leta0 = 9.84488741485959e-07 weta0 = 6.76753550404607e-14 peta0 = -6.79279866932551e-20
+ etab = 26.2401722495116 letab = -5.25793009294427e-05 wetab = -0.000131998135394453 petab = 2.64489019828688e-10
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.49847984671121 lpclm = 2.62070436991058e-06 wpclm = 1.18553181024263e-05 ppclm = -1.53923568341155e-11
+ pdiblc1 = 0.431783268677147 lpdiblc1 = -8.37225142962666e-08 wpdiblc1 = -1.6606027186633e-07 ppdiblc1 = 3.32740446727535e-13
+ pdiblc2 = -0.000253088986934233 lpdiblc2 = 6.85638958122458e-10 wpdiblc2 = 3.43623283533935e-09 ppdiblc2 = -3.44906029251367e-15
+ pdiblcb = -0.0493912705764652 lpdiblcb = 4.88735937659923e-08 wpdiblcb = 3.19009485350353e-10 ppdiblcb = -6.3920983310956e-16
+ drout = 0.646962994413163 ldrout = -1.74250621684469e-07 wdrout = -1.70931503334233e-06 pdrout = 3.42501093970412e-12
+ pscbe1 = 855105070.871389 lpscbe1 = -55.3107781009521 wpscbe1 = -393.612623923167 ppscbe1 = 0.000395081979848274
+ pscbe2 = 1.99688464655647e-09 lpscbe2 = 1.13211232871677e-14 wpscbe2 = 4.88530981731477e-14 ppscbe2 = -7.96641373446371e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -0.000157530460836959 lalpha0 = 3.15649183257523e-10 walpha0 = 7.92446805718298e-10 palpha0 = -1.58785181536234e-15
+ alpha1 = 4.5283384017013e-10 lalpha1 = -7.06984809065615e-16 walpha1 = -1.77490671084148e-15 palpha1 = 3.55643914843452e-21
+ beta0 = -67.0014310998223 lbeta0 = 0.000150185025897164 wbeta0 = 0.000374936153033959 pbeta0 = -7.48434655213907e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = -964031701.888411 lbgidl = 2770.31523947488 wbgidl = 12433.6185203275 pbgidl = -0.0155730495492178
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.456037107736268 lkt1 = -1.13118667908732e-08 wkt1 = -2.51756171730397e-09 pkt1 = -3.13304506781357e-14
+ kt2 = -0.0368006820787488 lkt2 = -9.71192141009485e-09 wkt2 = -2.55367836027181e-08 pkt2 = 1.93929425968899e-14
+ at = -86801.0111937397 lat = 0.343429370596988 wat = 1.11008783723494 pat = -2.27522212943894e-6
+ ute = 0.295079810589718 lute = -7.61449654079699e-07 wute = -3.24392604182502e-06 pute = 4.38507986763407e-12
+ ua1 = 2.2482129589609e-09 lua1 = -4.53516099026409e-16 wua1 = -5.81288674374355e-15 pua1 = 6.38178821400367e-21
+ ub1 = -4.39577686940451e-19 lub1 = -6.68188281648402e-25 wub1 = 2.92730128616082e-24 pub1 = -3.60486611338701e-30
+ uc1 = -6.78683826633964e-10 luc1 = 6.6888254545766e-16 wuc1 = 4.62038624447242e-15 puc1 = -4.63207673592072e-21
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.14 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.04174419892901+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.19834715282742e-09 wvth0 = -3.73996029679366e-08 pvth0 = 1.1830812046937e-13
+ k1 = 0.590051086441485 lk1 = -6.54707874047882e-08 wk1 = -2.05732838326371e-07 pk1 = 1.57838754192719e-13
+ k2 = -0.0485524385121944 lk2 = 3.52191227440656e-08 wk2 = 8.99802825370504e-08 pk2 = -7.71026942329772e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 269329.624477245 lvsat = -0.0895385141961657 wvsat = -1.47683601193054 pvsat = 7.14059602832683e-7
+ ua = 4.46435783152769e-11 lua = -6.50151134831569e-16 wua = -5.01734555433145e-15 pua = 2.24098150301335e-21
+ ub = 6.43508606088843e-19 lub = 3.4862150179018e-25 wub = 2.5929204237018e-24 pub = -1.22308301809334e-30
+ uc = -8.22977402087657e-11 luc = 3.33270513386032e-17 wuc = 1.69054964841836e-16 puc = -7.44165981411415e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.014062964865402 lu0 = -3.31443964899469e-09 wu0 = -2.58199790801936e-08 pu0 = 1.16248162264043e-14
+ a0 = 2.66327816297539 la0 = -8.73453529209019e-07 wa0 = -1.23982813559338e-05 pa0 = 6.17701356291206e-12
+ keta = 0.0786750059549647 lketa = -3.99981754578274e-08 wketa = -8.52134997246587e-07 pketa = 3.95709799360122e-13
+ a1 = 0.0
+ a2 = 1.51208289337108 la2 = -3.61907258641901e-07 wa2 = -3.59491514194466e-06 pa2 = 1.83342824932807e-12
+ ags = -2.68420466825445 lags = 1.71455045869e-06 wags = 2.22024426982389e-05 pags = -1.07611015003892e-11
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.245048037871199+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.40987805183888e-08 wvoff = -1.30859821189938e-07 pvoff = -8.12782259388541e-14
+ nfactor = {2.29568131661117+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.56841749950507e-07 wnfactor = -4.76456622227322e-06 pnfactor = 2.79375751859445e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = -52.4822060798878 letab = 2.64369480382604e-05 wetab = 0.000263995714068429 petab = -1.32983074674239e-10
+ dsub = 0.201690073605044 ldsub = 5.8527597350188e-08 wdsub = 1.31247954931104e-07 pdsub = -1.31737903546862e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.60741490517706 lpclm = -4.96784687086484e-07 wpclm = -6.99899751460254e-06 ppclm = 3.53234194311168e-12
+ pdiblc1 = 0.611162480983884 lpdiblc1 = -2.63771349202545e-07 wpdiblc1 = 6.76891952831219e-07 ppdiblc1 = -5.13358518624807e-13
+ pdiblc2 = 0.00043
+ pdiblcb = 0.225275741152931 lpdiblcb = -2.26818749918189e-07 wpdiblcb = -6.38018970700609e-10 ppdiblcb = 3.21391210167792e-16
+ drout = -0.0572110288263259 ldrout = 5.32552083183772e-07 wdrout = 3.41863006668465e-06 pdrout = -1.72207677938126e-12
+ pscbe1 = 800000000.0
+ pscbe2 = -3.20549135275597e-09 lpscbe2 = 1.65429197560856e-14 wpscbe2 = 8.38653457078619e-14 ppscbe2 = -1.14807085599398e-19
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.000315061221673918 lalpha0 = -1.58706684004168e-10 walpha0 = -1.5848936114366e-09 palpha0 = 7.98363213569792e-16
+ alpha1 = -6.0566768034026e-10 lalpha1 = 3.55468097620841e-16 walpha1 = 3.54981342168295e-15 palpha1 = -1.78815816434462e-21
+ beta0 = 156.416791355518 lbeta0 = -7.4067216782602e-05 wbeta0 = -0.000744368460059441 pbeta0 = 3.75048322000171e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 3096320386.42579 lbgidl = -1305.194143185 wbgidl = -9805.12833729631 pbgidl = 0.0067487145504255
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.425846559740641 lkt1 = -4.16151161021678e-08 wkt1 = -6.77148209066575e-08 pkt1 = 3.41101898797714e-14
+ kt2 = -0.037699927262087 lkt2 = -8.80931934448708e-09 wkt2 = -1.24783396380341e-08 pkt2 = 6.28575146088592e-15
+ at = 426608.654278905 lat = -0.171896853156867 wat = -2.24858254743059 pat = 1.09598617177255e-6
+ ute = -0.424183533321056 lute = -3.95013001061072e-08 wute = 1.3206590976698e-06 pute = -1.9654486818649e-13
+ ua1 = 3.12247212476655e-09 lua1 = -1.33103887429802e-15 wua1 = 1.27255470766576e-15 pua1 = -7.30103190343741e-22
+ ub1 = -2.54823985395907e-18 lub1 = 1.4483455212397e-24 wub1 = -1.94237193841447e-24 pub1 = 1.28298560133563e-30
+ uc1 = -4.91711889222574e-11 luc1 = 3.70199370693755e-17 wuc1 = 1.11148208046314e-17 puc1 = -5.5989020283794e-24
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.15 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.05636724546566+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.5564458253876e-08 wvth0 = 4.55233755568939e-07 pvth0 = -1.29847559126492e-13
+ k1 = 0.0868475978712553 lk1 = 1.88009415503159e-07 wk1 = 2.39928535486563e-07 pk1 = -6.66555866221941e-14
+ k2 = 0.153012015749869 lk2 = -6.63155444947266e-08 wk2 = -1.58816172151626e-07 pk2 = 4.8224290276714e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 22113.7369484139 lvsat = 0.0349922864763949 wvsat = 0.219158095538455 pvsat = -1.40268596904995e-7
+ ua = -3.33373096616676e-10 lua = -4.59731661118072e-16 wua = -1.61697134795934e-15 pua = 5.28100802914905e-22
+ ub = 8.87135225143802e-19 lub = 2.25898734093767e-25 wub = 1.57825321894989e-25 pub = 3.55474282511048e-33
+ uc = -3.25561055784428e-11 luc = 8.27054850136674e-18 wuc = 4.25615083775039e-17 puc = -1.0697669835994e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0111967335579596 lu0 = -1.87062435380277e-09 wu0 = -7.43580858573647e-09 pu0 = 2.36410287072001e-15
+ a0 = 1.24139616885342 la0 = -1.57204646663976e-07 wa0 = -5.13275015097785e-07 pa0 = 1.90143663823715e-13
+ keta = 0.0329539760785183 lketa = -1.69669839150754e-08 wketa = 2.08553228808248e-07 pketa = -1.38593862815159e-13
+ a1 = 0.0
+ a2 = 0.787169573938368 la2 = 3.25550249589605e-09 wa2 = 9.02034405234174e-08 pa2 = -2.28875895743286e-14
+ ags = -0.0816142642123276 lags = 4.03539786690653e-07 wags = -2.1588059894435e-06 pags = 1.51046338480315e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.163992098518546+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.67317709795409e-08 wvoff = -2.39704329484745e-07 pvoff = -2.64496552419865e-14
+ nfactor = {1.51806926236015+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 3.48671029735201e-08 wnfactor = -1.28457879010814e-06 pnfactor = 1.04077300942763e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 2.05660100940677 leta0 = -7.89148626271501e-07 weta0 = -7.52950305205238e-06 peta0 = 3.79285916091951e-12
+ etab = 0.0140625277106893 letab = -7.15483625102932e-09 wetab = -6.38347978996382e-08 petab = 3.24340548434633e-14
+ dsub = 0.229245027302589 ldsub = 4.46472578592628e-08 wdsub = -3.43861778215202e-07 pdsub = 1.07590547660126e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.261300708411208 lpclm = 1.81297455592968e-07 wpclm = 1.47685171026069e-06 ppclm = -7.37223014476352e-13
+ pdiblc1 = -0.390722190826025 lpdiblc1 = 2.40911022182277e-07 wpdiblc1 = 2.83985219114751e-07 ppdiblc1 = -3.15438430929611e-13
+ pdiblc2 = -0.0182732804499644 lpdiblc2 = 9.42145957090192e-09 wpdiblc2 = 6.25571715161098e-08 ppdiblc2 = -3.15121116793246e-14
+ pdiblcb = -0.24960113465974 lpdiblcb = 1.23924033655549e-08 wpdiblcb = -8.97354982773187e-07 ppdiblcb = 4.52027317537286e-13
+ drout = 2.25214637525071 ldrout = -6.30747450044167e-07 wdrout = -5.01287350110126e-06 pdrout = 2.52514980733024e-12
+ pscbe1 = 800012629.676785 lpscbe1 = -0.00636198497659279 wpscbe1 = -0.0635327327836421 ppscbe1 = 3.20035340815178e-8
+ pscbe2 = 6.30654195003831e-08 lpscbe2 = -1.68399249806988e-14 wpscbe2 = -3.77188570622473e-13 ppscbe2 = 1.1744098683543e-19
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -7.10671732919327e-09 lalpha0 = 3.63026134038652e-15 walpha0 = -6.68903838664835e-15 palpha0 = 3.36948937362154e-21
+ alpha1 = 2.014932e-10 lalpha1 = -5.11254741156e-17
+ beta0 = 3.13293609550798 lbeta0 = 3.14691947908859e-06 wbeta0 = -6.29619074417743e-08 pbeta0 = 1.17080499569982e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = -50543825.4421301 lbgidl = 279.98520685186 wbgidl = 3603.00631556265 pbgidl = -5.40534266311142e-6
+ cgidl = 468.721735145804 lcgidl = -8.49907058102016e-05 wcgidl = 0.000483598132329611 pcgidl = -2.43604337992792e-10
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.480497067011927 lkt1 = -1.40858521228809e-08 wkt1 = 1.63318606864722e-07 pkt1 = -8.22689717917865e-14
+ kt2 = 0.021924189806907 lkt2 = -3.88439547080027e-08 wkt2 = -6.56863847389971e-08 pkt2 = 3.30883996437294e-14
+ at = 14776.0530722971 lat = 0.0355568185467419 wat = 0.337775448328289 pat = -2.06847700505062e-7
+ ute = -0.483461141257362 lute = -9.64121282752766e-09 wute = 7.44191525945833e-07 pute = 9.38408711207407e-14
+ ua1 = 9.16709709775115e-10 lua1 = -2.19923555707135e-16 wua1 = -9.60400933551529e-16 pua1 = 3.94710253673558e-22
+ ub1 = 3.00392331791239e-19 lub1 = 1.33954844151359e-26 wub1 = 9.362460951418e-25 pub1 = -1.67069296561781e-31
+ uc1 = -4.79871323193846e-11 luc1 = 3.64234886846406e-17 wuc1 = 4.10845005312876e-16 puc1 = -2.06956187061271e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.16 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.752085361422663+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -6.16418970300059e-08 wvth0 = -5.0380414670359e-07 pvth0 = 1.13492004930827e-13
+ k1 = 0.402548019445497 lk1 = 1.07905800435862e-07 wk1 = -6.7946695194518e-07 pk1 = 1.66625388590326e-13
+ k2 = 0.0463787216430325 lk2 = -3.92591588811166e-08 wk2 = 2.26251882224597e-07 pk2 = -4.9480182364328e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 377699.797421018 lvsat = -0.0552316314055003 wvsat = -1.3485998663872 pvsat = 2.57523334048288e-7
+ ua = -1.81334425565846e-09 lua = -8.42141390209225e-17 wua = 1.76994848884881e-15 pua = -3.31272528037942e-22
+ ub = 1.38372678100913e-18 lub = 9.98970688493881e-26 wub = -2.41135689048691e-25 pub = 1.0478431701489e-31
+ uc = 1.60296732358923e-13 luc = -3.06824061599317e-20 wuc = -1.53403619582221e-18 puc = 4.90824975229764e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00413046609004372 lu0 = -7.76791103660845e-11 wu0 = 1.08722804803487e-08 pu0 = -2.28126349228498e-15
+ a0 = 0.778431492647826 la0 = -3.97352304763016e-08 wa0 = 1.42115998717191e-06 pa0 = -3.00686332607182e-13
+ keta = -0.231769866615295 lketa = 5.0202190863154e-08 wketa = -2.74203322980789e-08 pketa = -7.87195832349672e-14
+ a1 = 0.0
+ a2 = 0.805420971608987 la2 = -1.37547938926351e-09 wa2 = 4.84043202004885e-07 pa2 = -1.22817733774306e-13
+ ags = 2.18807577984666 lags = -1.72355477258567e-07 wags = 1.37529009240526e-05 pags = -2.52686174547895e-12
+ b0 = 0.0
+ b1 = 1.39123192780888e-23 lb1 = -3.53001450738731e-30 wb1 = -9.78096174293563e-29 pb1 = 2.48175276592029e-35
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.244640914059811+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -6.26850506580921e-09 wvoff = 1.04216848848363e-06 pvoff = -3.51703090963557e-13
+ nfactor = {2.02412486521204+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -9.35359033048966e-08 wnfactor = -8.9170542464456e-06 pnfactor = 2.97738390439051e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -4.08983213941502 leta0 = 7.70404295878499e-07 weta0 = 2.56438298811856e-05 peta0 = -4.62431012422977e-12
+ etab = 0.108548866178091 letab = -3.11291383693785e-08 wetab = 1.64543406723525e-07 petab = -2.55130321501858e-14
+ dsub = 0.85854118398817 ldsub = -1.1502594386504e-07 wdsub = -6.41832028953577e-07 pdsub = 1.83195433290727e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.87560948692154 lpclm = -2.28305953704795e-07 wpclm = -5.24054148209731e-06 ppclm = 9.67201312400219e-13
+ pdiblc1 = 1.56293106007215 lpdiblc1 = -2.5479527812787e-07 wpdiblc1 = -3.66960121677749e-06 ppdiblc1 = 6.87716916208636e-13
+ pdiblc2 = 0.0576976767070423 lpdiblc2 = -9.85487930141688e-09 wpdiblc2 = -2.25503114455354e-07 ppdiblc2 = 4.15782888610729e-14
+ pdiblcb = -0.530852376215214 lpdiblcb = 8.37551246391499e-08 wpdiblcb = 3.20483922418995e-06 ppdiblcb = -5.88834725178093e-13
+ drout = -3.59337263456052 ldrout = 8.52453624872266e-07 wdrout = 1.96843629658594e-05 pdrout = -3.74135409314109e-12
+ pscbe1 = 799954894.011478 lpscbe1 = 0.00828745858916591 wpscbe1 = 0.226902617076121 ppscbe1 = -4.16894985425659e-8
+ pscbe2 = -3.50445059549781e-08 lpscbe2 = 8.05380073486643e-15 wpscbe2 = 3.02927419244911e-13 ppscbe2 = -5.51268836215906e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.58382761756902e-08 lalpha0 = -4.72897069658809e-15 walpha0 = 2.38894228094585e-14 palpha0 = -4.38927532105022e-21
+ alpha1 = -2.62475714285714e-10 lalpha1 = 6.65987504128571e-17
+ beta0 = 33.5796656460607 lbeta0 = -4.57842054996179e-06 wbeta0 = 2.46881467504535e-06 pbeta0 = -5.25314768034245e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.99974125349601e-11 lagidl = 3.0447303474733e-17 wagidl = 6.03638847932548e-16 pagidl = -1.53163095802469e-22
+ bgidl = 1806746721.25756 lbgidl = -191.270695433894 wbgidl = 8659.62018859581 pbgidl = -0.00128843515050944
+ cgidl = -302.57762552073 lcgidl = 0.0001107133948698 wcgidl = -0.00172713618689147 pcgidl = 3.1733191302613e-10
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.536011533489999 wkt1 = -1.60915811960526e-7
+ kt2 = -0.131165690926 wkt2 = 6.47199859093978e-8
+ at = 562385.294062613 lat = -0.103389716997454 wat = -2.43795839920244 pat = 4.97447575830453e-7
+ ute = -1.10273369403117 lute = 1.47488669805429e-07 wute = 4.03809742247934e-06 pute = -7.41931753724397e-13
+ ua1 = -1.72259819668082e-10 lua1 = 5.63839499070758e-17 wua1 = 2.15749776572468e-15 pua1 = -3.96403536989892e-22
+ ub1 = 2.4947118339318e-19 lub1 = 2.6315860161621e-26 wub1 = 1.00696048424049e-24 pub1 = -1.85011870650957e-31
+ uc1 = 9.55633269611999e-11 wuc1 = -4.04800523890149e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.17 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.850923742713245+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -4.34820247203432e-08 wvth0 = 5.78845429245078e-07 pvth0 = -8.54264496069482e-14
+ k1 = -0.492330911058914 lk1 = 2.72324590974229e-07 wk1 = 1.0587659410571e-06 pk1 = -1.52745355539662e-13
+ k2 = 0.469618568939547 lk2 = -1.17022285744447e-07 wk2 = -5.49285381715923e-07 pk2 = 9.30116057512559e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 253560.091371957 lvsat = -0.0324230707939882 wvsat = -0.123964072931356 pvsat = 3.25173258092643e-8
+ ua = -1.69882046907165e-09 lua = -1.05255937901879e-16 wua = 5.0670854054829e-15 pua = -9.37065385141873e-22
+ ub = 1.38744704983717e-18 lub = 9.9213532696808e-26 wub = -5.14265373780624e-24 pub = 1.00535493266727e-30
+ uc = -6.06006134606363e-13 luc = 1.10112718496201e-19 wuc = 6.21605057064256e-18 puc = -9.33121716633109e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00491718546219112 lu0 = -2.2222542076884e-10 wu0 = 9.47939470488931e-09 pu0 = -2.02534441010249e-15
+ a0 = 1.20712043139365 la0 = -1.18499535258888e-07 wa0 = -1.47231579113891e-05 pa0 = 2.66555762784912e-12
+ keta = 0.291081587447803 lketa = -4.58628753462212e-08 wketa = -2.7249356443574e-06 pketa = 4.16902997595628e-13
+ a1 = 0.0
+ a2 = -2.40541921479392 la2 = 5.88561820579103e-07 wa2 = 1.41297381208853e-05 pa2 = -2.62998219830495e-12
+ ags = 1.25
+ b0 = 0.0
+ b1 = -3.24620783155406e-23 lb1 = 4.990492685683e-30 wb1 = 2.28222440668498e-28 pb1 = -3.50853204712902e-35
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.195650633742748+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -8.71645920182166e-08 wvoff = -3.24323655786297e-06 pvoff = 4.35667234416845e-13
+ nfactor = {-4.02206929016926+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 1.01734948744577e-06 wnfactor = 2.33123651026435e-05 pnfactor = -2.94422400087568e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -1.63337483502509 leta0 = 3.19072025971024e-07 weta0 = 6.74204147416827e-06 peta0 = -1.15142783484325e-12
+ etab = -0.243544075417125 letab = 3.35619540687353e-08 wetab = -1.20735257293199e-07 petab = 2.69020726255993e-14
+ dsub = 0.09152744975529 ldsub = 2.589979056677e-08 wdsub = 2.17565697049997e-06 pdsub = -3.34470273045871e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.93582810211273 lpclm = -6.06836100529717e-07 wpclm = -1.20242464252813e-05 ppclm = 2.21359177272623e-12
+ pdiblc1 = 0.978965416199412 lpdiblc1 = -1.475015184822e-07 wpdiblc1 = 4.49664120405898e-07 ppdiblc1 = -6.91280619880792e-14
+ pdiblc2 = 0.0361061133190584 lpdiblc2 = -5.88779658545242e-09 wpdiblc2 = -8.96249915396316e-08 ppdiblc2 = 1.66129937033985e-14
+ pdiblcb = -1.3704596315583 lpdiblcb = 2.38018684485101e-07 wpdiblcb = 6.51672184439101e-06 ppdiblcb = -1.19733685463549e-12
+ drout = 1.28331635355196 ldrout = -4.35550729806028e-08 wdrout = -4.15623441116152e-06 pdrout = 6.38950384731095e-13
+ pscbe1 = 1053745053.24314 lpscbe1 = -46.6213398675209 wpscbe1 = -1276.44728642498 ppscbe1 = 0.000234525489276721
+ pscbe2 = 1.16529804552043e-08 lpscbe2 = -5.26068535735616e-16 wpscbe2 = -1.0209878978835e-14 ppscbe2 = 2.40677159295291e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 19.380148875601 lbeta0 = -1.96950073517493e-06 wbeta0 = -3.15054521140616e-05 pbeta0 = 5.7168791919288e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 8.85369385140146e-10 lagidl = -1.35898454362507e-16 wagidl = -4.96149828902033e-15 pagidl = 8.69336245781294e-22
+ bgidl = -1260646407.09446 lbgidl = 372.310646217609 wbgidl = 14241.6751522008 pbgidl = -0.00231404285513747
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = 0.214424925572597 lkt1 = -1.37879941932948e-07 wkt1 = -7.13671233838841e-07 pkt1 = 1.01559411927967e-13
+ kt2 = -0.178339640363558 lkt2 = 8.66741125201095e-09 wkt2 = 3.96373239036382e-07 pkt2 = -6.09356471567802e-14
+ at = -196761.125448261 lat = 0.0360905320985374 wat = 1.65047217565969 pat = -2.53732038980691e-7
+ ute = -0.3
+ ua1 = 1.3462e-10
+ ub1 = 3.927e-19
+ uc1 = 3.90619624918739e-10 luc1 = -5.42115787926325e-17 wuc1 = -2.47917382186362e-15 puc1 = 3.81130829156561e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.18 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0551071475136+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = 5.31724104111628e-8
+ k1 = 0.44197932961901 wk1 = -5.74263556878937e-8
+ k2 = 0.0242577805060215 wk2 = -4.64812692873905e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 322250.46307945 wvsat = -0.814617943877277
+ ua = -1.08156655008669e-09 wua = 2.64261803363704e-15
+ ub = 1.12029676449825e-18 wub = -9.45213454097547e-25
+ uc = -9.6192749169918e-12 wuc = -2.69674382780597e-16
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00821518957419 wu0 = 1.16017382291903e-8
+ a0 = 1.3187341681914 wa0 = -7.78027611856234e-7
+ keta = -0.0122354112795964 wketa = 3.70936478479419e-8
+ a1 = 0.0
+ a2 = 1.07610503033547 wa2 = -8.36717574510579e-7
+ ags = 0.371042957725606 wags = -5.83421315510329e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.259638531068819+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = -8.29158037068265e-8
+ nfactor = {1.44930088139524+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor = 8.55145900212889e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.346247533159597 wpclm = -5.9843939635282e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000133562314706127 wpdiblc2 = 1.76758095666019e-10
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 864959920.378692 wpscbe1 = -326.776475182409
+ pscbe2 = 7.8706837911503e-09 wpscbe2 = 6.06861384804025e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.24526776033921e-10 walpha0 = -6.26423503923224e-16
+ alpha1 = 2.51521514455741e-10 walpha1 = -7.62218705310926e-16
+ beta0 = 1.30770589641956 wbeta0 = 2.53707735405587e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1830081692.44049 wbgidl = -1447.15620639806
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.423527863674774 wkt1 = -6.3010068556414e-8
+ kt2 = -0.0473098436534728 wkt2 = -1.622728060345e-8
+ at = 90000.0
+ ute = -0.154818536779372 wute = -4.97689493021047e-8
+ ua1 = 1.73130733108857e-09 wua1 = 1.14718789464818e-15
+ ub1 = -7.7356927328652e-19 wub1 = 1.06353967452558e-25
+ uc1 = 1.1395029153969e-10 wuc1 = -1.0159619529392e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.19 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0551071475136+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = 5.31724104111628e-8
+ k1 = 0.44197932961901 wk1 = -5.74263556878946e-8
+ k2 = 0.0242577805060215 wk2 = -4.64812692873903e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 322250.46307945 wvsat = -0.814617943877276
+ ua = -1.08156655008669e-09 wua = 2.64261803363704e-15
+ ub = 1.12029676449825e-18 wub = -9.45213454097547e-25
+ uc = -9.61927491699185e-12 wuc = -2.69674382780597e-16
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00821518957419 wu0 = 1.16017382291903e-8
+ a0 = 1.3187341681914 wa0 = -7.78027611856234e-7
+ keta = -0.0122354112795964 wketa = 3.70936478479419e-8
+ a1 = 0.0
+ a2 = 1.07610503033547 wa2 = -8.36717574510581e-7
+ ags = 0.371042957725606 wags = -5.83421315510329e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.259638531068819+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = -8.29158037068265e-8
+ nfactor = {1.44930088139524+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor = 8.55145900212885e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.346247533159597 wpclm = -5.9843939635282e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000133562314706127 wpdiblc2 = 1.76758095666019e-10
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 864959920.378692 wpscbe1 = -326.776475182409
+ pscbe2 = 7.87068379115031e-09 wpscbe2 = 6.06861384804028e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.24526776033921e-10 walpha0 = -6.26423503923224e-16
+ alpha1 = 2.51521514455741e-10 walpha1 = -7.62218705310926e-16
+ beta0 = 1.30770589641956 wbeta0 = 2.53707735405587e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1830081692.44049 wbgidl = -1447.15620639805
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.423527863674774 wkt1 = -6.30100685564148e-8
+ kt2 = -0.0473098436534728 wkt2 = -1.622728060345e-8
+ at = 90000.0
+ ute = -0.154818536779372 wute = -4.97689493021047e-8
+ ua1 = 1.73130733108857e-09 wua1 = 1.14718789464817e-15
+ ub1 = -7.7356927328652e-19 wub1 = 1.06353967452558e-25
+ uc1 = 1.1395029153969e-10 wuc1 = -1.01596195293922e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.20 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.06176714994021+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.330488120191e-08 wvth0 = 5.73303817832914e-08 pvth0 = -3.3279292684119e-14
+ k1 = 0.530487020412317 lk1 = -7.08391925556188e-07 wk1 = -4.23961526530476e-07 pk1 = 2.93364964253341e-12
+ k2 = -0.00675130069498674 lk2 = 2.48188406508189e-07 wk2 = 1.26644885004757e-07 pk2 = -1.05083421228151e-12
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 547124.508078514 lvsat = -1.7998318148025 wvsat = -1.42445042383115 pvsat = 4.88093634427864e-6
+ ua = -1.59424064035679e-09 lua = 4.10330653453978e-15 wua = 4.43053832322399e-15 pua = -1.43100366231366e-20
+ ub = 1.35855186448395e-18 lub = -1.90693020617386e-24 wub = -1.66131889111918e-24 pub = 5.7315167177695e-30
+ uc = 5.54441825142105e-12 luc = -1.21366151413901e-16 wuc = -3.56187080621841e-16 puc = 6.92424534630989e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00576142778001046 lu0 = 1.9639254246214e-08 wu0 = 2.03380556938115e-08 pu0 = -6.99231523900644e-14
+ a0 = 1.37609085268896 la0 = -4.59067588483716e-07 wa0 = -9.84957258693119e-07 pa0 = 1.65620964306674e-12
+ keta = -0.0128892221103971 lketa = 5.2329273222373e-09 wketa = 6.84815462387128e-08 pketa = -2.5122035815086e-13
+ a1 = 0.0
+ a2 = 1.3524677356905 la2 = -2.21193330481932e-06 wa2 = -1.67421601569757e-06 pa2 = 6.70311391117688e-12
+ ags = 0.441157948017916 lags = -5.61181661597241e-07 wags = -1.36594717903995e-06 pags = 6.26312807728552e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.254915029127204+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -3.78056483656642e-08 wvoff = -1.21858219182343e-07 pvoff = 3.1168469584111e-13
+ nfactor = {1.52070887623684+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.71530524777563e-07 wnfactor = 6.20283840921654e-07 pnfactor = 1.87977321439719e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.210473138764475 lpclm = 1.08670200097526e-06 wpclm = -9.87598051284599e-07 ppclm = 3.11472196871309e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000322686695925676 lpdiblc2 = -1.51370105107148e-09 wpdiblc2 = -4.66469165694935e-10 ppdiblc2 = 5.1482192582543e-15
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 929980464.603077 lpscbe1 = -520.407075486673 wpscbe1 = -653.857914510281 ppscbe1 = 0.00261787250963599
+ pscbe2 = 6.34412702422363e-09 lpscbe2 = 1.22181527718244e-14 wpscbe2 = 1.17928045361014e-14 ppscbe2 = -4.58148939083278e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.19589532094321e-10 lalpha0 = 3.95163822484289e-17 walpha0 = -6.01587033030204e-16 palpha0 = -1.98784481690005e-22
+ alpha1 = 2.5286424956465e-10 lalpha1 = -1.07468933014344e-17 walpha1 = -7.68973243238853e-16 palpha1 = 5.40615181134988e-23
+ beta0 = -9.62571745476535 lbeta0 = 8.75082012788493e-05 wbeta0 = 7.8765053928818e-05 pbeta0 = -4.27353563954763e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.54202375684171e-10 lagidl = -4.33821342941799e-16 wagidl = -2.72661375958152e-16 pagidl = 2.18230885258167e-21
+ bgidl = 1435806602.16471 lbgidl = 3155.67255111826 wbgidl = 817.014843550642 pbgidl = -0.0181218205501191
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.368985021702377 lkt1 = -4.3654634420826e-07 wkt1 = -2.02371993958821e-07 pkt1 = 1.11541564128678e-12
+ kt2 = -0.043188243409902 lkt2 = -3.2988187882276e-08 wkt2 = -3.24697053165232e-08 pkt2 = 1.3000003067604e-13
+ at = 12875.9883250619 lat = 0.617279997335087 wat = 0.366206652957658 pat = -2.93102027309675e-6
+ ute = -0.0281670312461897 lute = -1.01368483433561e-06 wute = -4.81049608973706e-07 pute = 3.45185524807536e-12
+ ua1 = 1.28085206676243e-09 lua1 = 3.60532366411086e-15 wua1 = 2.29544640239903e-15 pua1 = -9.19035451101631e-21
+ ub1 = -6.23808352507214e-19 lub1 = -1.19864642375171e-24 wub1 = 2.1280718974524e-25 pub1 = -8.5202316822028e-31
+ uc1 = 3.58470258571152e-10 luc1 = -1.95707252928862e-15 wuc1 = -2.03287205237099e-17 puc1 = 8.13907692085563e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.21 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.05850891776324+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.02597895133367e-08 wvth0 = 5.57052985937478e-08 pvth0 = -2.67728934904185e-14
+ k1 = 0.373212429032384 lk1 = -7.87064539868342e-08 wk1 = 7.38324917106177e-08 pk1 = 9.40615304498942e-13
+ k2 = 0.0456371716177361 lk2 = 3.84389510901547e-08 wk2 = -4.20428893015999e-08 pk2 = -3.75453403594602e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 98061.5722514518 lvsat = -0.00190371955480373 wvsat = -0.190982319486844 pvsat = -5.75406095320924e-8
+ ua = 1.1965190759705e-10 lua = -2.75866161815711e-15 wua = 3.43268601005354e-16 pua = 2.05430004361093e-21
+ ub = 4.60455906063701e-19 lub = 1.68880621971992e-24 wub = 2.54771866038559e-25 pub = -1.93999907765794e-30
+ uc = -6.07921508805809e-11 luc = 1.44227759526677e-16 wuc = -1.37006910002429e-16 puc = -1.8511434742358e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0135427828588655 lu0 = -1.15152138677157e-08 wu0 = 1.38751925576714e-09 pu0 = 5.94973571463616e-15
+ a0 = 1.0012757541528 la0 = 1.04159199042377e-06 wa0 = 7.77987914604482e-07 pa0 = -5.40215212445558e-12
+ keta = -0.0140622345732879 lketa = 9.92935602932465e-09 wketa = 4.99778146083035e-08 pketa = -1.77136357199046e-13
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.367681303341791 lags = -2.67000794578166e-07 wags = -8.17080357391235e-07 pags = 4.06561187084545e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.261120292038855+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.29614324726126e-08 wvoff = -5.84712415954529e-08 pvoff = 5.79001619062136e-14
+ nfactor = {1.65163121968883+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.09570863169361e-06 wnfactor = 6.00698507978873e-07 pnfactor = 1.95818765821619e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.280332899879597 leta0 = -8.02079442233639e-07 weta0 = -6.07095270514508e-07 peta0 = 2.43064736870286e-12
+ etab = -0.245133796125758 letab = 7.01188958963969e-07 wetab = 5.30731095087732e-07 petab = -2.12490559952889e-12
+ dsub = 1.3159732252552 ldsub = -3.02671494907066e-06 wdsub = -2.2909256041512e-06 pdsub = 9.17225444188509e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.0145528229692635 lpclm = 1.98764586982536e-06 wpclm = 1.28550228297201e-06 ppclm = -5.98616485186115e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -0.000868056947899335 lpdiblc2 = 3.25371857025096e-09 wpdiblc2 = 3.28213064934787e-09 ppdiblc2 = -9.86017352502647e-15
+ pdiblcb = 0.0109204723674743 lpdiblcb = -1.43815980593245e-07 wpdiblcb = -1.80695500836553e-07 ppdiblcb = 7.23456539650834e-13
+ drout = 0.56
+ pscbe1 = 829102575.257112 lpscbe1 = -116.518940941881 wpscbe1 = -88.1933811620747 ppscbe1 = 0.000353102750540176
+ pscbe2 = 8.69645746427683e-09 lpscbe2 = 2.80004976207878e-15 wpscbe2 = 3.92026939850948e-15 ppscbe2 = -1.42953651842915e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.83915422542303e-10 lalpha0 = -2.18027308092544e-16 walpha0 = -9.25174063633408e-16 palpha0 = 1.09677159110805e-21
+ alpha1 = 4.00640373600396e-10 lalpha1 = -6.02403037715442e-16 walpha1 = -1.51235101597946e-15 palpha1 = 3.03034763830158e-21
+ beta0 = 13.6318519792571 lbeta0 = -5.6088969639376e-06 wbeta0 = -4.28963321509202e-05 pbeta0 = 5.97461423184248e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 8.10275466949416e-11 lagidl = -1.40848865348264e-16 wagidl = 9.54396400187618e-17 pagidl = 7.08530667581372e-22
+ bgidl = 2580326219.96692 lbgidl = -1426.67841182384 wbgidl = -4789.07146349204 pbgidl = 0.00432345219823584
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.504948820482291 lkt1 = 1.0781640377224e-07 wkt1 = 2.23900633987395e-07 pkt1 = -5.91266146218203e-13
+ kt2 = -0.0753745832487117 lkt2 = 9.58773230795813e-08 wkt2 = 8.70621679172569e-08 pkt2 = -3.48573674741863e-13
+ at = 175303.16561431 lat = -0.0330350524747263 wat = -0.33289316940324 pat = -1.32011244016291e-7
+ ute = -1.41002231293085 lute = 4.51889475816957e-06 wute = 6.50816835747906e-06 pute = -2.45311073684045e-11
+ ua1 = 3.21248919943146e-10 lua1 = 7.44731844993507e-15 wua1 = 1.27935938539862e-14 pua1 = -5.12221339018018e-20
+ ub1 = 4.67871847788181e-19 lub1 = -5.56944246712099e-24 wub1 = -8.8846617979768e-24 pub1 = 3.5571813634399e-29
+ uc1 = -5.33045177925385e-10 luc1 = 1.61231724382197e-15 wuc1 = 7.93963108427395e-16 puc1 = -3.17881629799334e-21
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.22 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0340896596396+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -8.669883824527e-09 wvth0 = -4.21283629971866e-08 pvth0 = 1.69259642750171e-13
+ k1 = 0.0996745177206462 lk1 = 4.69390485659568e-07 wk1 = 1.35178669146604e-06 pk1 = -1.62006369803959e-12
+ k2 = 0.160729449161298 lk2 = -1.92175243469039e-07 wk2 = -5.60093186701856e-07 pk2 = 6.62581072966105e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 251856.57490261 lvsat = -0.310067841602018 wvsat = -0.869511687881406 pvsat = 1.30205107738925e-6
+ ua = -1.66804499263397e-09 lua = 8.23405654833496e-16 wua = 4.30211435754029e-15 pua = -5.87816984066808e-21
+ ub = 1.55924906713604e-18 lub = -5.12881897295037e-25 wub = -2.51898886989039e-24 pub = 3.61787684302719e-30
+ uc = 5.29525612667361e-11 luc = -8.3686273778403e-17 wuc = -4.60629378232021e-16 puc = 4.63338671709504e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00606337850448048 lu0 = 3.47151545750934e-09 wu0 = 1.67661918704429e-08 pu0 = -2.48650180995859e-14
+ a0 = 3.18675321918251 la0 = -3.33752132701261e-06 wa0 = -7.32791157297951e-06 pa0 = 1.08399061734995e-11
+ keta = 0.10150378234503 lketa = -2.21634085748467e-07 wketa = -4.15827770394485e-07 pketa = 7.56213665055345e-13
+ a1 = 0.0
+ a2 = 0.8
+ ags = -1.79059333263795 lags = 4.05760531659743e-06 wags = 7.20278869206839e-06 pags = -1.20040643992354e-11
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.281502279525606+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.78786284601767e-08 wvoff = 3.86193924179184e-08 pvoff = -1.36643545457302e-13
+ nfactor = {0.519267133514538+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.17324665578866e-06 wnfactor = 3.87793821155857e-06 pnfactor = -4.60852568475668e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.732196329759194 leta0 = 1.22675878865819e-06 weta0 = 1.21419054102901e-06 peta0 = -1.21872311431868e-12
+ etab = -34.4225440615545 letab = 6.91835937623422e-05 wetab = 0.000173161546076199 petab = -3.48030966394076e-10
+ dsub = -0.650826550510391 ldsub = 9.14226666023446e-07 wdsub = 4.58185120830239e-06 pdsub = -4.59895525886299e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.8499049361474 lpclm = -1.74822966922274e-06 wpclm = -4.98850452725569e-06 ppclm = 6.58526963601685e-12
+ pdiblc1 = 0.39092545198256 lpdiblc1 = -1.85435867737242e-09 wpdiblc1 = 3.94722048558198e-08 ppdiblc1 = -7.90917594523653e-14
+ pdiblc2 = 0.00108275902786578 lpdiblc2 = -6.55195777316803e-10 wpdiblc2 = -3.28366003261672e-09 ppdiblc2 = 3.29591793551847e-15
+ pdiblcb = -0.121190811114683 lpdiblcb = 1.20899757792309e-07 wpdiblcb = 3.61501730154008e-07 ppdiblcb = -3.62961944593576e-13
+ drout = 0.227351650137107 ldrout = 6.66538476015825e-07 wdrout = 4.0151138438923e-07 pdrout = -8.04521610776385e-13
+ pscbe1 = 741794849.485777 lpscbe1 = 58.4224303410929 wpscbe1 = 176.386762324149 ppscbe1 = -0.000177045214107904
+ pscbe2 = 1.32282972846764e-08 lpscbe2 = -6.28054723676987e-15 wpscbe2 = -7.64576161313776e-15 ppscbe2 = 8.87987283276946e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.50490093264413e-10 lalpha0 = -1.51051872782569e-16 walpha0 = -7.57030210938307e-16 palpha0 = 7.59856204715739e-22
+ alpha1 = 1.0e-10
+ beta0 = 12.6604182177895 lbeta0 = -3.66240307877091e-06 wbeta0 = -2.57973788849036e-05 pbeta0 = 2.54844053938496e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -7.88645961265686e-11 lagidl = 1.79532297663909e-16 wagidl = 8.99766223795085e-16 pagidl = -9.03125051108512e-22
+ bgidl = 2578620710.96468 lbgidl = -1423.26102715426 wbgidl = -5387.45425069637 pbgidl = 0.00552245153558914
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.391040993952746 lkt1 = -1.20424467203285e-07 wkt1 = -3.29476105368793e-07 pkt1 = 5.17553087862189e-13
+ kt2 = -0.0110390401760913 lkt2 = -3.30339276479498e-08 wkt2 = -1.55128976554716e-07 pkt2 = 1.36712713744396e-13
+ at = 352601.957742806 lat = -0.388294493122733 wat = -1.10029900647906 pat = 1.40566515612516e-6
+ ute = 1.68054780296696 lute = -1.67378257186869e-06 wute = -1.02134288427488e-05 pute = 8.97450875439978e-12
+ ua1 = 3.66577333706654e-09 lua1 = 7.45784506039159e-16 wua1 = -1.29438281152103e-14 pua1 = 3.48787832802347e-22
+ ub1 = -7.28757950103794e-19 lub1 = -3.17171585230151e-24 wub1 = 4.38200299358217e-24 pub1 = 8.98895959161418e-30
+ uc1 = 7.16144639608873e-10 luc1 = -8.90725616835407e-16 wuc1 = -2.39620378559216e-15 puc1 = 3.21342638306114e-21
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.23 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.08623799204969+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.36731183104509e-08 wvth0 = 1.86423406646476e-07 pvth0 = -6.01453106495699e-14
+ k1 = 0.606815551743725 lk1 = -3.96437058435189e-08 wk1 = -2.90065344398547e-07 pk1 = 2.79173714748844e-14
+ k2 = -0.0550044072733476 lk2 = 2.43639474516768e-08 wk2 = 1.22436473946549e-07 pk2 = -2.24964709055003e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -137660.654577621 lvsat = 0.0809034556958634 wvsat = 0.570500992914045 pvsat = -1.43337170743611e-7
+ ua = -1.13305594033347e-10 lua = -7.37137585942105e-16 wua = -4.22279295178559e-15 pua = 2.67856094764351e-21
+ ub = 6.74206831586564e-19 lub = 3.75464200919743e-25 wub = 2.43849508167521e-24 pub = -1.35811339612961e-30
+ uc = -4.18463324797036e-11 luc = 1.14665042383922e-17 wuc = -3.44330991337664e-17 puc = 3.5551401901376e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0127554090486587 lu0 = -3.24549643669028e-09 wu0 = -1.92424081963505e-08 pu0 = 1.12780020712568e-14
+ a0 = -1.02990401711006 la0 = 8.94876690743043e-07 wa0 = 6.18002120323431e-06 pa0 = -2.71845171576789e-12
+ keta = -0.223041851712473 lketa = 1.04123077160973e-07 wketa = 6.65631198846509e-07 pketa = -3.29282390517825e-13
+ a1 = 0.0
+ a2 = 0.856465725237901 la2 = -5.66765117902138e-08 wa2 = -2.96877428494723e-07 pa2 = 2.97985671935294e-13
+ ags = 3.80494453248637 lags = -1.5588206913774e-06 wags = -1.0440782391772e-05 pags = 5.70537013546093e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.285334852206834+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 3.17255081352239e-08 wvoff = 7.18002668794606e-08 pvoff = -1.69948284123209e-13
+ nfactor = {1.57110751369142+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.17479755472577e-07 wnfactor = -1.11964683278924e-06 pnfactor = 4.07715344561683e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = 69.264468660018 letab = -3.48904825777199e-05 wetab = -0.00034844267878612 petab = 1.75520407039654e-10
+ dsub = 0.223730129051379 ldsub = 3.64052663768723e-08 wdsub = 2.03769503240768e-08 pdsub = -2.04530174796367e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.41290574631516 lpclm = 5.23028085517448e-07 wpclm = 3.16408854498889e-06 ppclm = -1.59775706616642e-12
+ pdiblc1 = 1.02035620663085 lpdiblc1 = -6.33634778332764e-07 wpdiblc1 = -1.38152934070124e-06 ppdiblc1 = 1.34721438487426e-12
+ pdiblc2 = 0.00067029686719512 lpdiblc2 = -2.4119389540036e-10 wpdiblc2 = -1.20879709829746e-09 ppdiblc2 = 1.2133095378654e-15
+ pdiblcb = 0.22519293275947 lpdiblcb = -2.26777036597726e-07 wpdiblcb = -2.21456961805826e-10 ppdiblcb = 1.11555179741311e-16
+ drout = 0.782011659725787 ldrout = 1.0980792061135e-07 wdrout = -8.03022768778461e-07 pdrout = 4.0450906838508e-13
+ pscbe1 = 800000000.0
+ pscbe2 = 2.56924744567959e-08 lpscbe2 = -1.87912531822729e-14 wpscbe2 = -6.1503912015007e-14 ppscbe2 = 6.29390757100889e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.5642599555547 lbeta0 = 4.4904614225683e-07 wbeta0 = -6.06325253554694e-07 pbeta0 = 1.99313559294857e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.64191885543993e-10 lagidl = -1.64804813852729e-16 wagidl = -8.25956148019218e-16 pagidl = 8.29039442319774e-22
+ bgidl = 766583401.446103 lbgidl = 395.54061764075 wbgidl = 1914.45560947643 pbgidl = -0.00180671635409168
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.513594272012911 lkt1 = 2.58630224388011e-09 wkt1 = 3.73694096384108e-07 pkt1 = -1.88242048253856e-13
+ kt2 = -0.0326283195140367 lkt2 = -1.13640555302358e-08 wkt2 = -3.79907185595965e-08 pkt2 = 1.91371786321812e-14
+ at = -135582.148513139 lat = 0.101712004401865 wat = 0.57948016947836 pat = -2.80384635496112e-7
+ ute = 0.346078857673474 lute = -3.34332054002432e-07 wute = -2.55409363643807e-06 pute = 1.28658124976386e-12
+ ua1 = 8.57200325689244e-09 lua1 = -4.17876037007745e-15 wua1 = -2.61409421742828e-14 pua1 = 1.35951667186573e-20
+ ub1 = -8.30240290353452e-18 lub1 = 4.43020151774037e-24 wub1 = 2.70035551502201e-23 pub1 = -1.37170388192245e-29
+ uc1 = -3.68316791693746e-10 luc1 = 1.97784108990266e-16 wuc1 = 1.61655513747474e-15 puc1 = -8.14312169065562e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.24 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.965433361769523+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.71801605144682e-08 wvth0 = -2.20298104716986e-09 pvth0 = 3.48720255025132e-14
+ k1 = 0.147745055347055 lk1 = 1.91605252517865e-07 wk1 = -6.64119954978304e-08 pk1 = -8.47442009269212e-14
+ k2 = 0.118642381937682 lk2 = -6.31076706179627e-08 wk2 = 1.40779404794095e-08 pk2 = 3.20872982335023e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 19343.0972682559 lvsat = 0.00181548476728438 wvsat = 0.23309561060012 pvsat = 2.66250547055294e-8
+ ua = -9.50702928494548e-10 lua = -3.1531291446196e-16 wua = 1.48846451633969e-15 pua = -1.98387910547637e-22
+ ub = 9.53544090140247e-19 lub = 2.3475280565672e-25 wub = -1.7623997094857e-25 pub = -4.0985063866274e-32
+ uc = -4.86489445123201e-11 luc = 1.48932044054183e-17 wuc = 1.23515443539894e-16 puc = -4.40124913452549e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00868111508935995 lu0 = -1.19314011769086e-09 wu0 = 5.21883956162168e-09 pu0 = -1.04393564560978e-15
+ a0 = 0.567434212241447 la0 = 9.02447124571195e-08 wa0 = 2.87704491301812e-06 pa0 = -1.05463356016841e-12
+ keta = 0.10646695516567 lketa = -6.18613826541747e-08 wketa = -1.61248828309685e-07 pketa = 8.72443662016456e-14
+ a1 = 0.0
+ a2 = 0.687068549524198 la2 = 2.86544357235767e-08 wa2 = 5.93754856989447e-07 pa2 = -1.50655201128504e-13
+ ags = -2.95447004901742 lags = 1.84611949400725e-06 wags = 1.22929002563963e-05 pags = -5.74633602594882e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.166891398871197+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -2.79383679438966e-08 wvoff = -2.25119595633298e-07 pvoff = -2.03799510200697e-14
+ nfactor = {1.57614431778768+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 1.14942551034755e-07 wnfactor = -1.57672141894755e-06 pnfactor = 6.37958897070968e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.362463978475422 leta0 = 6.42441027306404e-08 weta0 = 9.92738419557072e-07 peta0 = -5.00075102298742e-13
+ etab = 0.0047984347493751 letab = -2.10111613465856e-09 wetab = -1.72324063632499e-08 petab = 7.01165844028411e-15
+ dsub = 0.293145869470594 ldsub = 1.43826720828011e-09 wdsub = -6.6531063226425e-07 pdsub = 3.24950445560329e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.799815236488979 lpclm = -8.78594933134296e-08 wpclm = -1.23210911194954e-06 ppclm = 6.16752768156145e-13
+ pdiblc1 = -0.822741600675803 lpdiblc1 = 2.94794409435239e-07 wpdiblc1 = 2.45722956944807e-06 ppdiblc1 = -5.8649515721198e-13
+ pdiblc2 = -0.00452878511617366 lpdiblc2 = 2.37775526932795e-09 wpdiblc2 = -6.58358038374091e-09 ppdiblc2 = 3.92076524659169e-15
+ pdiblcb = -0.581394451588941 lpdiblcb = 1.79527646282252e-07 wpdiblcb = 7.71708802452271e-07 ppdiblcb = -3.88735190185689e-13
+ drout = 1.00618024871377 ldrout = -3.11319522533504e-09 wdrout = 1.25487462193944e-06 pdrout = -6.32121757933417e-13
+ pscbe1 = 800000000.0
+ pscbe2 = -4.42466276765124e-08 lpscbe2 = 1.64393805526449e-14 wpscbe2 = 1.62637406944101e-13 ppscbe2 = -4.99683033131396e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.13709706478601e-08 lalpha0 = 1.08156364573585e-14 walpha0 = 6.50663208165302e-14 palpha0 = -3.27760529838732e-20
+ alpha1 = 3.5527733068052e-10 lalpha1 = -1.28591615615691e-16 walpha1 = -7.73600642824297e-16 palpha1 = 3.89688172611812e-22
+ beta0 = -7.08646322853708 lbeta0 = 8.33283188394892e-06 wbeta0 = 5.13450335168927e-05 pbeta0 = -2.59703002482189e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.55915112773427e-09 lagidl = -1.82458451779896e-15 wagidl = -1.74010252176208e-14 pagidl = 9.17844870995736e-21
+ bgidl = 159158414.273688 lbgidl = 701.520628704073 wbgidl = 2548.11341648408 pbgidl = -0.00212591070218907
+ cgidl = 598.285985109728 lcgidl = -0.000150256494137278 wcgidl = -0.000168166042657757 pcgidl = 8.47107851661195e-11
+ egidl = 2.04672624427771 legidl = -9.80630251208742e-07 wegidl = -9.79287438379964e-06 pegidl = 4.93299399197454e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.396036534136916 lkt1 = -5.66314097296087e-08 wkt1 = -2.61554377338894e-07 pkt1 = 1.31753571160053e-13
+ kt2 = 0.0972092200947318 lkt2 = -7.67675088699795e-08 wkt2 = -4.44402625276846e-07 pkt2 = 2.23860267638581e-13
+ at = 66933.3315454859 lat = -0.00030172591450614 wat = 0.0754017952323933 pat = -2.64637238020681e-8
+ ute = -0.33552325116 lute = 9.01342108658029e-9
+ ua1 = 4.37917789120984e-10 lua1 = -8.13530951405335e-17 wua1 = 1.44812936120685e-15 pua1 = -3.02359053129504e-22
+ ub1 = 5.53360918686954e-19 lub1 = -3.07389597187192e-26 wub1 = -3.36295229966893e-25 pub1 = 5.49460323382655e-32
+ uc1 = 1.13975355330602e-11 luc1 = 6.50947179332496e-18 wuc1 = 1.12114459961633e-16 puc1 = -5.64757532598531e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.25 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.900937819654219+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -3.35448079020102e-08 wvth0 = 2.44988052233577e-07 pvth0 = -2.78484969449119e-14
+ k1 = 0.566402449992247 lk1 = 8.53780558023564e-08 wk1 = -1.50372555548022e-06 pk1 = 2.7994968058809e-13
+ k2 = -0.0160274574314221 lk2 = -2.89374882653218e-08 wk2 = 5.40181934919699e-07 pk2 = -1.01402646587816e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -138136.494517651 lvsat = 0.041773254029898 wvsat = 1.24627962650968 pvsat = -2.30453165203251e-7
+ ua = -1.81720911050816e-09 lua = -9.54517013811011e-17 wua = 1.78939037913309e-15 pua = -2.74742732491794e-22
+ ub = 1.68420104103326e-18 lub = 4.93610255357845e-26 wub = -1.75265108194523e-24 pub = 3.59002456560239e-31
+ uc = 3.59746036749668e-11 luc = -6.57858234678662e-18 wuc = -1.816954790606e-16 puc = 3.34295916789364e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00575367371017647 lu0 = -4.50351634226492e-10 wu0 = 2.70684460074756e-09 pu0 = -4.06559628202304e-16
+ a0 = 3.46045617752574 la0 = -6.43810429860361e-07 wa0 = -1.20705833488328e-05 pa0 = 2.73807300159581e-12
+ keta = -0.078258230061916 lketa = -1.49905072308237e-08 wketa = -7.99650211890896e-07 pketa = 2.49227864461857e-13
+ a1 = 0.0
+ a2 = 0.546101151806532 la2 = 6.44225164486733e-08 wa2 = 1.78853397363736e-06 pa2 = -4.53810090732927e-13
+ ags = 12.3829527865701 lags = -2.04549081433489e-06 wags = -3.75317366456088e-05 pags = 6.89581856910764e-12
+ b0 = 0.0
+ b1 = -1.39123192780888e-23 lb1 = 3.5300145073873e-30 wb1 = 4.2160340317001e-29 pb1 = -1.06974696296536e-35
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.142387050742026+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -1.06412516799609e-07 wvoff = -9.04749447955994e-07 pvoff = 1.52064570299325e-13
+ nfactor = {-1.00231239108507+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 7.69182107147165e-07 wnfactor = 6.30723317891103e-06 pnfactor = -1.36246055490748e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 1.65034549965664 leta0 = -2.62533939283234e-07 weta0 = -3.23174454812048e-06 peta0 = 5.71815634538986e-13
+ etab = 0.0439506870827838 letab = -1.20353345759714e-08 wetab = 4.89500166905924e-07 petab = -1.21563117573023e-13
+ dsub = 0.162639854992526 ldsub = 3.45519497798437e-08 wdsub = 2.8588524244489e-06 pdsub = -5.6924601930867e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.0569572764084025 lpclm = 1.29531966701562e-07 wpclm = 4.48110459280743e-06 ppclm = -8.32878084792955e-13
+ pdiblc1 = 0.688821684443156 lpdiblc1 = -8.87390775878504e-08 wpdiblc1 = 7.27546732708484e-07 ppdiblc1 = -1.47617541997536e-13
+ pdiblc2 = 0.00571633822123033 lpdiblc2 = -2.21770610441582e-10 wpdiblc2 = 3.59854844627738e-08 ppdiblc2 = -6.88041128410903e-15
+ pdiblcb = 0.951634991989341 lpdiblcb = -2.09452513525196e-07 wpdiblcb = -4.2527129689195e-06 ppdiblcb = 8.86126419129784e-13
+ drout = 1.56314854819377 ldrout = -1.44434432757294e-07 wdrout = -6.25516723184988e-06 pdrout = 1.27342369175411e-12
+ pscbe1 = 800000000.0
+ pscbe2 = 5.03350718637853e-08 lpscbe2 = -7.55911781681351e-15 wpscbe2 = -1.26568758237003e-13 ppscbe2 = 2.34128445967575e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.67820380280716e-08 lalpha0 = -1.40890208930117e-14 walpha0 = -2.32379717201893e-13 palpha0 = 4.26958225806554e-20
+ alpha1 = -8.11704752430428e-10 lalpha1 = 1.675102492783e-16 walpha1 = 2.7628594386582e-15 palpha1 = -5.07628453242986e-22
+ beta0 = 70.8148186515871 lbeta0 = -1.14332940713406e-05 wbeta0 = -0.000184840097975882 pbeta0 = 3.39576617208373e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.26252502173615e-08 lagidl = 2.28193218869622e-15 wagidl = 6.40135084464723e-14 pagidl = -1.1479105160234e-20
+ bgidl = 7358952436.22714 lbgidl = -1125.30470786824 wbgidl = -19270.3742210112 pbgidl = 0.00341015962153552
+ cgidl = -765.307089677598 lcgidl = 0.000195732067507734 wcgidl = 0.000600593009491985 pcgidl = -1.10348755412991e-10
+ egidl = -6.85259372956321 legidl = 1.27742090371384e-06 wegidl = 3.49745513707129e-05 pegidl = -6.42597924699519e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.873006566240141 lkt1 = 6.43916274260388e-08 wkt1 = 1.53431485202584e-06 pkt1 = -3.23917716014349e-13
+ kt2 = -0.448366205122709 lkt2 = 6.16629804967173e-08 wkt2 = 1.66037566638108e-06 pkt2 = -3.10191442638659e-13
+ at = 158526.980063159 lat = -0.0235420571338409 wat = -0.406376532221878 pat = 9.57793365578867e-8
+ ute = -0.3
+ ua1 = 7.18137540928753e-11 lua1 = 1.15395799792537e-17 wua1 = 9.29702201108482e-16 pua1 = -1.70816974516265e-22
+ ub1 = 5.3592881660682e-19 lub1 = -2.6315860161621e-26 wub1 = -4.34045217813203e-25 pub1 = 7.97484300044735e-32
+ uc1 = 3.7052345090055e-11 wuc1 = -1.10464996631925e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.26 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.775591869012523+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -5.65749954512611e-08 wvth0 = 1.99893546094628e-07 pvth0 = -1.9563148048484e-14
+ k1 = -0.113408247847117 lk1 = 2.10281714748476e-07 wk1 = -8.47378825273275e-07 pk1 = 1.5935712680698e-13
+ k2 = 0.297166161326424 lk2 = -8.64814914205572e-08 wk2 = 3.18224762508653e-07 pk2 = -6.06217894292168e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 166862.39521737 lvsat = -0.0142651069777868 wvsat = 0.312162809470494 pvsat = -5.88250800581903e-8
+ ua = -4.76562519885256e-10 lua = -3.4177272141602e-16 wua = -1.08140033881034e-15 pua = 2.52716258488103e-22
+ ub = -6.75575037889693e-20 lub = 3.71216878251606e-25 wub = 2.17664801990124e-24 pub = -3.62939455319319e-31
+ uc = 7.71753528304655e-13 luc = -1.10657080789949e-19 wuc = -7.14676001526163e-19 puc = 1.77445790483477e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00751190127067766 lu0 = -7.73396058600056e-10 wu0 = -3.57314724797038e-09 pu0 = 7.47282114138189e-16
+ a0 = -5.994167542703 la0 = 1.09331595012843e-06 wa0 = 2.15024329949795e-05 pa0 = -3.43039801030185e-12
+ keta = -0.741470907779387 lketa = 1.0686354768424e-07 wketa = 2.4692496758238e-06 pketa = -3.51376918607627e-13
+ a1 = 0.0
+ a2 = 2.54055202682437 la2 = -3.0202392617098e-07 wa2 = -1.07506348732254e-05 pa2 = 1.8500490190077e-12
+ ags = 1.25
+ b0 = 0.0
+ b1 = 3.24620783155406e-23 lb1 = -4.990492685683e-30 wb1 = -9.83741274063359e-29 pb1 = 1.51233497285582e-35
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.320877448527282+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -2.12955405553608e-08 wvoff = -6.4487706060756e-07 pvoff = 1.04317436954635e-13
+ nfactor = {4.87702645390899+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -3.1104645686013e-07 wnfactor = -2.14539326792507e-05 pnfactor = 3.73818173171015e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.141935608382891 leta0 = 1.4610735270166e-08 weta0 = -2.18853734534751e-06 peta0 = 3.80144045551901e-13
+ etab = -0.0536884802369407 letab = 5.90420255318363e-09 wetab = -1.07579095663776e-06 petab = 1.66032516429029e-13
+ dsub = 0.815455941906182 ldsub = -8.5391908317063e-08 wdsub = -1.46601622691332e-06 pdsub = 2.25375072612066e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.47553996410237 lpclm = -1.52038348789204e-07 wpclm = 3.52066245444073e-07 ppclm = -7.42374821168419e-14
+ pdiblc1 = 1.16074606021093 lpdiblc1 = -1.75447158920791e-07 wpdiblc1 = -4.64771084566387e-07 ppdiblc1 = 7.14505875238289e-14
+ pdiblc2 = 0.0119734504462039 lpdiblc2 = -1.37140861087264e-09 wpdiblc2 = 3.17727328477203e-08 ppdiblc2 = -6.10638979162041e-15
+ pdiblcb = -0.187223741544138 lpdiblcb = -2.06581836889634e-10 wpdiblcb = 5.64533923068111e-07 ppdiblcb = 1.03919592422475e-15
+ drout = -0.36551535173359 ldrout = 2.0992477156806e-07 wdrout = 4.1381016914878e-06 pdrout = -6.36162787337493e-13
+ pscbe1 = 800000000.0
+ pscbe2 = 1.04794862508309e-08 lpscbe2 = -2.36331505388553e-16 wpscbe2 = -4.3066959466416e-15 ppscbe2 = 9.4926910596262e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 10.6863326345987 lbeta0 = -3.85706949981313e-07 wbeta0 = 1.2228201045559e-05 pbeta0 = -2.2502880632691e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -9.43592389047907e-10 lagidl = 1.35626150926684e-16 wagidl = 4.23896991242438e-15 pagidl = -4.96549871757744e-22
+ bgidl = 2434823336.56926 lbgidl = -220.579696000802 wbgidl = -4348.13484045091 pbgidl = 0.000668451813427041
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = 0.33542011858788 lkt1 = -1.57636232657468e-07 wkt1 = -1.32232934882813e-06 pkt1 = 2.00942092941153e-13
+ kt2 = -0.0655803596364415 lkt2 = -8.66741125201095e-09 wkt2 = -1.70854677582147e-07 pkt2 = 2.62660021487363e-14
+ at = -8575.78352988337 lat = 0.00716023492939957 wat = 0.703818572105475 pat = -1.08200140545491e-7
+ ute = -0.3
+ ua1 = 1.3462e-10
+ ub1 = 3.927e-19
+ uc1 = 3.22730171810359e-11 luc1 = 8.78120254707823e-19 wuc1 = -6.76535507539113e-16 puc1 = 1.04005833180511e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.27 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 2e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.037561+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.42302944
+ k2 = 0.022723964
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 53438.0
+ ua = -2.0953977e-10
+ ub = 8.0838962e-19
+ uc = -9.8608028e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0120436
+ a0 = 1.061996
+ keta = 4.9707517e-6
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.17852213
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.28699958+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.731487+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.14877095
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00019189
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 757128280.0
+ pscbe2 = 9.873241e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.7815831e-11
+ alpha1 = 6.3056523e-17
+ beta0 = 9.6797043
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1352540500.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.4443203
+ kt2 = -0.052664618
+ at = 90000.0
+ ute = -0.17124159
+ ua1 = 2.1098632e-9
+ ub1 = -7.3847396e-19
+ uc1 = 1.1059776e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.28 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 2e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.037561+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.42302944
+ k2 = 0.022723964
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 53438.0
+ ua = -2.0953977e-10
+ ub = 8.0838962e-19
+ uc = -9.8608028e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0120436
+ a0 = 1.061996
+ keta = 4.9707517e-6
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.17852213
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.28699958+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.731487+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.14877095
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00019189
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 757128280.0
+ pscbe2 = 9.873241e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.7815831e-11
+ alpha1 = 6.3056523e-17
+ beta0 = 9.6797043
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1352540500.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.4443203
+ kt2 = -0.052664618
+ at = 90000.0
+ ute = -0.17124159
+ ua1 = 2.1098632e-9
+ ub1 = -7.3847396e-19
+ uc1 = 1.1059776e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.29 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 2e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.04284893035975+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.23231827220295e-8
+ k1 = 0.390585680091792 lk1 = 2.59671191821398e-7
+ k2 = 0.0350397299721097 lk2 = -9.85721025312519e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 77075.9045060112 lvsat = -0.189191476345611
+ ua = -1.32225313558197e-10 lua = -6.18804266400317e-16
+ ub = 8.10339998493619e-19 lub = -1.56103087118768e-26
+ uc = -1.11992308233283e-10 luc = 1.07124205384377e-16
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.012472700084275 lu0 = -3.43440250481465e-9
+ a0 = 1.05106881170975 la0 = 8.74582975158882e-8
+ keta = 0.00970872488828937 lketa = -7.76662572069069e-08 wketa = 1.80945758995975e-25 pketa = 4.42748183055293e-29
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.00958540767898763 lags = 1.50556250687006e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.295126527402052+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 6.50459171110712e-8
+ nfactor = {1.72539381884062+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.87681951202713e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.115420326624588 lpclm = 2.11451643903234e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0001687584325925 lpdiblc2 = 1.85138889401132e-10
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 714216549.967309 lpscbe1 = 343.454029749733
+ pscbe2 = 1.02355866437793e-08 lpscbe2 = -2.90011778652299e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.1074273105783e-11 lalpha0 = -2.60797006106449e-17
+ alpha1 = -8.86104341585482e-13 lalpha1 = 7.092647247765e-18 walpha1 = 2.69799463400731e-34 palpha1 = -1.0058856688555e-39
+ beta0 = 16.365642434038 lbeta0 = -5.35124636793581e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.42279568675574e-11 lagidl = 2.86309882096553e-16
+ bgidl = 1705410008.42162 lbgidl = -2824.27332924794
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.435764933148282 lkt1 = -6.84748719981981e-8
+ kt2 = -0.0539027894461152 lkt2 = 9.90999366293038e-9
+ at = 133719.032745477 lat = -0.349915465113059
+ ute = -0.18690663577313 lute = 1.25378843800912e-7
+ ua1 = 2.03831709184995e-09 lua1 = 5.72635946822119e-16
+ ub1 = -5.53584973233049e-19 lub1 = -1.4798020847232e-24
+ uc1 = 3.51762066741712e-10 luc1 = -1.93021472029077e-15 wuc1 = 1.97215226305253e-31
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.30 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 2e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.04012695277695+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.14251112484953e-8
+ k1 = 0.397576112770505 lk1 = 2.31683365821358e-7
+ k2 = 0.0317636095226659 lk2 = -8.54553909758389e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 35040.0931743605 lvsat = -0.020891311335307
+ ua = 2.32925717519395e-10 lua = -2.0807714995097e-15
+ ub = 5.44527038240345e-19 lub = 1.04863381208185e-24
+ uc = -1.06002504044869e-10 luc = 8.31426286916824e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.01400064469645 lu0 = -9.55188477075187e-9
+ a0 = 1.2580008228095 la0 = -7.41042224080547e-07 wa0 = -1.6940658945086e-21
+ keta = 0.0024297412604903 lketa = -4.8523150249828e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.0980562784389951 lags = 1.07459393598385e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.280414979310015+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 6.14480653389412e-9
+ nfactor = {1.8498532779084+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.49534248311533e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.409644848561555 lpclm = 1.22956699888001e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000215
+ pdiblcb = -0.0487065012492107 lpdiblcb = 9.49145013660063e-8
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 9.99009122335234e-09 lpscbe2 = -1.91721967041058e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.1379004976454e-11 lalpha0 = 1.43891889805384e-16 palpha0 = -9.4039548065783e-38
+ alpha1 = -9.84141889730421e-11 lalpha1 = 3.97569058113521e-16 walpha1 = -9.24446373305873e-33 palpha1 = 1.32243114467507e-37
+ beta0 = -0.523334251578298 lbeta0 = 1.41064896130743e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.12521285449025e-10 lagidl = 9.29562887750888e-17
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.431064760648385 lkt1 = -8.72931077417295e-8
+ kt2 = -0.0466452924507665 lkt2 = -1.91470865547483e-8
+ at = 65453.102180045 lat = -0.0765969061325282
+ ute = 0.737581701268525 lute = -3.57602561932789e-06 wute = -4.2351647362715e-22 pute = -8.07793566946316e-28
+ ua1 = 4.5429549373179e-09 lua1 = -9.45526524812681e-15 pua1 = -6.01853107621011e-36
+ ub1 = -2.46394157406524e-18 lub1 = 6.16875567979647e-24
+ uc1 = -2.71048520013885e-10 luc1 = 5.63352578651982e-16 puc1 = -3.76158192263132e-37
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.31 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 2e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.04799142685194+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.7183417480208e-8
+ k1 = 0.5457451116993 lk1 = -6.52077469092333e-8
+ k2 = -0.0240934241905149 lk2 = 2.64671907573741e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -35070.051563874 lvsat = 0.11959069931147 pvsat = 5.29395592033938e-23
+ ua = -2.4840776810201e-10 lua = -1.11630771036507e-15
+ ub = 7.28018172120339e-19 lub = 6.80966571919086e-25
+ uc = -9.9048654346014e-11 luc = 6.92089705730477e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0115959859888 lu0 = -4.73359076449619e-9
+ a0 = 0.76864547436 la0 = 2.39495236334213e-7
+ keta = -0.0357135328598723 lketa = 2.79057868331885e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.58622562145988 lags = 9.64329137845811e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.26875842324731+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.72118195152978e-8
+ nfactor = {1.7989321963259+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.47501996748984e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.33153053 leta0 = 8.2459730346849e-07 peta0 = 4.03896783473158e-28
+ etab = 22.718330456674 letab = -4.56617297509428e-05 wetab = 1.30231315640349e-20 petab = 1.41363874215605e-26
+ dsub = 0.8611199 ldsub = -6.033638805867e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.20376861036004 lpclm = 4.24816682389036e-7
+ pdiblc1 = 0.40395072436972 lpdiblc1 = -2.79535267935125e-8
+ pdiblc2 = -8.02595000000059e-07 lpdiblc2 = 4.32410781087135e-10
+ pdiblcb = -0.00190032504012002 lpdiblcb = 1.12742149203631e-9
+ drout = 0.359844759334281 ldrout = 4.01057660844845e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.07053034974741e-08 lpscbe2 = -3.35031410607337e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 6.80772026899032e-13 lalpha0 = 9.96899866511246e-17
+ alpha1 = 1.0e-10
+ beta0 = 4.1476460511977 lbeta0 = 4.74709223805208e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.1804560163172e-10 lagidl = -1.18486265862611e-16
+ bgidl = 800836588.0609 lbgidl = 399.070300894969
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.49976347432 lkt1 = 5.03607718996363e-8
+ kt2 = -0.062229420398 lkt2 = 1.20793448893457e-8
+ at = -10481.237611 lat = 0.0755552363400019
+ ute = -1.68974005325 lute = 1.28767908181878e-6
+ ua1 = -6.0550787332e-10 lua1 = 8.60879584821104e-16 wua1 = 3.94430452610506e-31
+ ub1 = 7.1724140061e-19 lub1 = -2.05485625598477e-25
+ uc1 = -7.4568904681e-11 luc1 = 1.69659889582174e-16 wuc1 = 2.46519032881566e-32 puc1 = -7.05296610493373e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.32 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 2e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.02472089008434+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.38260117988551e-8
+ k1 = 0.511098068145661 lk1 = -3.04313659420077e-8
+ k2 = -0.014602093060032 lk2 = 1.69404284877811e-08 wk2 = -3.30872245021211e-24
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 50596.6484282161 lvsat = 0.0336042055283096
+ ua = -1.5067678703996e-09 lua = 1.46749850194402e-16
+ ub = 1.4788759087153e-18 lub = -7.26941166065844e-26
+ uc = -5.32087708585482e-11 luc = 2.31979668005232e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0064056850072 lu0 = 4.7608561066812e-10
+ a0 = 1.0094160519 la0 = -2.17413777174299e-9
+ keta = -0.00339291884853741 lketa = -4.53548003025071e-9
+ a1 = 0.0
+ a2 = 0.758500349706741 la2 = 4.16545684878049e-8
+ ags = 0.359633203042341 lags = 3.23871201700074e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.26164177407776+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.43550351361978e-8
+ nfactor = {1.2016398078014+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.52020084261877e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = -45.7167141515031 letab = 2.30287828787567e-5
+ dsub = 0.23045423603654 ldsub = 2.96560583003356e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.631198967523641 lpclm = -4.20927229785539e-9
+ pdiblc1 = 0.5644709567641 lpdiblc1 = -1.8907298121542e-7
+ pdiblc2 = 0.00027141082767328 lpdiblc2 = 1.59181185707016e-10
+ pdiblcb = 0.225119855077083 lpdiblcb = -2.26740224957544e-07 wpdiblcb = -4.96308367531817e-23 ppdiblcb = -2.91878534931774e-29
+ drout = 0.51702544133144 ldrout = 2.4329022336179e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 5.397048604666e-09 lpscbe2 = 1.97775650224959e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.36418115044081 lbeta0 = 5.14816813283503e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -8.36202541933992e-12 lagidl = 1.0876654086023e-16
+ bgidl = 1398326823.8782 lbgidl = -200.650365972638
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.39028047658 lkt1 = -5.9530925870927e-8
+ kt2 = -0.0451647222620001 lkt2 = -5.04905576479597e-9
+ at = 55638.156458 lat = 0.00918901857294227
+ ute = -0.49673611652 lute = 9.02216613929694e-8
+ ua1 = -5.41399626399999e-11 lua1 = 3.07453417730535e-16 pua1 = 1.88079096131566e-37
+ ub1 = 6.0839046456e-19 lub1 = -9.62283490042026e-26
+ uc1 = 1.6512366524e-10 luc1 = -7.0927452702341e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.33 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 2e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.966160314528+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -5.67288260786694e-9
+ k1 = 0.125830030982599 lk1 = 1.63640858222252e-7
+ k2 = 0.123287904275852 lk2 = -5.25193135402158e-08 pk2 = 2.52435489670724e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 96261.3700479999 lvsat = 0.0106013783126108
+ ua = -4.595305748152e-10 lua = -3.80778134422215e-16
+ ub = 8.95387378715201e-19 lub = 2.21228311075956e-25
+ uc = -7.890585509966e-12 luc = 3.69701340325803e-19
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0104032587366 lu0 = -1.53762419676373e-9
+ a0 = 1.51681856508 la0 = -2.57769527943444e-7
+ keta = 0.0532571099463361 lketa = -3.30719689851787e-08 wketa = 2.64697796016969e-23
+ a1 = 0.0
+ a2 = 0.88299930058652 la2 = -2.10596615357195e-8
+ ags = 1.102014123899 lags = -5.0090566705815e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.24117769890236+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -3.46634651165276e-8
+ nfactor = {1.0558484276676+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 3.25460013550817e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.69005369309008 leta0 = -1.00773646981345e-7
+ etab = -0.000888016959806824 letab = 2.12632524784841e-10 petab = -1.97215226305253e-31
+ dsub = 0.0736027190697197 ldsub = 1.08667343496583e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.39323656036828 lpclm = 1.15660244945735e-7
+ pdiblc1 = -0.0118904061009604 lpdiblc1 = 1.01259257184685e-7
+ pdiblc2 = -0.00670127403829537 lpdiblc2 = 3.671552651296e-09 wpdiblc2 = 8.27180612553028e-25 ppdiblc2 = -7.88860905221012e-31
+ pdiblcb = -0.3267414016206 lpdiblcb = 5.12505014625497e-8
+ drout = 1.42027122291192 ldrout = -2.1170448393109e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 9.4214289604588e-09 lpscbe2 = -4.94566875149892e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.85667561380121 lbeta0 = -2.37001900228421e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.18294243160052e-09 lagidl = 1.2041744526071e-15 wagidl = 3.94430452610506e-31 pagidl = -2.82118644197349e-37
+ bgidl = 1000000000.0
+ cgidl = 542.793556452932 lcgidl = -0.000122303126572705
+ egidl = -1.1847845559968 legidl = 6.47188378745936e-07 wegidl = 2.11758236813575e-22 pegidl = 3.53409685539013e-28
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.48234579964 lkt1 = -1.31545844899438e-8
+ kt2 = -0.049437395288 lkt2 = -2.8967693633899e-9
+ at = 91814.8633720001 lat = -0.00903438253096768
+ ute = -0.33552325116 lute = 9.01342108658023e-9
+ ua1 = 9.1578010896e-10 lua1 = -1.81127329696748e-16
+ ub1 = 4.4238822312e-19 lub1 = -1.2607541916907e-26
+ uc1 = 4.83937303206e-11 luc1 = -1.21267323955868e-17 puc1 = -1.17549435082229e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.34 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 2e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.820095208414285+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -4.27344201774182e-8
+ k1 = 0.0701941680580003 lk1 = 1.77757512629699e-7
+ k2 = 0.162224982903557 lk2 = -6.23989353116592e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 273118.252085714 lvsat = -0.0342730489374645
+ ua = -1.22673545492428e-09 lua = -1.86112938577496e-16
+ ub = 1.10585083674714e-18 lub = 1.67826786479138e-25
+ uc = -2.39823486899798e-11 luc = 4.45271268728026e-18
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00664689435399999 lu0 = -5.84510592873481e-10
+ a0 = -0.522666542999999 la0 = 2.59715146985019e-7
+ keta = -0.342131552121685 lketa = 6.72511824073267e-08 wketa = -2.11758236813575e-22 pketa = -5.04870979341448e-29
+ a1 = 0.0
+ a2 = 1.136292205623 la2 = -8.53284302093407e-8
+ ags = -0.00199238580785632 lags = 2.30032317021635e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.156167540895428+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -5.62333475381002e-8
+ nfactor = {1.07898584053714+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 3.1958928837119e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.583915256432428 leta0 = -7.38428230328893e-8
+ etab = 0.205478856861974 letab = -5.2149453470637e-08 wetab = -6.57608586979657e-23 petab = 4.43734259186819e-30
+ dsub = 1.10602094249843 ldsub = -1.53291229588654e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.42174420808857 lpclm = -1.45306086033278e-7
+ pdiblc1 = 0.928901872578856 lpdiblc1 = -1.37450790061581e-7
+ pdiblc2 = 0.0175910419228257 lpdiblc2 = -2.49220955446714e-9
+ pdiblcb = -0.451700469176725 lpdiblcb = 8.29567405507681e-8
+ drout = -0.500968653256857 ldrout = 2.75777473568842e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 8.56916195924999e-09 lpscbe2 = 1.66791575502721e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.8201862767457 lbeta0 = -2.27743351269319e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 8.49830715721771e-09 lagidl = -1.50601104931252e-15
+ bgidl = 1000000000.0
+ cgidl = -567.119844474757 lcgidl = 0.000159318530384881 pcgidl = -5.16987882845642e-26
+ egidl = 4.68851627141714 legidl = -8.43061860096286e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.366704246714286 lkt1 = -4.24966626384441e-8
+ kt2 = 0.0995344099714284 lkt2 = -4.06958324272805e-8
+ at = 24428.4405142858 lat = 0.00806377669998873
+ ute = -0.3
+ ua1 = 3.78602403285714e-10 lua1 = -4.48276189028941e-17
+ ub1 = 3.927e-19
+ uc1 = 6.0045e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.35 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 2e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.208875994416047+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -2.31790386187043e-07 wvth0 = -2.7834695671045e-06 pvth0 = 5.11415213972811e-13
+ k1 = 1.15643073584539 lk1 = -2.18199906795816e-08 wk1 = -4.69553977027035e-06 pk1 = 8.62725608611082e-13
+ k2 = 0.119823736710078 lk2 = -5.46084271447928e-08 wk2 = 8.55648956492103e-07 pk2 = -1.57210949723163e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 222186.466857196 lvsat = -0.0249151992420732 wvsat = 0.14450696133806 pvsat = -2.65506975275258e-8
+ ua = -4.05291913092332e-09 lua = 3.33150266764836e-16 wua = 9.75650589396231e-15 pua = -1.79259209741538e-21
+ ub = 2.32313606196624e-18 lub = -5.5828679806043e-26 wub = -5.06818674209617e-24 pub = 9.31193154685556e-31
+ uc = -4.31995271148543e-13 luc = 1.25735602578125e-19 wuc = 2.93320312104815e-18 puc = -5.3892620903954e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.00660879931834962 lu0 = 1.85099777262833e-09 wu0 = 3.92186785035768e-08 pu0 = -7.20576545749768e-15
+ a0 = -1.80848854444369 la0 = 4.95963080776273e-07 wa0 = 8.81801657979073e-06 pa0 = -1.62016064025469e-12
+ keta = -0.479725425066231 lketa = 9.25317174650468e-08 wketa = 1.67604773680531e-06 pketa = -3.0794527882645e-13
+ a1 = 0.0
+ a2 = -1.00700626312034 la2 = 3.08466227348278e-7
+ ags = -11.0894596329466 lags = 2.26716593674017e-06 wags = 3.73938958022814e-05 pags = -6.87049265744057e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.0341360153477357+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -9.11983908373257e-08 wvoff = -1.72072129296795e-06 pvoff = 3.1615328532088e-13
+ nfactor = {-13.6996854751647+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 3.03491890521903e-06 wnfactor = 3.48415333207382e-05 pnfactor = -6.40153944161919e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -1.09769099009137 leta0 = 2.35123737459668e-07 weta0 = 1.56806701464535e-06 peta0 = -2.88105656801834e-13
+ etab = -0.26413953704898 letab = 3.41349428978042e-08 wetab = -4.3803329755053e-07 petab = 8.04811718588515e-14
+ dsub = 0.334801623211045 ldsub = -1.1592790398025e-08 wdsub = -9.42590247052046e-09 pdsub = 1.73184933861628e-15
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.55264404279076 lpclm = -3.53089705362615e-07 wpclm = -2.91202463736455e-06 ppclm = 5.35035022696901e-13
+ pdiblc1 = 1.007378139765 lpdiblc1 = -1.51869470060493e-7
+ pdiblc2 = 0.0224580053713133 lpdiblc2 = -3.38643134974811e-9
+ pdiblcb = -0.260549789124617 lpdiblcb = 4.78360526527541e-08 wpdiblcb = 7.86743538754726e-07 ppdiblcb = -1.44550750606022e-13
+ drout = 1.0
+ pscbe1 = 606504475.033627 lpscbe1 = 35.5515132886462 wpscbe1 = 586.375069413996 ppscbe1 = -0.000107736450628642
+ pscbe2 = 6.35212816725501e-09 lpscbe2 = 5.74133845207332e-16 wpscbe2 = 8.20098289075684e-15 ppscbe2 = -1.50679118946743e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 15.3789648910716 lbeta0 = -1.24907442241526e-06 wbeta0 = -1.99250284721502e-06 pbeta0 = 3.6608852562735e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -8.33768970119201e-10 lagidl = 2.08599293791471e-16 wagidl = 3.90615748738873e-15 pagidl = -7.17690033630394e-22
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.254505027900745 lkt1 = -6.31113617087124e-08 wkt1 = 4.65398810680724e-07 pkt1 = -8.55091196828018e-14
+ kt2 = -0.101566563684363 lkt2 = -3.74694723458086e-09 wkt2 = -6.18009260795552e-08 pkt2 = 1.13548695513748e-14
+ at = 97661.7376020369 lat = -0.00539159667383504 wat = 0.381872967219124 pat = -7.01626658860714e-8
+ ute = 0.61114960110219 lute = -1.67408249659309e-07 wute = -2.76117709019724e-06 pute = 5.07319350313209e-13
+ ua1 = 1.39406214645506e-10 lua1 = -8.79385575462877e-19 wua1 = -1.45042989778545e-17 pua1 = 2.66491836409807e-24
+ ub1 = 2.98744525545817e-19 lub1 = 1.72627211878903e-26 wub1 = 2.84725695152235e-25 pub1 = -5.23135061474055e-32
+ uc1 = -5.19106655453149e-10 luc1 = 9.54873456062233e-17 wuc1 = 9.94383206836978e-16 puc1 = -1.82701009741778e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.36 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.037561+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.42302944
+ k2 = 0.022723964
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 53438.0
+ ua = -2.0953977e-10
+ ub = 8.0838962e-19
+ uc = -9.8608028e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0120436
+ a0 = 1.061996
+ keta = 4.9707517e-6
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.17852213
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.28699958+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.731487+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.14877095
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00019189
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 757128280.0
+ pscbe2 = 9.873241e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.7815831e-11
+ alpha1 = 6.3056523e-17
+ beta0 = 9.6797043
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1352540500.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.4443203
+ kt2 = -0.052664618
+ at = 90000.0
+ ute = -0.17124159
+ ua1 = 2.1098632e-9
+ ub1 = -7.3847396e-19
+ uc1 = 1.1059776e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.37 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.037561+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.42302944
+ k2 = 0.022723964
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 53438.0
+ ua = -2.0953977e-10
+ ub = 8.0838962e-19
+ uc = -9.8608028e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0120436
+ a0 = 1.061996
+ keta = 4.9707517e-6
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.17852213
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.28699958+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.731487+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.14877095
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00019189
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 757128280.0
+ pscbe2 = 9.873241e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.7815831e-11
+ alpha1 = 6.3056523e-17
+ beta0 = 9.6797043
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1352540500.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.4443203
+ kt2 = -0.052664618
+ at = 90000.0
+ ute = -0.17124159
+ ua1 = 2.1098632e-9
+ ub1 = -7.3847396e-19
+ uc1 = 1.1059776e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.38 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.04284893035975+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.23231827220363e-8
+ k1 = 0.390585680091792 lk1 = 2.59671191821396e-7
+ k2 = 0.0350397299721097 lk2 = -9.85721025312519e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 77075.9045060112 lvsat = -0.189191476345611
+ ua = -1.32225313558197e-10 lua = -6.18804266400319e-16
+ ub = 8.10339998493619e-19 lub = -1.56103087118768e-26
+ uc = -1.11992308233283e-10 luc = 1.07124205384377e-16
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.012472700084275 lu0 = -3.4344025048146e-9
+ a0 = 1.05106881170975 la0 = 8.74582975158916e-8
+ keta = 0.00970872488828937 lketa = -7.76662572069069e-08 wketa = -4.04543018326715e-24 pketa = 2.73143088432775e-29
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.00958540767898786 lags = 1.50556250687006e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.295126527402052+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 6.50459171110729e-8
+ nfactor = {1.72539381884062+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.87681951202645e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.115420326624587 lpclm = 2.11451643903234e-06 ppclm = 1.61558713389263e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0001687584325925 lpdiblc2 = 1.85138889401132e-10
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 714216549.96731 lpscbe1 = 343.45402974973
+ pscbe2 = 1.02355866437794e-08 lpscbe2 = -2.90011778652299e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.1074273105783e-11 lalpha0 = -2.60797006106449e-17
+ alpha1 = -8.86104341585482e-13 lalpha1 = 7.09264724776501e-18 walpha1 = 5.73077005912882e-34 palpha1 = -1.75850625846278e-39
+ beta0 = 16.365642434038 lbeta0 = -5.35124636793582e-05 wbeta0 = -2.71050543121376e-20 pbeta0 = 1.03397576569128e-25
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.42279568675575e-11 lagidl = 2.86309882096554e-16
+ bgidl = 1705410008.42162 lbgidl = -2824.27332924795 wbgidl = -3.63797880709171e-12
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.435764933148282 lkt1 = -6.84748719981998e-8
+ kt2 = -0.0539027894461152 lkt2 = 9.90999366293017e-9
+ at = 133719.032745477 lat = -0.349915465113059 wat = -2.22044604925031e-16
+ ute = -0.18690663577313 lute = 1.2537884380091e-7
+ ua1 = 2.03831709184995e-09 lua1 = 5.72635946822126e-16
+ ub1 = -5.53584973233049e-19 lub1 = -1.4798020847232e-24
+ uc1 = 3.51762066741712e-10 luc1 = -1.93021472029077e-15 puc1 = -1.50463276905253e-36
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.39 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.04012695277694+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.1425111248497e-8
+ k1 = 0.397576112770504 lk1 = 2.31683365821358e-7
+ k2 = 0.031763609522666 lk2 = -8.54553909758389e-08 wk2 = 2.64697796016969e-23
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 35040.0931743605 lvsat = -0.0208913113353069
+ ua = 2.32925717519395e-10 lua = -2.0807714995097e-15 pua = -1.50463276905253e-36
+ ub = 5.44527038240346e-19 lub = 1.04863381208185e-24
+ uc = -1.06002504044869e-10 luc = 8.3142628691682e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.01400064469645 lu0 = -9.55188477075184e-9
+ a0 = 1.2580008228095 la0 = -7.4104222408055e-7
+ keta = 0.0024297412604903 lketa = -4.8523150249828e-08 pketa = -5.04870979341448e-29
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.0980562784389951 lags = 1.07459393598385e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.280414979310016+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 6.14480653389497e-9
+ nfactor = {1.8498532779084+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.49534248311533e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.409644848561555 lpclm = 1.22956699888001e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000215
+ pdiblcb = -0.0487065012492108 lpdiblcb = 9.49145013660063e-8
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 9.99009122335236e-09 lpscbe2 = -1.91721967041056e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.1379004976454e-11 lalpha0 = 1.43891889805384e-16 palpha0 = -9.4039548065783e-38
+ alpha1 = -9.8414188973042e-11 lalpha1 = 3.9756905811352e-16 walpha1 = -5.23852944873328e-32 palpha1 = 2.4685381367268e-37
+ beta0 = -0.523334251578298 lbeta0 = 1.41064896130743e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.12521285449025e-10 lagidl = 9.29562887750888e-17
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.431064760648384 lkt1 = -8.72931077417295e-8
+ kt2 = -0.0466452924507665 lkt2 = -1.91470865547484e-8
+ at = 65453.102180045 lat = -0.0765969061325282
+ ute = 0.737581701268526 lute = -3.57602561932788e-06 wute = -4.2351647362715e-22 pute = 3.23117426778526e-27
+ ua1 = 4.5429549373179e-09 lua1 = -9.45526524812681e-15
+ ub1 = -2.46394157406524e-18 lub1 = 6.16875567979646e-24
+ uc1 = -2.71048520013885e-10 luc1 = 5.63352578651982e-16 puc1 = -7.52316384526264e-37
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.40 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.04799142685194+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.71834174802088e-8
+ k1 = 0.545745111699301 lk1 = -6.52077469092329e-8
+ k2 = -0.0240934241905149 lk2 = 2.64671907573741e-08 pk2 = 5.04870979341448e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -35070.0515638739 lvsat = 0.11959069931147 pvsat = -1.05879118406788e-22
+ ua = -2.48407768102012e-10 lua = -1.11630771036507e-15
+ ub = 7.28018172120341e-19 lub = 6.80966571919086e-25
+ uc = -9.9048654346014e-11 luc = 6.92089705730477e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0115959859888 lu0 = -4.73359076449619e-9
+ a0 = 0.768645474360001 la0 = 2.39495236334215e-7
+ keta = -0.0357135328598723 lketa = 2.79057868331885e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.586225621459881 lags = 9.64329137845803e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.26875842324731+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.72118195152978e-8
+ nfactor = {1.7989321963259+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.47501996748984e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.33153053 leta0 = 8.24597303468489e-07 weta0 = 2.11758236813575e-22 peta0 = 2.01948391736579e-28
+ etab = 22.718330456674 letab = -4.56617297509427e-05 wetab = -6.35274710440725e-21 petab = -3.25136910695892e-26
+ dsub = 0.861119900000001 ldsub = -6.033638805867e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.203768610360041 lpclm = 4.24816682389036e-7
+ pdiblc1 = 0.403950724369721 lpdiblc1 = -2.79535267935121e-8
+ pdiblc2 = -8.02594999999625e-07 lpdiblc2 = 4.32410781087135e-10
+ pdiblcb = -0.00190032504012002 lpdiblcb = 1.12742149203631e-9
+ drout = 0.359844759334281 ldrout = 4.01057660844845e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.07053034974741e-08 lpscbe2 = -3.35031410607337e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 6.80772026899032e-13 lalpha0 = 9.96899866511246e-17
+ alpha1 = 1.0e-10
+ beta0 = 4.1476460511977 lbeta0 = 4.74709223805209e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.1804560163172e-10 lagidl = -1.18486265862611e-16
+ bgidl = 800836588.0609 lbgidl = 399.070300894969
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.499763474320001 lkt1 = 5.03607718996376e-8
+ kt2 = -0.0622294203980002 lkt2 = 1.20793448893456e-8
+ at = -10481.237611 lat = 0.0755552363400018
+ ute = -1.68974005325 lute = 1.28767908181878e-06 wute = -3.3881317890172e-21
+ ua1 = -6.05507873320001e-10 lua1 = 8.60879584821103e-16 wua1 = 7.88860905221012e-31
+ ub1 = 7.1724140061e-19 lub1 = -2.05485625598477e-25
+ uc1 = -7.4568904681e-11 luc1 = 1.69659889582174e-16 wuc1 = -2.46519032881566e-32 puc1 = -9.4039548065783e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.41 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.02472089008434+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.38260117988547e-8
+ k1 = 0.51109806814566 lk1 = -3.04313659420077e-8
+ k2 = -0.014602093060032 lk2 = 1.69404284877811e-08 wk2 = -1.32348898008484e-23 pk2 = 6.31088724176809e-30
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 50596.6484282161 lvsat = 0.0336042055283096
+ ua = -1.5067678703996e-09 lua = 1.46749850194403e-16
+ ub = 1.4788759087153e-18 lub = -7.26941166065852e-26
+ uc = -5.32087708585482e-11 luc = 2.31979668005231e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0064056850072 lu0 = 4.76085610668126e-10
+ a0 = 1.0094160519 la0 = -2.1741377717413e-9
+ keta = -0.0033929188485374 lketa = -4.5354800302507e-9
+ a1 = 0.0
+ a2 = 0.758500349706742 la2 = 4.16545684878049e-8
+ ags = 0.359633203042339 lags = 3.23871201700074e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.261641774077761+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.43550351361974e-8
+ nfactor = {1.2016398078014+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.52020084261877e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = -45.7167141515032 letab = 2.30287828787567e-5
+ dsub = 0.23045423603654 ldsub = 2.96560583003356e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.63119896752364 lpclm = -4.20927229785624e-9
+ pdiblc1 = 0.564470956764101 lpdiblc1 = -1.8907298121542e-7
+ pdiblc2 = 0.00027141082767328 lpdiblc2 = 1.59181185707015e-10
+ pdiblcb = 0.225119855077083 lpdiblcb = -2.26740224957544e-07 wpdiblcb = 8.27180612553028e-23 ppdiblcb = -7.25752032803331e-29
+ drout = 0.517025441331441 ldrout = 2.43290223361789e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 5.39704860466602e-09 lpscbe2 = 1.97775650224958e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.3641811504408 lbeta0 = 5.14816813283503e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -8.36202541933982e-12 lagidl = 1.08766540860231e-16
+ bgidl = 1398326823.8782 lbgidl = -200.650365972637
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.390280476580001 lkt1 = -5.95309258709272e-8
+ kt2 = -0.0451647222620002 lkt2 = -5.04905576479592e-9
+ at = 55638.1564580002 lat = 0.0091890185729423
+ ute = -0.49673611652 lute = 9.02216613929696e-8
+ ua1 = -5.41399626399993e-11 lua1 = 3.07453417730535e-16
+ ub1 = 6.0839046456e-19 lub1 = -9.62283490042024e-26
+ uc1 = 1.6512366524e-10 luc1 = -7.0927452702341e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.42 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.966160314527999+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -5.67288260786673e-9
+ k1 = 0.125830030982599 lk1 = 1.63640858222252e-7
+ k2 = 0.123287904275852 lk2 = -5.25193135402158e-08 wk2 = 5.29395592033938e-23 pk2 = 1.26217744835362e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 96261.370048 lvsat = 0.0106013783126108
+ ua = -4.59530574815197e-10 lua = -3.80778134422215e-16
+ ub = 8.95387378715198e-19 lub = 2.21228311075956e-25
+ uc = -7.890585509966e-12 luc = 3.69701340325802e-19
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0104032587366 lu0 = -1.53762419676373e-9
+ a0 = 1.51681856508 la0 = -2.57769527943444e-7
+ keta = 0.0532571099463361 lketa = -3.30719689851787e-08 wketa = -5.29395592033938e-23 pketa = 2.52435489670724e-29
+ a1 = 0.0
+ a2 = 0.882999300586521 la2 = -2.10596615357197e-8
+ ags = 1.102014123899 lags = -5.00905667058152e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.241177698902359+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -3.46634651165276e-8
+ nfactor = {1.0558484276676+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 3.25460013550817e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.69005369309008 leta0 = -1.00773646981345e-7
+ etab = -0.000888016959806824 letab = 2.12632524784841e-10
+ dsub = 0.0736027190697195 ldsub = 1.08667343496583e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.39323656036828 lpclm = 1.15660244945735e-7
+ pdiblc1 = -0.0118904061009601 lpdiblc1 = 1.01259257184685e-7
+ pdiblc2 = -0.00670127403829537 lpdiblc2 = 3.671552651296e-09 wpdiblc2 = 4.96308367531817e-24 ppdiblc2 = 2.36658271566304e-30
+ pdiblcb = -0.3267414016206 lpdiblcb = 5.12505014625496e-8
+ drout = 1.42027122291192 ldrout = -2.1170448393109e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 9.42142896045879e-09 lpscbe2 = -4.9456687514986e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.8566756138012 lbeta0 = -2.3700190022842e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.18294243160052e-09 lagidl = 1.20417445260709e-15 wagidl = 7.88860905221012e-31 pagidl = -5.64237288394698e-37
+ bgidl = 1000000000.0
+ cgidl = 542.793556452932 lcgidl = -0.000122303126572705
+ egidl = -1.1847845559968 legidl = 6.47188378745937e-07 wegidl = 8.470329472543e-22
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.482345799639999 lkt1 = -1.31545844899437e-8
+ kt2 = -0.049437395288 lkt2 = -2.8967693633899e-9
+ at = 91814.8633720001 lat = -0.00903438253096769
+ ute = -0.33552325116 lute = 9.01342108658045e-9
+ ua1 = 9.15780108959999e-10 lua1 = -1.81127329696748e-16
+ ub1 = 4.4238822312e-19 lub1 = -1.2607541916907e-26
+ uc1 = 4.83937303206e-11 luc1 = -1.21267323955868e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.43 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.820095208414287+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -4.27344201774174e-8
+ k1 = 0.070194168058002 lk1 = 1.77757512629699e-7
+ k2 = 0.162224982903557 lk2 = -6.23989353116592e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 273118.252085715 lvsat = -0.0342730489374645
+ ua = -1.22673545492429e-09 lua = -1.86112938577496e-16
+ ub = 1.10585083674714e-18 lub = 1.67826786479138e-25
+ uc = -2.39823486899799e-11 luc = 4.45271268728026e-18
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00664689435400001 lu0 = -5.84510592873479e-10
+ a0 = -0.522666542999998 la0 = 2.59715146985019e-7
+ keta = -0.342131552121685 lketa = 6.72511824073267e-08 wketa = 4.2351647362715e-22
+ a1 = 0.0
+ a2 = 1.136292205623 la2 = -8.53284302093402e-8
+ ags = -0.00199238580785632 lags = 2.30032317021635e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.15616754089543+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -5.62333475381003e-8
+ nfactor = {1.07898584053715+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 3.19589288371187e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.583915256432428 leta0 = -7.38428230328895e-8
+ etab = 0.205478856861974 letab = -5.2149453470637e-08 wetab = -9.05762770745565e-23 petab = 1.5580002878115e-29
+ dsub = 1.10602094249843 ldsub = -1.53291229588654e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.42174420808857 lpclm = -1.45306086033277e-7
+ pdiblc1 = 0.928901872578858 lpdiblc1 = -1.37450790061581e-07 wpdiblc1 = 1.6940658945086e-21
+ pdiblc2 = 0.0175910419228257 lpdiblc2 = -2.49220955446714e-9
+ pdiblcb = -0.451700469176726 lpdiblcb = 8.29567405507681e-8
+ drout = -0.500968653256855 ldrout = 2.75777473568842e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 8.56916195925002e-09 lpscbe2 = 1.66791575502718e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.82018627674574 lbeta0 = -2.27743351269322e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 8.49830715721772e-09 lagidl = -1.50601104931252e-15
+ bgidl = 1000000000.0
+ cgidl = -567.119844474757 lcgidl = 0.00015931853038488 pcgidl = -5.16987882845642e-26
+ egidl = 4.68851627141714 legidl = -8.43061860096286e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.366704246714288 lkt1 = -4.24966626384439e-8
+ kt2 = 0.0995344099714282 lkt2 = -4.06958324272804e-8
+ at = 24428.4405142858 lat = 0.00806377669998876
+ ute = -0.3
+ ua1 = 3.78602403285715e-10 lua1 = -4.48276189028941e-17
+ ub1 = 3.927e-19
+ uc1 = 6.0045e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.44 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.02951871587319+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 3.63209589118529e-07 wvth0 = 3.79187132897642e-06 pvth0 = -6.96691894886828e-13
+ k1 = -4.99841257623531 lk1 = 1.10902783557894e-06 wk1 = 7.80145227653297e-06 pk1 = -1.43338423112423e-12
+ k2 = 1.29980005899153 lk2 = -2.71409016766532e-07 wk2 = -1.54021296350575e-06 pk2 = 2.82987948423801e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 497721.103229597 lvsat = -0.0755400045866835 wvsat = -0.414947436567754 pvsat = 7.62395373629031e-8
+ ua = 8.69448233649641e-09 lua = -2.0089680470486e-15 wua = -1.6126228511814e-14 pua = 2.96292034316113e-21
+ ub = -2.95927250641151e-18 lub = 9.14724093687709e-25 wub = 5.65738570869396e-24 pub = -1.03944844841547e-30
+ uc = 6.73463650189835e-13 luc = -7.73736814161388e-20 wuc = 6.88643731385437e-19 puc = -1.26526578698641e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0430767969287639 lu0 = -7.27788588264258e-09 wu0 = -6.16645559927617e-08 pu0 = 1.13298138662181e-14
+ a0 = 9.07418202811084 la0 = -1.50354263153089e-06 wa0 = -1.32785081727164e-05 pa0 = 2.43970014209771e-12
+ keta = 2.17409332885046 lketa = -3.95062363648329e-07 wketa = -3.71235131411102e-06 pketa = 6.82081443995561e-13
+ a1 = 0.0
+ a2 = -1.00700626312033 la2 = 3.08466227348278e-7
+ ags = 39.8108113529578 lags = -7.08489355231299e-06 wags = -6.59556533962246e-05 pags = 1.21182300654485e-11
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-2.63327789597624+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 3.98893569331962e-07 wvoff = 3.6952818033122e-06 pvoff = -6.7894521156796e-13
+ nfactor = {36.2325711572154+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -6.13928440261805e-06 wnfactor = -6.65425283643098e-05 pnfactor = 1.22260583639597e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.222017693822973 leta0 = -7.35029816196609e-09 weta0 = -1.11151199179395e-06 peta0 = 2.04221432788278e-13
+ etab = -1.44781488319242 letab = 2.51615165270777e-07 wetab = 1.96533923960526e-06 petab = -3.61097674510392e-13
+ dsub = 0.32197116038436 ldsub = -9.23541097148937e-09 wdsub = 1.66254823936906e-08 pdsub = -3.0546497566396e-15
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.40870440954069 lpclm = 1.910077298296e-07 wpclm = 3.10079261566939e-06 ppclm = -5.69717929654785e-13
+ pdiblc1 = 1.007378139765 lpdiblc1 = -1.51869470060493e-7
+ pdiblc2 = 0.0224580053713133 lpdiblc2 = -3.38643134974811e-9
+ pdiblcb = 0.811027924477753 lpdiblcb = -1.4904813540055e-07 wpdiblcb = -1.38902235574591e-06 ppdiblcb = 2.55209244488262e-13
+ drout = 1.0
+ pscbe1 = 1404673515.51991 lpscbe1 = -111.098479027019 wpscbe1 = -1034.25305143245 ppscbe1 = 0.000190026415898837
+ pscbe2 = 1.10517844909409e-08 lpscbe2 = -2.89348110112432e-16 wpscbe2 = -1.34135063778841e-15 ppscbe2 = 2.46450376732787e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 16.922391402336 lbeta0 = -1.53265280560938e-06 wbeta0 = -5.12632573401966e-06 pbeta0 = 9.41875206088639e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 4.77162058812081e-09 lagidl = -8.2129574591264e-16 wagidl = -7.47520596520556e-15 pagidl = 1.37344201760511e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.0252933306666669 lkt1 = -1.05225114476621e-7
+ kt2 = -0.132003889333333 lkt2 = 1.8453939188814e-9
+ at = 651017.656601777 lat = -0.107061339739414 wat = -0.741678708778541 pat = 1.36270854200008e-7
+ ute = -0.748746627000003 lute = 8.2449564018591e-8
+ ua1 = 9.4439440091532e-10 lua1 = -1.48782280003374e-16 wua1 = -1.64897823299968e-15 pua1 = 3.0297171768373e-22
+ ub1 = 3.46882026435061e-20 lub1 = 6.57785815637008e-26 wub1 = 8.20874155786687e-25 pub1 = -1.50821671265156e-31
+ uc1 = -2.93669799116667e-11 luc1 = 5.50600579996025e-18 wuc1 = 6.16297582203915e-33 puc1 = 2.93873587705572e-39
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.45 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.037561+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.42302944
+ k2 = 0.022723964
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 53438.0
+ ua = -2.0953977e-10
+ ub = 8.0838962e-19
+ uc = -9.8608028e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0120436
+ a0 = 1.061996
+ keta = 4.9707517e-6
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.17852213
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.28699958+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.731487+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.14877095
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00019189
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 757128280.0
+ pscbe2 = 9.873241e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.7815831e-11
+ alpha1 = 6.3056523e-17
+ beta0 = 9.6797043
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1352540500.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.4443203
+ kt2 = -0.052664618
+ at = 90000.0
+ ute = -0.17124159
+ ua1 = 2.1098632e-9
+ ub1 = -7.3847396e-19
+ uc1 = 1.1059776e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.46 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.037561+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.42302944
+ k2 = 0.022723964
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 53438.0
+ ua = -2.0953977e-10
+ ub = 8.0838962e-19
+ uc = -9.8608028e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0120436
+ a0 = 1.061996
+ keta = 4.9707517e-6
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.17852213
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.28699958+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.731487+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.14877095
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00019189
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 757128280.0
+ pscbe2 = 9.873241e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.7815831e-11
+ alpha1 = 6.3056523e-17
+ beta0 = 9.6797043
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1352540500.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.4443203
+ kt2 = -0.052664618
+ at = 90000.0
+ ute = -0.17124159
+ ua1 = 2.1098632e-9
+ ub1 = -7.3847396e-19
+ uc1 = 1.1059776e-10
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.47 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.04284893035975+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.23231827220228e-8
+ k1 = 0.390585680091796 lk1 = 2.596711918214e-7
+ k2 = 0.0350397299721097 lk2 = -9.85721025312506e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 77075.9045060119 lvsat = -0.189191476345606
+ ua = -1.32225313558196e-10 lua = -6.18804266400337e-16
+ ub = 8.10339998493616e-19 lub = -1.56103087118886e-26
+ uc = -1.11992308233285e-10 luc = 1.07124205384379e-16
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0124727000842748 lu0 = -3.43440250481375e-9
+ a0 = 1.05106881170974 la0 = 8.74582975158916e-8
+ keta = 0.00970872488828944 lketa = -7.76662572069065e-08 wketa = 3.7843513024301e-23 pketa = 3.09233474846637e-28
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.00958540767899052 lags = 1.50556250687004e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.295126527402061+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 6.50459171110899e-8
+ nfactor = {1.72539381884062+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.87681951202509e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.115420326624591 lpclm = 2.11451643903234e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000168758432592502 lpdiblc2 = 1.85138889401121e-10
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 714216549.967316 lpscbe1 = 343.454029749788
+ pscbe2 = 1.02355866437794e-08 lpscbe2 = -2.90011778652339e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.10742731057832e-11 lalpha0 = -2.60797006106445e-17 walpha0 = -3.94430452610506e-31
+ alpha1 = -8.86104341585485e-13 lalpha1 = 7.09264724776499e-18 walpha1 = -5.10672361816428e-33 palpha1 = 4.54470911611859e-38
+ beta0 = 16.3656424340381 lbeta0 = -5.35124636793583e-05 wbeta0 = 2.16840434497101e-19
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.42279568675583e-11 lagidl = 2.86309882096552e-16
+ bgidl = 1705410008.42163 lbgidl = -2824.27332924795
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.435764933148285 lkt1 = -6.84748719981829e-8
+ kt2 = -0.0539027894461155 lkt2 = 9.90999366293186e-9
+ at = 133719.032745479 lat = -0.349915465113064
+ ute = -0.186906635773127 lute = 1.2537884380091e-7
+ ua1 = 2.03831709184994e-09 lua1 = 5.7263594682176e-16
+ ub1 = -5.53584973233049e-19 lub1 = -1.47980208472318e-24
+ uc1 = 3.51762066741714e-10 luc1 = -1.93021472029078e-15
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.48 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.04012695277694+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.14251112485038e-8
+ k1 = 0.397576112770516 lk1 = 2.3168336582136e-7
+ k2 = 0.0317636095226659 lk2 = -8.54553909758387e-08 wk2 = 4.2351647362715e-22 pk2 = -8.07793566946316e-28
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 35040.0931743607 lvsat = -0.0208913113353066
+ ua = 2.32925717519392e-10 lua = -2.08077149950967e-15
+ ub = 5.44527038240359e-19 lub = 1.04863381208184e-24
+ uc = -1.06002504044869e-10 luc = 8.31426286916824e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.01400064469645 lu0 = -9.55188477075195e-9
+ a0 = 1.25800082280952 la0 = -7.41042224080527e-7
+ keta = 0.00242974126049034 lketa = -4.85231502498277e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.098056278438996 lags = 1.07459393598383e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.28041497931002+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 6.14480653389666e-9
+ nfactor = {1.84985327790841+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.49534248311574e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.409644848561555 lpclm = 1.229566998879e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000215
+ pdiblcb = -0.0487065012492107 lpdiblcb = 9.4914501366006e-8
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 9.99009122335228e-09 lpscbe2 = -1.91721967041076e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.13790049764537e-11 lalpha0 = 1.43891889805384e-16 palpha0 = -1.50463276905253e-36
+ alpha1 = -9.84141889730412e-11 lalpha1 = 3.9756905811352e-16 walpha1 = -5.66993775627602e-31 palpha1 = 9.4039548065783e-38
+ beta0 = -0.523334251578262 lbeta0 = 1.41064896130743e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.12521285449026e-10 lagidl = 9.29562887750873e-17
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.43106476064839 lkt1 = -8.72931077417329e-8
+ kt2 = -0.0466452924507674 lkt2 = -1.91470865547493e-8
+ at = 65453.1021800451 lat = -0.0765969061325276
+ ute = 0.737581701268525 lute = -3.57602561932787e-06 wute = -3.3881317890172e-21 pute = -1.29246970711411e-26
+ ua1 = 4.54295493731791e-09 lua1 = -9.45526524812688e-15
+ ub1 = -2.46394157406523e-18 lub1 = 6.16875567979648e-24 wub1 = -2.35098870164458e-38 pub1 = 4.48415508583941e-44
+ uc1 = -2.71048520013887e-10 luc1 = 5.63352578651987e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.49 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.04799142685194+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.71834174802004e-8
+ k1 = 0.545745111699297 lk1 = -6.52077469092346e-8
+ k2 = -0.0240934241905149 lk2 = 2.64671907573739e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -35070.0515638734 lvsat = 0.119590699311471 pvsat = 8.470329472543e-22
+ ua = -2.48407768102021e-10 lua = -1.11630771036506e-15
+ ub = 7.28018172120314e-19 lub = 6.80966571919109e-25
+ uc = -9.90486543460148e-11 luc = 6.92089705730479e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0115959859888002 lu0 = -4.73359076449638e-9
+ a0 = 0.76864547436 la0 = 2.3949523633421e-7
+ keta = -0.0357135328598726 lketa = 2.79057868331884e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.586225621459889 lags = 9.64329137845938e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.268758423247309+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.72118195152936e-8
+ nfactor = {1.79893219632589+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.47501996748981e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.331530530000002 leta0 = 8.24597303468484e-07 peta0 = 6.46234853557053e-27
+ etab = 22.718330456674 letab = -4.56617297509423e-05 wetab = 1.60936259978317e-19 petab = -3.36042123849667e-25
+ dsub = 0.861119899999998 ldsub = -6.03363880586694e-07 wdsub = 1.35525271560688e-20
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.203768610360044 lpclm = 4.24816682389034e-7
+ pdiblc1 = 0.403950724369714 lpdiblc1 = -2.79535267935121e-8
+ pdiblc2 = -8.02594999998324e-07 lpdiblc2 = 4.32410781087133e-10
+ pdiblcb = -0.00190032504012003 lpdiblcb = 1.1274214920363e-9
+ drout = 0.35984475933428 ldrout = 4.01057660844834e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.07053034974739e-08 lpscbe2 = -3.3503141060733e-15 wpscbe2 = 2.01948391736579e-28
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 6.8077202690017e-13 lalpha0 = 9.96899866511236e-17
+ alpha1 = 1.0e-10
+ beta0 = 4.14764605119763 lbeta0 = 4.74709223805209e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.18045601631723e-10 lagidl = -1.18486265862614e-16
+ bgidl = 800836588.060913 lbgidl = 399.070300894993
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.499763474319998 lkt1 = 5.03607718996401e-8
+ kt2 = -0.0622294203980003 lkt2 = 1.20793448893464e-8
+ at = -10481.237611 lat = 0.0755552363400023
+ ute = -1.68974005325001 lute = 1.28767908181876e-06 wute = -2.71050543121376e-20
+ ua1 = -6.0550787332e-10 lua1 = 8.608795848211e-16
+ ub1 = 7.17241400609996e-19 lub1 = -2.05485625598478e-25
+ uc1 = -7.45689046810001e-11 luc1 = 1.69659889582173e-16 wuc1 = -3.94430452610506e-31 puc1 = -3.76158192263132e-37
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.50 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.02472089008434+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.3826011798853e-8
+ k1 = 0.511098068145657 lk1 = -3.04313659420081e-8
+ k2 = -0.014602093060032 lk2 = 1.69404284877811e-08 pk2 = -7.57306469012171e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 50596.6484282166 lvsat = 0.0336042055283094
+ ua = -1.50676787039959e-09 lua = 1.46749850194402e-16
+ ub = 1.47887590871529e-18 lub = -7.26941166065749e-26
+ uc = -5.32087708585479e-11 luc = 2.3197966800523e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00640568500719996 lu0 = 4.7608561066814e-10
+ a0 = 1.00941605189999 la0 = -2.17413777174553e-9
+ keta = -0.00339291884853732 lketa = -4.5354800302507e-9
+ a1 = 0.0
+ a2 = 0.75850034970675 la2 = 4.16545684878066e-8
+ ags = 0.359633203042335 lags = 3.23871201700072e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.261641774077759+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.43550351361967e-8
+ nfactor = {1.2016398078014+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.52020084261874e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = -45.7167141515029 letab = 2.30287828787569e-5
+ dsub = 0.230454236036536 ldsub = 2.96560583003345e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.631198967523645 lpclm = -4.20927229785709e-9
+ pdiblc1 = 0.564470956764097 lpdiblc1 = -1.89072981215419e-7
+ pdiblc2 = 0.000271410827673277 lpdiblc2 = 1.5918118570702e-10
+ pdiblcb = 0.225119855077083 lpdiblcb = -2.26740224957545e-07 wpdiblcb = -1.64112633530521e-21 ppdiblcb = -8.07793566946316e-28
+ drout = 0.517025441331441 ldrout = 2.43290223361786e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 5.39704860466608e-09 lpscbe2 = 1.97775650224962e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.3641811504408 lbeta0 = 5.14816813283422e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -8.36202541934002e-12 lagidl = 1.08766540860229e-16
+ bgidl = 1398326823.8782 lbgidl = -200.65036597263
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.390280476579996 lkt1 = -5.95309258709255e-8
+ kt2 = -0.0451647222620002 lkt2 = -5.04905576479592e-9
+ at = 55638.1564579988 lat = 0.00918901857294285
+ ute = -0.496736116520005 lute = 9.022166139297e-8
+ ua1 = -5.41399626400005e-11 lua1 = 3.07453417730534e-16
+ ub1 = 6.08390464559995e-19 lub1 = -9.62283490042079e-26
+ uc1 = 1.65123665239999e-10 luc1 = -7.09274527023411e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.51 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.966160314527997+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -5.67288260786588e-9
+ k1 = 0.125830030982598 lk1 = 1.63640858222251e-7
+ k2 = 0.123287904275853 lk2 = -5.25193135402156e-08 pk2 = -4.03896783473158e-28
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 96261.3700479995 lvsat = 0.0106013783126104
+ ua = -4.59530574815174e-10 lua = -3.80778134422207e-16
+ ub = 8.95387378715192e-19 lub = 2.21228311075962e-25
+ uc = -7.89058550996593e-12 luc = 3.6970134032578e-19
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0104032587366 lu0 = -1.53762419676372e-9
+ a0 = 1.51681856508 la0 = -2.57769527943447e-7
+ keta = 0.0532571099463366 lketa = -3.30719689851789e-08 pketa = 1.0097419586829e-28
+ a1 = 0.0
+ a2 = 0.882999300586519 la2 = -2.10596615357202e-8
+ ags = 1.10201412389901 lags = -5.00905667058152e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.241177698902362+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -3.46634651165269e-8
+ nfactor = {1.05584842766763+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 3.25460013550819e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.690053693090078 leta0 = -1.00773646981345e-7
+ etab = -0.000888016959806823 letab = 2.12632524784841e-10
+ dsub = 0.0736027190697186 ldsub = 1.08667343496583e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.39323656036828 lpclm = 1.15660244945737e-7
+ pdiblc1 = -0.0118904061009601 lpdiblc1 = 1.01259257184685e-7
+ pdiblc2 = -0.0067012740382954 lpdiblc2 = 3.67155265129602e-09 wpdiblc2 = -5.29395592033938e-23 ppdiblc2 = 2.52435489670724e-29
+ pdiblcb = -0.326741401620598 lpdiblcb = 5.125050146255e-08 wpdiblcb = 6.7762635780344e-21
+ drout = 1.42027122291192 ldrout = -2.11704483931093e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 9.421428960459e-09 lpscbe2 = -4.94566875149545e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.85667561380137 lbeta0 = -2.37001900228447e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.18294243160054e-09 lagidl = 1.2041744526071e-15 pagidl = -9.02779661431517e-36
+ bgidl = 1000000000.0
+ cgidl = 542.79355645294 lcgidl = -0.000122303126572704
+ egidl = -1.1847845559968 legidl = 6.47188378745936e-07 wegidl = 6.7762635780344e-21 pegidl = 1.61558713389263e-27
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.482345799640001 lkt1 = -1.31545844899464e-8
+ kt2 = -0.0494373952879998 lkt2 = -2.89676936338988e-9
+ at = 91814.8633719999 lat = -0.00903438253096756
+ ute = -0.335523251159998 lute = 9.01342108658002e-9
+ ua1 = 9.15780108959991e-10 lua1 = -1.81127329696749e-16
+ ub1 = 4.42388223120001e-19 lub1 = -1.26075419169083e-26
+ uc1 = 4.83937303205998e-11 luc1 = -1.21267323955868e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.52 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.820095208414273+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -4.27344201774072e-8
+ k1 = 0.0701941680579523 lk1 = 1.77757512629699e-7
+ k2 = 0.16222498290356 lk2 = -6.23989353116595e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 273118.252085712 lvsat = -0.0342730489374645
+ ua = -1.22673545492422e-09 lua = -1.86112938577494e-16
+ ub = 1.10585083674707e-18 lub = 1.67826786479138e-25
+ uc = -2.39823486899797e-11 luc = 4.45271268728027e-18 puc = 4.70197740328915e-38
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00664689435400001 lu0 = -5.84510592873483e-10
+ a0 = -0.522666543 la0 = 2.59715146985019e-7
+ keta = -0.342131552121685 lketa = 6.7251182407327e-08 wketa = 3.3881317890172e-21 pketa = 8.07793566946316e-28
+ a1 = 0.0
+ a2 = 1.13629220562296 la2 = -8.53284302093423e-8
+ ags = -0.00199238580788119 lags = 2.30032317021627e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.156167540895424+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -5.62333475381009e-8
+ nfactor = {1.07898584053709+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 3.19589288371187e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.583915256432427 leta0 = -7.38428230328895e-8
+ etab = 0.205478856861975 letab = -5.21494534706368e-08 wetab = -1.49885126994609e-21 petab = 1.82621299558664e-28
+ dsub = 1.1060209424984 ldsub = -1.53291229588656e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.42174420808854 lpclm = -1.45306086033282e-7
+ pdiblc1 = 0.928901872578848 lpdiblc1 = -1.37450790061581e-7
+ pdiblc2 = 0.0175910419228256 lpdiblc2 = -2.49220955446717e-9
+ pdiblcb = -0.451700469176728 lpdiblcb = 8.2956740550768e-8
+ drout = -0.500968653256891 ldrout = 2.75777473568842e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 8.56916195924962e-09 lpscbe2 = 1.66791575502724e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.82018627674574 lbeta0 = -2.2774335126937e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 8.49830715721768e-09 lagidl = -1.50601104931252e-15
+ bgidl = 1000000000.0
+ cgidl = -567.119844474768 lcgidl = 0.00015931853038488 wcgidl = 3.46944695195361e-18
+ egidl = 4.68851627141714 legidl = -8.43061860096295e-7
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.366704246714264 lkt1 = -4.2496662638446e-8
+ kt2 = 0.0995344099714313 lkt2 = -4.06958324272798e-8
+ at = 24428.4405142851 lat = 0.0080637766999887
+ ute = -0.3
+ ua1 = 3.78602403285712e-10 lua1 = -4.48276189028925e-17
+ ub1 = 3.927e-19
+ uc1 = 6.0045e-13
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.53 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.58062345640172+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.03502466262007e-06 wvth0 = -9.22476088906058e-06 pvth0 = 1.69489299242978e-12
+ k1 = -0.437312594293303 lk1 = 2.71003252596805e-7
+ k2 = -1.07788640245405 lk2 = 1.65450449854247e-07 wk2 = 2.52665852165483e-06 pk2 = -4.64230550159208e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -81921.7253226042 lvsat = 0.030959511231698 wvsat = 0.576492321887002 pvsat = -1.05920663777266e-7
+ ua = 1.88357210175783e-09 lua = -7.57579076889378e-16 wua = -4.47662833500772e-15 pua = 8.22504353875938e-22
+ ub = 4.72282569583753e-18 lub = -4.96730855306083e-25 wub = -7.48232241999482e-24 pub = 1.37474954519291e-30
+ uc = 1.07607752251136e-12 luc = -1.5134713601939e-19
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0192269245310499 lu0 = -2.89587727739342e-09 wu0 = -2.08709662778205e-08 pu0 = 3.83468524712279e-15
+ a0 = 1.31093471978932 la0 = -7.71779138310601e-8
+ keta = 0.00367621783546568 lketa = 3.7148834097892e-9
+ a1 = 0.0
+ a2 = -1.0070062631203 la2 = 3.08466227348277e-7
+ ags = 1.25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.524508009358215+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 1.14429517539678e-08 wvoff = 8.83738868503298e-08 pvoff = -1.62371993526758e-14
+ nfactor = {8.15013168399594+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -9.7961355088503e-07 wnfactor = -1.85094196347643e-05 pnfactor = 3.40079119775418e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.427825072113002 leta0 = 1.12047262751746e-7
+ etab = -0.298784106289798 letab = 4.05002935381285e-8
+ dsub = 0.331691207980327 ldsub = -1.10213044764397e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.40416640502266 lpclm = -1.42076463542576e-7
+ pdiblc1 = 1.007378139765 lpdiblc1 = -1.51869470060491e-7
+ pdiblc2 = 0.0224580053713135 lpdiblc2 = -3.38643134974814e-9
+ pdiblcb = -0.00106059662580517 lpdiblcb = 1.5932484736986e-10
+ drout = 1.0
+ pscbe1 = 800000000.0
+ pscbe2 = 1.02675671230797e-08 lpscbe2 = -1.45261500463247e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 13.925297606967 lbeta0 = -9.8198777130485e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 4.01259713713989e-10 lagidl = -1.83162313752573e-17
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.0252933306666705 lkt1 = -1.0522511447662e-7
+ kt2 = -0.132003889333333 lkt2 = 1.84539391888119e-9
+ at = 217397.014533333 lat = -0.0273909183102528
+ ute = -0.748746627000003 lute = 8.24495640185907e-8
+ ua1 = -1.96766876666683e-11 lua1 = 2.83493933150585e-17
+ ub1 = 5.14610268999982e-19 lub1 = -2.23989394541766e-26
+ uc1 = -2.93669799116669e-11 luc1 = 5.50600579996025e-18 wuc1 = -9.86076131526265e-32 puc1 = 1.17549435082229e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.54 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.13096512967641+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = 1.56959307121216e-7
+ k1 = 0.19558057364442 wk1 = 3.82212398877412e-7
+ k2 = 0.106152758287165 wk2 = -1.40196432327327e-7
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 47482.7645874169 wvsat = 0.0100073693458849
+ ua = 3.73691070795186e-09 wua = -6.63174245885569e-15
+ ub = -1.41791159199137e-18 wub = 3.74114824352933e-24
+ uc = -2.96115068812591e-10 wuc = 3.31897191108192e-16
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0286798347166373 wu0 = -2.79560645045952e-8
+ a0 = 0.549753975009232 wa0 = 8.60787992987693e-7
+ keta = -0.0219498026060158 wketa = 3.68935080940078e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.173246511271507 wags = 5.9112335174289e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.295306886183523+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = 1.39598648060513e-8
+ nfactor = {2.05437034220267+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor = -5.42583565080981e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.635266257177647 wpclm = -8.17522379330209e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00105204806018602 wpdiblc2 = 2.09035357114213e-9
+ pdiblcb = 0.636760102564102 wpdiblcb = -1.11204298502402e-6
+ drout = 0.56
+ pscbe1 = 615322983.334046 wpscbe1 = 238.294186648021
+ pscbe2 = 6.89952271511282e-09 wpscbe2 = 4.9971319596532e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.67648617491236e-11 walpha0 = -9.90598494296174e-17
+ alpha1 = 2.71697978639078e-16 walpha1 = -3.50607820310779e-22
+ beta0 = -57.5561005328244 wbeta0 = 0.000112985211433994
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -5.45472558247896e-11 wagidl = 2.59706185109614e-16
+ bgidl = 2519026687.19 wbgidl = -1960.2009498093
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.109172888696564 wkt1 = -5.63192501700938e-7
+ kt2 = -0.0532622469310246 wkt2 = 1.00427489934535e-9
+ at = 354704.041025641 wat = -0.444817194009608
+ ute = 3.42958839508923 wute = -6.05095065366947e-6
+ ua1 = 9.93819800944882e-09 wua1 = -1.31549858861787e-14
+ ub1 = -4.81760942306028e-18 wub1 = 6.85471058028841e-24
+ uc1 = 4.49427733922184e-10 wuc1 = -5.69380798503999e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.55 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.13096512967641+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = 1.56959307121216e-7
+ k1 = 0.195580573644421 wk1 = 3.82212398877413e-7
+ k2 = 0.106152758287165 wk2 = -1.40196432327327e-7
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 47482.7645874169 wvsat = 0.0100073693458849
+ ua = 3.73691070795186e-09 wua = -6.6317424588557e-15
+ ub = -1.41791159199137e-18 wub = 3.74114824352933e-24
+ uc = -2.96115068812591e-10 wuc = 3.31897191108192e-16
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0286798347166373 wu0 = -2.79560645045952e-8
+ a0 = 0.549753975009232 wa0 = 8.60787992987693e-7
+ keta = -0.0219498026060158 wketa = 3.68935080940078e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.173246511271507 wags = 5.9112335174289e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.295306886183523+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = 1.39598648060508e-8
+ nfactor = {2.05437034220267+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor = -5.42583565080982e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.635266257177647 wpclm = -8.17522379330209e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00105204806018602 wpdiblc2 = 2.09035357114213e-9
+ pdiblcb = 0.636760102564102 wpdiblcb = -1.11204298502402e-6
+ drout = 0.56
+ pscbe1 = 615322983.334046 wpscbe1 = 238.294186648021
+ pscbe2 = 6.89952271511282e-09 wpscbe2 = 4.9971319596532e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.67648617491236e-11 walpha0 = -9.90598494296174e-17
+ alpha1 = 2.71697978639078e-16 walpha1 = -3.50607820310779e-22
+ beta0 = -57.5561005328244 wbeta0 = 0.000112985211433994
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -5.45472558247897e-11 wagidl = 2.59706185109614e-16
+ bgidl = 2519026687.19 wbgidl = -1960.2009498093
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.109172888696564 wkt1 = -5.63192501700938e-7
+ kt2 = -0.0532622469310247 wkt2 = 1.00427489934529e-9
+ at = 354704.041025641 wat = -0.444817194009608
+ ute = 3.42958839508923 wute = -6.05095065366947e-6
+ ua1 = 9.93819800944882e-09 wua1 = -1.31549858861787e-14
+ ub1 = -4.81760942306028e-18 wub1 = 6.85471058028841e-24
+ uc1 = 4.49427733922184e-10 wuc1 = -5.69380798503999e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.56 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.15268933315917+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.73874724313652e-07 wvth0 = 1.84579349725112e-07 pvth0 = -2.21063446450198e-13
+ k1 = -0.0833504842219526 lk1 = 2.23248971257e-06 wk1 = 7.96417591257308e-07 pk1 = -3.31518776702232e-12
+ k2 = 0.200620284903445 lk2 = -7.56092860207099e-07 wk2 = -2.78246896200484e-07 pk2 = 1.10491905336689e-12
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 107961.513457532 lvsat = -0.484055758130451 wvsat = -0.0519011717987432 pvsat = 4.95499433741118e-7
+ ua = 5.96260590324293e-09 lua = -1.78138700824926e-14 wua = -1.02419506302778e-14 pua = 2.88951422784807e-20
+ ub = -2.49963760973955e-18 lub = 8.65784622520965e-24 wub = 5.562192954154e-24 pub = -1.45751556449021e-29
+ uc = -4.05629646953081e-10 luc = 8.76525443044119e-16 wuc = 4.93437639107055e-16 puc = -1.29292661448328e-21
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0388037424036403 lu0 = -8.10290540434194e-08 wu0 = -4.42475313730242e-08 pu0 = 1.30392550993251e-13
+ a0 = 0.23032437751773 la0 = 2.55662921061944e-06 wa0 = 1.37920537518705e-06 pa0 = -4.14927430968263e-12
+ keta = 0.00854221681154138 lketa = -2.44049982048944e-07 wketa = 1.96023773372737e-09 pketa = 2.79596568780498e-13
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.789087290608182 lags = 4.92902516832266e-06 wags = 1.30990006403485e-06 pags = -5.75289689180265e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.27019923169411+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.00954962789513e-07 wvoff = -4.18886303665484e-08 pvoff = 4.46996443813276e-13
+ nfactor = {3.27343975022941+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -9.75710605031412e-06 wnfactor = -2.60138623018471e-06 pnfactor = 1.64781068311787e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.382980916699502 lpclm = 8.14977850771728e-06 wpclm = 4.49617431012888e-07 ppclm = -1.01418487156568e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000405029040398884 lpdiblc2 = -1.16620560734957e-08 wpdiblc2 = -3.9703673727142e-10 ppdiblc2 = 1.99084078953297e-14
+ pdiblcb = 0.636760102564102 wpdiblcb = -1.11204298502402e-6
+ drout = 0.56
+ pscbe1 = 430473550.60452 lpscbe1 = 1479.48550476859 wpscbe1 = 476.810872653812 ppscbe1 = -0.00190902387083518
+ pscbe2 = 4.25771064718526e-09 lpscbe2 = 2.11443584278701e-14 wpscbe2 = 1.00454153122838e-14 ppscbe2 = -4.04051120628001e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 9.08048387655173e-11 lalpha0 = -1.12372227365352e-16 walpha0 = -1.17177487858832e-16 palpha0 = 1.45008740577972e-22
+ alpha1 = -3.81804684143601e-12 lalpha1 = 3.05608020984248e-17 walpha1 = 4.92693058529732e-18 palpha1 = -3.9436643085635e-23
+ beta0 = -28.7477268721954 lbeta0 = -0.000230574530943907 wbeta0 = 7.58099584326862e-05 pbeta0 = 2.97540799229915e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.73010662274819e-10 lagidl = 9.48149475496512e-16 wagidl = 3.98663414690386e-16 pagidl = -1.1121765639842e-21
+ bgidl = 4039471006.03582 lbgidl = -12169.2303694088 wbgidl = -3922.23125715502 pbgidl = 0.015703566717903
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = 0.206982033445805 lkt1 = -2.53041958346331e-06 wkt1 = -1.08009269911703e-06 pkt1 = 4.13713116776569e-12
+ kt2 = 0.026657351810039 lkt2 = -6.39655129790609e-07 wkt2 = -1.3537585540339e-07 pkt2 = 1.0915501494483e-12
+ at = 693004.854078897 lat = -2.70766938136118 wat = -0.939841903172125 pat = 3.96204560053944e-6
+ ute = 7.3015821501731 lute = -3.09904041933586e-05 wute = -1.25838976852429e-05 pute = 5.22879637438567e-11
+ ua1 = 1.68354302101602e-08 lua1 = -5.52036049734964e-14 wua1 = -2.4865545351051e-14 pua1 = 9.37281912374608e-20
+ ub1 = -9.02138132076949e-18 lub1 = 3.36458678621678e-23 wub1 = 1.42295576454426e-23 pub1 = -5.90263068253279e-29
+ uc1 = 1.19646428936899e-09 luc1 = -5.97908113103591e-15 wuc1 = -1.41946481431444e-15 puc1 = 6.80384549011456e-21
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.57 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.12795846071278+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 7.48589141812741e-08 wvth0 = 1.47594894109938e-07 pvth0 = -7.29875610166889e-14
+ k1 = 0.262962843733705 lk1 = 8.45943613094112e-07 wk1 = 2.26208471836701e-07 pk1 = -1.0322226986971e-12
+ k2 = 0.0930776850968266 lk2 = -3.25521004455549e-07 wk2 = -1.03034146908053e-07 pk2 = 4.03413987004058e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 44986.3782493797 lvsat = -0.231920131118111 wvsat = -0.0167140577104419 pvsat = 3.54619623891021e-7
+ ua = 3.10262333166134e-09 lua = -6.36326348122651e-15 wua = -4.82233227506731e-15 pua = 7.19643742231874e-21
+ ub = -9.34731136817085e-19 lub = 2.39237853765638e-24 wub = 2.48579306947974e-24 pub = -2.2580719054356e-30
+ uc = -2.4456119525243e-10 luc = 2.3165036771132e-16 wuc = 2.32838486295044e-16 puc = -2.49557186597795e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0267858009959204 lu0 = -3.29124254372647e-08 wu0 = -2.14845883276629e-08 pu0 = 3.92558047454177e-14
+ a0 = 1.48948521864268 la0 = -2.48471460130029e-06 wa0 = -3.88993832555628e-07 pa0 = 2.9301232089306e-12
+ keta = -0.0268341771817933 lketa = -1.02412345996828e-07 wketa = 4.91760308485872e-08 pketa = 9.05571397653612e-14
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.447936202865201 lags = 3.56314730034019e-06 wags = 9.17503346541472e-07 pags = -4.18184520488274e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.332420120866248+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 4.8160864478318e-08 wvoff = 8.73911144366522e-08 pvoff = -7.06051366868769e-14
+ nfactor = {0.28001400669724+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.22777138211518e-06 wnfactor = 2.63800846016776e-06 pnfactor = -4.49903059061034e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.183540622923726 leta0 = 1.05514628884028e-06 weta0 = 4.42862148769088e-07 peta0 = -1.77310179947771e-12
+ etab = 0.160390854094634 letab = -9.22423465436873e-07 wetab = -3.87156209806126e-07 petab = 1.55007009335571e-12
+ dsub = -0.434492916693306 ldsub = 3.98168410883124e-06 wdsub = 1.67117791988335e-06 pdsub = -6.69095018670832e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.68117485306635 lpclm = -4.11828306483465e-06 wpclm = -3.817152162836e-06 ppclm = 6.9411575106326e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00523561526674618 lpdiblc2 = 1.09215776802831e-08 wpdiblc2 = 9.15938940405188e-09 ppdiblc2 = -1.83529708087491e-14
+ pdiblcb = 0.534613517824323 lpdiblcb = 4.08967652159951e-07 wpdiblcb = -9.8022974295578e-07 ppdiblcb = -5.277450271056e-13
+ drout = 0.56
+ pscbe1 = 800000132.475538 lpscbe1 = -0.000265445605691639 wpscbe1 = -0.000222616159589961 ppscbe1 = 4.46063345982406e-10
+ pscbe2 = 1.1168753746831e-08 lpscbe2 = -6.52561289460364e-15 wpscbe2 = -1.98066245738667e-15 ppscbe2 = 7.74409236419584e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -8.20105476908372e-11 lalpha0 = 5.79534438297708e-16 walpha0 = 1.01887196712925e-16 palpha0 = -7.32067766176562e-22
+ alpha1 = -4.2405680044438e-10 lalpha1 = 1.7130845677774e-15 walpha1 = 5.47220330008526e-16 palpha1 = -2.2106346220386e-21
+ beta0 = -191.02332077859 lbeta0 = 0.000419133619473724 wbeta0 = 0.000320122311459557 pbeta0 = -6.80620630891417e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.65110715812428e-10 lagidl = -8.05971543956877e-16 wagidl = -2.56416192162321e-16 pagidl = 1.51058727559901e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.363210682395961 lkt1 = -2.47520190688011e-07 wkt1 = -1.14024177996694e-07 pkt1 = 2.69250749495003e-13
+ kt2 = -0.174779778138403 lkt2 = 1.66845354809257e-07 wkt2 = 2.15321315679944e-07 pkt2 = -3.12547687424687e-13
+ at = -59333.7870843834 lat = 0.304493663439408 wat = 0.20969590685778 pat = -6.40396864225022e-7
+ ute = 0.674687178844237 lute = -4.45808610911521e-06 wute = 1.05689980685395e-07 pute = 1.4822428493864e-12
+ ua1 = 6.35146539274984e-09 lua1 = -1.32286090631915e-14 wua1 = -3.0390792033445e-15 pua1 = 6.34084844850554e-21
+ ub1 = -1.41492755423026e-18 lub1 = 3.19165790410035e-24 wub1 = -1.76279693718214e-24 pub1 = 5.00281096482813e-30
+ uc1 = -4.32907520610718e-10 luc1 = 5.44488553849572e-16 wuc1 = 2.71993076462738e-16 puc1 = 3.16997146995681e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.58 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.16184614327083+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.4276078201636e-07 wvth0 = 1.91325131592172e-07 pvth0 = -1.60611280957685e-13
+ k1 = 0.800042927328011 lk1 = -2.30221474046558e-07 wk1 = -4.27330237772149e-07 pk1 = 2.77294380523574e-13
+ k2 = -0.118599424517932 lk2 = 9.86234054241614e-08 wk2 = 1.58810926043403e-07 pk2 = -1.21253626556182e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -409713.432117915 lvsat = 0.67917688400858 wvsat = 0.629562800199865 pvsat = -9.40346643440171e-7
+ ua = 3.17707810037381e-09 lua = -6.51245095830304e-15 wua = -5.75629675403173e-15 pua = 9.06785286964756e-21
+ ub = -1.92473730551581e-18 lub = 4.37608656808158e-24 wub = 4.45777572334617e-24 pub = -6.20939862441533e-30
+ uc = -2.89891397292771e-10 luc = 3.22479989436217e-16 wuc = 3.20698290384053e-16 puc = -4.25604775424478e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0219673920086448 lu0 = -2.32576203419641e-08 wu0 = -1.74284446350211e-08 pu0 = 3.11283757757294e-14
+ a0 = -2.1946860631406 la0 = 4.89738097366116e-06 wa0 = 4.97967773489151e-06 pa0 = -7.82726117692495e-12
+ keta = -0.247639255010535 lketa = 3.40022075016191e-07 wketa = 3.56126807510227e-07 pketa = -5.24490260807197e-13
+ a1 = 0.0
+ a2 = 0.8
+ ags = 4.02162087128858 lags = -5.39265170452518e-06 wags = -5.77294879753919e-06 pags = 9.22403454113243e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.288576718625007+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -3.96896074247314e-08 wvoff = 3.3303301701792e-08 pvoff = 3.77723985877833e-14
+ nfactor = {2.18422657147463+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.58776217294391e-06 wnfactor = -6.47461074478801e-07 pnfactor = 2.08417313645563e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -1.16612171285784 leta0 = 3.02397644391724e-06 weta0 = 1.40247389751041e-06 peta0 = -3.6959075276184e-12
+ etab = 97.8688208425544 letab = -0.000196704029011503 wetab = -0.000126285303890224 petab = 2.53816343239482e-10
+ dsub = 3.84645141292708 ldsub = -4.59618531559199e-06 wdsub = -5.01664720199737e-06 pdsub = 6.7096657082331e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.224252861369861 lpclm = 1.70341832569575e-06 wpclm = 7.19261063386316e-07 ppclm = -2.14860337238552e-12
+ pdiblc1 = 0.424336521569003 lpdiblc1 = -6.88012213730229e-08 wpdiblc1 = -3.42569500363451e-08 ppdiblc1 = 6.86417812671749e-14
+ pdiblc2 = -0.000714850332003997 lpdiblc2 = 1.86317179529736e-09 wpdiblc2 = 1.19990880959865e-09 ppdiblc2 = -2.40429687878353e-15
+ pdiblcb = 1.40052244690419 lpdiblcb = -1.32608264403205e-06 wpdiblcb = -2.35667638398848e-06 ppdiblcb = 2.23028653027078e-12
+ drout = 0.864135028730798 ldrout = -6.09405393523848e-07 wdrout = -8.47425606840583e-07 pdrout = 1.6980146534715e-12
+ pscbe1 = 800000000.0
+ pscbe2 = 1.19206346111005e-08 lpscbe2 = -8.03218139440919e-15 wpscbe2 = -2.04228153699977e-15 ppscbe2 = 7.86756054744621e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.14833897541503e-10 lalpha0 = -2.15635872481026e-16 walpha0 = -5.27913027845383e-16 palpha0 = 5.2988372717833e-22
+ alpha1 = 7.63014662852583e-10 lalpha1 = -6.65489696589011e-16 walpha1 = -1.11415118852962e-15 palpha1 = 1.1183103149164e-21
+ beta0 = 27.5431844246873 lbeta0 = -1.88152996967546e-05 wbeta0 = -3.93146160191475e-05 pbeta0 = 3.95950021162695e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.75133754029893e-10 lagidl = 4.76907428333686e-16 wagidl = 9.96797689629026e-16 pagidl = -1.00051873540441e-21
+ bgidl = 141844588.501722 lbgidl = 1719.51431714768 wbgidl = 1107.39137560163 pbgidl = -0.00221891664320837
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.737435485876977 lkt1 = 5.02326397465415e-07 wkt1 = 3.99391701259115e-07 pkt1 = -7.59497590493878e-13
+ kt2 = -0.178419001103814 lkt2 = 1.74137385959408e-07 wkt2 = 1.95248712722548e-07 pkt2 = -2.72327550483055e-13
+ at = -18397.0476652952 lat = 0.22246736775298 wat = 0.0133019821043213 pat = -2.46875876197e-7
+ ute = -5.3101813035763 lute = 7.53399236977073e-06 wute = 6.08390605525657e-06 pute = -1.04965059803623e-11
+ ua1 = -2.39118691876407e-09 lua1 = 4.28933188091521e-15 wua1 = 3.00071256682948e-15 pua1 = -5.76128163452047e-21
+ ub1 = -2.66182660577006e-19 lub1 = 8.89879852105835e-25 wub1 = 1.65257745867341e-24 pub1 = -1.84068741950271e-30
+ uc1 = -5.73927101458302e-10 luc1 = 8.27054141640043e-16 wuc1 = 8.39137593198514e-16 puc1 = -1.10470646925296e-21
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.59 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.00984295615293+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -9.80983299905289e-09 wvth0 = -2.50013592478149e-08 pvth0 = 5.65227566726069e-14
+ k1 = 0.886335072031763 lk1 = -3.16835747326488e-07 wk1 = -6.30560343961732e-07 pk1 = 4.81283144699561e-13
+ k2 = -0.140330413602454 lk2 = 1.20435516290936e-07 wk2 = 2.11277918291408e-07 pk2 = -1.73916478086248e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 323513.680742197 lvsat = -0.0567873656638388 wvsat = -0.458618569028855 pvsat = 1.51896906839878e-7
+ ua = -5.15325049847805e-09 lua = 1.84897475720833e-15 wua = 6.12766682496365e-15 pua = -2.86047354538821e-21
+ ub = 3.50814664785413e-18 lub = -1.07707834108629e-24 wub = -3.4100518925667e-24 pub = 1.68779959198773e-30
+ uc = 2.14193978527617e-11 luc = 1.00070710924064e-17 wuc = -1.25407577729518e-16 puc = 2.21664058947612e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.00984879722284161 lu0 = 8.67733872392346e-09 wu0 = 2.73145553336897e-08 pu0 = -1.37816498118645e-14
+ a0 = 4.81042244136562 la0 = -2.13387760089237e-06 wa0 = -6.38733352926377e-06 pa0 = 3.58218314027942e-12
+ keta = 0.125535544892604 lketa = -3.45457864149867e-08 wketa = -2.16655541967146e-07 pketa = 5.04302851807759e-14
+ a1 = 0.0
+ a2 = 0.621186285534529 la2 = 1.7948122606157e-07 wa2 = 2.30746974947848e-07 pa2 = -2.31608353405329e-13
+ ags = -2.68841261231614 lags = 1.34243033407384e-06 wags = 5.12203433520365e-06 pags = -1.71161956364494e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.258322495173483+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.00567698923991e-08 wvoff = -5.57782315152712e-09 pvoff = 7.67986666801801e-14
+ nfactor = {0.454058274395418+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.48864842388289e-07 wnfactor = 1.25626008086078e-06 pnfactor = 1.73345390043164e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 3.21334485741059 leta0 = -1.37183867505801e-06 weta0 = -4.57639639009717e-06 peta0 = 2.30528188277282e-12
+ etab = -196.937726083154 letab = 9.92030307538784e-05 wetab = 0.00025411665776653 petab = -1.28005658940136e-10
+ dsub = -1.66859342824252 ldsub = 9.39447187969692e-07 wdsub = 3.19122084438933e-06 pdsub = -1.52884230957076e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.34044477998998 lpclm = -8.70853331959288e-07 wpclm = -2.8722717009836e-06 ppclm = 1.45633658379379e-12
+ pdiblc1 = 0.410441363260046 lpdiblc1 = -5.48541924380977e-08 wpdiblc1 = 2.58836288677125e-07 ppdiblc1 = -2.25545574506411e-13
+ pdiblc2 = 0.00151542464288602 lpdiblc2 = -3.75428796073915e-10 wpdiblc2 = -2.09048087232834e-09 ppdiblc2 = 8.9837582782609e-16
+ pdiblcb = 1.05271655982273 lpdiblcb = -9.76978397574105e-07 wpdiblcb = -1.39072015126847e-06 ppdiblcb = 1.26072438293403e-12
+ drout = -0.491555097461596 ldrout = 7.51345523909622e-07 wdrout = 1.69485121368117e-06 pdrout = -8.53752486421255e-13
+ pscbe1 = 800000000.0
+ pscbe2 = -1.54727645675521e-09 lpscbe2 = 5.48600538546286e-15 wpscbe2 = 1.16694674404792e-14 ppscbe2 = -5.89537438896565e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.02408397721993 lbeta0 = 1.7803985526831e-06 wbeta0 = 2.25194244100931e-06 pbeta0 = -2.1267243066191e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 5.61020661795334e-10 lagidl = -4.62741651925816e-16 wagidl = -9.56809001718067e-16 pagidl = 9.6038076972148e-22
+ bgidl = 2716310822.99655 lbgidl = -864.562399800522 wbgidl = -2214.78275120325 pbgidl = 0.00111565915961187
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = 0.0365322921993196 lkt1 = -2.7453060232644e-07 wkt1 = -7.17229920027923e-07 pkt1 = 3.61292379305426e-13
+ kt2 = 0.0457047270569474 lkt2 = -5.08229960785773e-08 wkt2 = -1.52699948631827e-07 pkt2 = 7.69200032241563e-14
+ at = 303970.184062551 lat = -0.101103260850906 wat = -0.417305135477977 pat = 1.85338697755233e-7
+ ute = 4.98465755369996 lute = -2.79927712095974e-06 wute = -9.2111104243138e-06 pute = 4.85560679572628e-12
+ ua1 = 3.21807465890679e-09 lua1 = -1.34086907022509e-15 wua1 = -5.49873481535804e-15 pua1 = 2.76989418474475e-21
+ ub1 = 1.27212061749461e-18 lub1 = -6.54165912102817e-25 wub1 = -1.11535352110223e-24 pub1 = 9.37576246620443e-31
+ uc1 = 4.77467567503995e-10 luc1 = -2.2826538362149e-16 wuc1 = -5.2487275083807e-16 puc1 = 2.64395725397913e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.60 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.981978318361394+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -2.38461705876974e-08 wvth0 = 2.65810829813602e-08 pvth0 = 3.05389783011791e-14
+ k1 = -0.903508253159703 lk1 = 5.84767400402184e-07 wk1 = 1.72973319736548e-06 pk1 = -7.07674601753817e-13
+ k2 = 0.508139235230788 lk2 = -2.0622004532478e-07 wk2 = -6.46716568749531e-07 pk2 = 2.58283658854345e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 320334.969845211 lvsat = -0.0551861440875674 wvsat = -0.376540492269147 pvsat = 1.10551470999481e-7
+ ua = 3.02897582694716e-10 lua = -8.99467084165071e-16 wua = -1.28120882606633e-15 pua = 8.71621612932078e-22
+ ub = 4.15510093331442e-19 lub = 4.80784748433084e-25 wub = 8.06401242407454e-25 pub = -4.36166995052202e-31
+ uc = 1.11507821781192e-10 luc = -3.53734409583336e-17 wuc = -2.00640928240777e-16 puc = 6.00639272478493e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0143839513337989 lu0 = -3.52949640475873e-09 wu0 = -6.68928401863467e-09 pu0 = 3.3472061965999e-15
+ a0 = 1.69384829980688 la0 = -5.63956358842563e-07 wa0 = -2.97486466592505e-07 pa0 = 5.14526209858835e-13
+ keta = 0.418383597390542 lketa = -1.8206301444393e-07 wketa = -6.13570306574139e-07 pketa = 2.5036935030055e-13
+ a1 = 0.0
+ a2 = 0.229832802487768 la2 = 3.76618890137164e-07 wa2 = 1.09760201536638e-06 pa2 = -6.68271843480478e-13
+ ags = -2.58668385850566 lags = 1.29118620373062e-06 wags = 6.19860686570783e-06 pags = -2.2539246741534e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.462754456201644+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 3.29223551321994e-08 wvoff = 3.72344717737302e-07 pvoff = -1.13573388609373e-13
+ nfactor = {-0.264213898928766+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 5.10682239073404e-07 wnfactor = 2.21827523961945e-06 pnfactor = -3.11253391923814e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 1.35199145537817 leta0 = -4.34213541792014e-07 weta0 = -1.11234153014486e-06 peta0 = 5.6032313600446e-13
+ etab = -0.00399450710172071 letab = 1.01134587900693e-09 wetab = 5.22024606345467e-09 petab = -1.3421836390048e-15
+ dsub = 0.30986317483247 ldsub = -5.71666920670837e-08 wdsub = -3.97019677450401e-07 pdsub = 2.7867285321713e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.340989343402781 lpclm = 4.79873523319717e-07 wpclm = 1.23381685077099e-06 ppclm = -6.12035720647203e-13
+ pdiblc1 = 0.465694320785025 lpdiblc1 = -8.26869304910286e-08 wpdiblc1 = -8.02548753287416e-07 ppdiblc1 = 3.09109096837512e-13
+ pdiblc2 = 0.00474415708928271 lpdiblc2 = -2.00184787749465e-09 wpdiblc2 = -1.92332710096645e-08 ppdiblc2 = 9.53376493207684e-15
+ pdiblcb = -1.99678501045761 lpdiblcb = 5.59156176927921e-07 wpdiblcb = 2.80639505569392e-06 ppdiblcb = -8.53501051614759e-13
+ drout = 0.902326984994161 ldrout = 4.92011208679362e-08 wdrout = 8.70370175201463e-07 pdrout = -4.38434179464758e-13
+ pscbe1 = 799761097.116879 lpscbe1 = 0.120343266023156 wpscbe1 = 0.401460097467861 ppscbe1 = -2.02228699278193e-7
+ pscbe2 = 9.4055268074146e-09 lpscbe2 = -3.1283061207172e-17 wpscbe2 = 2.67224900248169e-17 ppscbe2 = -3.05395468384256e-23
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 13.4631732957545 lbeta0 = -1.46318322701028e-06 wbeta0 = -6.0604748339797e-06 pbeta0 = 2.06051458456296e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.15926055450049e-08 lagidl = 5.65944093810431e-15 wagidl = 1.5812300886917e-14 pagidl = -7.48677326181034e-21
+ bgidl = 1931421692.05947 lbgidl = -469.187843206192 wbgidl = -1565.19100311522 pbgidl = 0.000788438359572237
+ cgidl = 1346.14900055391 lcgidl = -0.000526979774496022 wcgidl = -0.00134998435631258 pcgidl = 6.80031669758406e-10
+ egidl = -5.43588035374289 legidl = 2.78860561823196e-06 wegidl = 7.14367826381721e-06 pegidl = -3.59850648286743e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.408062249251635 lkt1 = -5.05736601777259e-08 wkt1 = -1.2482847000293e-07 pkt1 = 6.28802196799858e-14
+ kt2 = 0.0958453785321361 lkt2 = -7.60804968681285e-08 wkt2 = -2.44137851232674e-07 pkt2 = 1.22980292214988e-13
+ at = 185765.267952839 lat = -0.0415595438442128 wat = -0.157877285060669 pat = 5.46563283809714e-8
+ ute = -0.463595720839178 lute = -5.48121542163133e-08 wute = 2.15217101982415e-07 pute = 1.07254551922507e-13
+ ua1 = 1.58947011996406e-09 lua1 = -5.20487220009854e-16 wua1 = -1.13209038730957e-15 pua1 = 5.70271287070612e-22
+ ub1 = -2.96505896489419e-19 lub1 = 1.36003027665898e-25 wub1 = 1.24166147098232e-24 pub1 = -2.49729986387285e-31
+ uc1 = 4.82993311071544e-11 luc1 = -1.20791803966002e-17 wuc1 = 1.58631477928674e-19 puc1 = -7.99079102714413e-26
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.61 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.856218409482713+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -5.57556095472118e-08 wvth0 = 6.07025902424543e-08 pvth0 = 2.18812258992994e-14
+ k1 = 3.14533704828126 lk1 = -4.42558264468334e-07 wk1 = -5.1675691155279e-06 pk1 = 1.04239860600356e-12
+ k2 = -0.947268468808864 lk2 = 1.63064917644313e-07 wk2 = 1.8644285219467e-06 pk2 = -3.78876718443281e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 51264.0648297486 lvsat = 0.0130860238547209 wvsat = 0.372810919969754 pvsat = -7.95837108821321e-8
+ ua = -6.81973044036041e-09 lua = 9.07778692008775e-16 wua = 9.3986488679654e-15 pua = -1.83821071934767e-21
+ ub = 4.88874324679449e-18 lub = -6.54222119294554e-25 wub = -6.35689421497917e-24 pub = 1.38139745123688e-30
+ uc = -1.02009959094472e-10 luc = 1.88030661365914e-17 wuc = 1.31120109012764e-16 puc = -2.41147960176034e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.00972879047338698 lu0 = 2.58870191220397e-09 wu0 = 2.75182280809925e-08 pu0 = -5.33236847097481e-15
+ a0 = -2.5518117911484 la0 = 5.13307713015792e-07 wa0 = 3.40984101346556e-06 pa0 = -4.26145113638737e-13
+ keta = -1.119048423742 lketa = 2.08034224574093e-07 wketa = 1.30555612779404e-06 pketa = -2.36576357270992e-13
+ a1 = 0.0
+ a2 = 4.57933269347308 la2 = -7.26992765702212e-07 wa2 = -5.78579610168698e-06 pa2 = 1.07827341095382e-12
+ ags = 5.78846997514865 lags = -8.33866703943988e-07 wags = -9.73047940423934e-06 pags = 1.78781017237911e-12
+ b0 = 0.0
+ b1 = 1.83018425978837e-23 lb1 = -4.64378142788883e-30 wb1 = -3.07550056208155e-29 pb1 = 7.80355984118637e-36
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.186871258147022+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -3.70783163597937e-08 wvoff = 5.15955151292737e-08 pvoff = -3.21887311840299e-14
+ nfactor = {3.12524512136215+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -3.49335366522072e-07 wnfactor = -3.43859998504718e-06 pnfactor = 1.12408252945652e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -1.52518770339428 leta0 = 2.95821757700797e-07 weta0 = 3.54420452680811e-06 peta0 = -6.21196264664387e-13
+ etab = 0.612070259368403 letab = -1.55304615511757e-07 wetab = -6.83249285014964e-07 petab = 1.73345255890116e-13
+ dsub = -0.4259168102941 ldsub = 1.29524970899036e-07 wdsub = 2.5743175281882e-06 pdsub = -4.7525344998117e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.88670821701493 lpclm = -5.92832861777749e-07 wpclm = -4.14220489244094e-06 ppclm = 7.52038404323189e-13
+ pdiblc1 = -0.215798692771996 lpdiblc1 = 9.02303363178349e-08 wpdiblc1 = 1.92359168937378e-06 ppdiblc1 = -3.8260269610024e-13
+ pdiblc2 = -0.0368377928346984 lpdiblc2 = 8.54886502256684e-09 wpdiblc2 = 9.14639665350227e-08 ppdiblc2 = -1.85537772418493e-14
+ pdiblcb = 0.100912569201927 lpdiblcb = 2.69010769481674e-08 wpdiblcb = -9.28628743831323e-07 ppdiblcb = 9.41977421101783e-14
+ drout = 1.34883219644943 ldrout = -6.40919859502426e-08 wdrout = -3.1084649114338e-06 pdrout = 5.71127583572466e-13
+ pscbe1 = 800853224.582573 lpscbe1 = -0.156765512230322 wpscbe1 = -1.43378606238912 ppscbe1 = 2.63433814600908e-7
+ pscbe2 = 8.00152215600707e-09 lpscbe2 = 3.24959251008408e-16 wpscbe2 = 9.53880203371062e-16 ppscbe2 = -2.65790054918909e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.21472771990992 lbeta0 = 1.22253614285507e-07 wbeta0 = 4.37829645467242e-06 pbeta0 = -5.8814617082062e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.62866301858439e-08 lagidl = -6.48910118159115e-15 wagidl = -4.66963928013049e-14 pagidl = 8.37374511378328e-21
+ bgidl = -2300856361.30515 lbgidl = 604.680764108172 wbgidl = 5546.86531711201 pbgidl = -0.00101612502672798
+ cgidl = -3436.24643054968 lcgidl = 0.000686471765424184 wcgidl = 0.00482137270111637 pcgidl = -8.85845270494214e-10
+ egidl = 19.8710012633675 legidl = -3.63258537512229e-06 wegidl = -2.551313665649e-05 pegidl = 4.68760513730689e-12
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.980089335993471 lkt1 = 9.45684886225404e-08 wkt1 = 1.03075205502462e-06 pkt1 = -2.30328693676829e-13
+ kt2 = -0.402310435736784 lkt2 = 5.03180723537673e-08 wkt2 = 8.43316238132111e-07 pkt2 = -1.52942696241807e-13
+ at = -179334.971063617 lat = 0.0510784351021497 wat = 0.342410597997361 pat = -7.22832170509918e-8
+ ute = -0.947892086269828 lute = 6.80698154735016e-08 wute = 1.088738723893e-06 pute = -1.1438670976973e-13
+ ua1 = -1.8895187615488e-09 lua1 = 3.62247065863048e-16 wua1 = 3.81142383888943e-15 pua1 = -6.84061408085539e-22
+ ub1 = 2.39502536256411e-19 wub1 = 2.57437951033061e-25
+ uc1 = 3.89823761132943e-12 luc1 = -8.13157740624048e-19 wuc1 = -5.54170849083906e-18 puc1 = 1.3664564510239e-24
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.62 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.56567624281669+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 7.45952065447403e-08 wvth0 = 1.10367903635643e-06 pvth0 = -1.69747965474557e-13
+ k1 = -2.45493284911526 lk1 = 5.86396124590019e-07 wk1 = 3.39047404357496e-06 pk1 = -5.29996337747888e-13
+ k2 = 1.33410837317936 lk2 = -2.5609929366471e-07 wk2 = -1.52653516555132e-06 pk2 = 2.44155212751793e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 803847.932513579 lvsat = -0.125188467906432 wvsat = -0.911983532923894 pvsat = 1.56475428331376e-7
+ ua = 2.66977959082302e-09 lua = -8.35757454550653e-16 wua = -5.79779671551387e-15 pua = 9.53877817041721e-22
+ ub = -3.64192025150027e-18 lub = 9.13142277237636e-25 wub = 6.57406601473101e-24 pub = -9.94446664648461e-31
+ uc = 2.72879257770752e-12 luc = -4.40898924393286e-19 wuc = -2.77727559617639e-18 puc = 4.86572148751079e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0178518903487222 lu0 = -2.47877931728462e-09 wu0 = -1.85603145617363e-08 pu0 = 3.13378040440169e-15
+ a0 = -0.900936199117321 la0 = 2.09987387865146e-07 wa0 = 3.71689911437433e-06 pa0 = -4.82561819693009e-13
+ keta = -0.880788130246744 lketa = 1.64257946069329e-07 wketa = 1.48628237026936e-06 pketa = -2.69781731979709e-13
+ a1 = 0.0
+ a2 = -3.44275966782512 la2 = 7.46930330116191e-07 wa2 = 4.09311845252556e-06 pa2 = -7.3680919683531e-13
+ ags = 1.25
+ b0 = 0.0
+ b1 = -4.27042993950619e-23 lb1 = 6.56506005890105e-30 wb1 = 7.17616797819026e-29 pb1 = -1.10321383179112e-35
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.084715375680311+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -8.69777433527911e-08 wvoff = -9.35384706361355e-07 pvoff = 1.49152105851108e-13
+ nfactor = {-13.3318234189756+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 2.67437120759981e-06 wnfactor = 1.75895494392235e-05 pnfactor = -2.739482448713e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -2.55504315318391 leta0 = 4.85040189056996e-07 weta0 = 3.57464575985378e-06 peta0 = -6.26789323735567e-13
+ etab = -0.897692107971719 letab = 1.22088553526746e-07 wetab = 1.00642429086395e-06 petab = -1.37103539226845e-13
+ dsub = 0.376647253109009 ldsub = -1.79325321622072e-08 wdsub = -7.55455858188785e-08 pdsub = 1.16138495446936e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.89438342328049 lpclm = -5.9424305045054e-07 wpclm = -4.18464086246844e-06 ppclm = 7.59835292404252e-13
+ pdiblc1 = 3.66574502734349 lpdiblc1 = -6.22937336010143e-07 wpdiblc1 = -4.46720531730067e-06 ppdiblc1 = 7.91597610327076e-13
+ pdiblc2 = 0.0948050946725187 lpdiblc2 = -1.56382776277967e-08 wpdiblc2 = -1.21574378438021e-07 ppdiblc2 = 2.0588396995083e-14
+ pdiblcb = -1.06009642187104 lpdiblcb = 2.40216741904977e-07 wpdiblcb = 1.77963790169567e-06 ppdiblcb = -4.03400213472433e-13
+ drout = 1.0
+ pscbe1 = 800000000.0
+ pscbe2 = 9.6239320007883e-09 lpscbe2 = 2.68690229972105e-17 wpscbe2 = 1.08158518454985e-15 ppscbe2 = -2.89253674225825e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 16.4248694146139 lbeta0 = -1.56995334970753e-06 wbeta0 = -4.20036095178245e-06 pbeta0 = 9.88036290439571e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.49817556120657e-09 lagidl = -1.01597904804267e-15 wagidl = -1.02454537108168e-14 pagidl = 1.67650472187062e-21
+ bgidl = 940150742.549778 lbgidl = 9.20080589559575 wbgidl = 100.572619365448 pbgidl = -1.54613304929087e-5
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = 0.786908957748391 lkt1 = -2.30087408881534e-07 wkt1 = -1.36485087836635e-06 pkt1 = 2.09822620083894e-13
+ kt2 = -0.171722364515308 lkt2 = 7.95143426403179e-09 wkt2 = 6.67442046306901e-08 pkt2 = -1.02607868104899e-14
+ at = 601953.792063103 lat = -0.0924700932134119 wat = -0.646221591689261 pat = 1.093611410567e-7
+ ute = -2.44772466743709 lute = 3.43638555109106e-07 wute = 2.85501740624339e-06 pute = -4.38910390914014e-13
+ ua1 = -3.11875789184375e-11 lua1 = 2.0810302684823e-17 wua1 = 1.93432723101731e-17 pua1 = 1.26689306537679e-23
+ ub1 = -4.23637384533365e-19 lub1 = 1.21840687066468e-25 wub1 = 1.57666156857191e-24 pub1 = -2.42384912921265e-31
+ uc1 = -3.62751575593886e-11 luc1 = 6.56802067427748e-18 wuc1 = 1.16087241625521e-17 puc1 = -1.78464399168162e-24
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.63 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1e-06 wmax = 1.26e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.009332+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.49177002
+ k2 = -0.002490247
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 55237.817
+ ua = -1.4022531e-9
+ ub = 1.481232e-18
+ uc = -3.8916596e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0070157252
+ a0 = 1.216808
+ keta = 0.0066402373
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.28483517
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.28448891+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.6339038+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0017402344
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00056783834
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 799985290.0
+ pscbe2 = 1.0771971e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.4670794e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.54561
+ kt2 = -0.052484
+ at = 10000.0
+ ute = -1.2595
+ ua1 = -2.5605e-10
+ ub1 = 4.9434e-19
+ uc1 = 8.1951e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.64 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1e-06 wmax = 1.26e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.009332+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.49177002
+ k2 = -0.002490247
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 55237.817
+ ua = -1.4022531e-9
+ ub = 1.481232e-18
+ uc = -3.8916596e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0070157252
+ a0 = 1.216808
+ keta = 0.0066402373
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.28483517
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.28448891+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.6339038+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0017402344
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00056783834
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 799985290.0
+ pscbe2 = 1.0771971e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.4670794e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.54561
+ kt2 = -0.052484
+ at = 10000.0
+ ute = -1.2595
+ ua1 = -2.5605e-10
+ ub1 = 4.9434e-19
+ uc1 = 8.1951e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.65 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1e-06 wmax = 1.26e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.00965248881732+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.56510692328967e-9
+ k1 = 0.533820717223042 lk1 = -3.36562553037073e-7
+ k2 = -0.015002741397731 lk2 = 1.00146664323435e-07 wk2 = 3.30872245021211e-24 pk2 = 1.26217744835362e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 67741.5222028627 lvsat = -0.100076317954424
+ ua = -1.97423156119557e-09 lua = 4.5779628851602e-15
+ ub = 1.81069574535962e-18 lub = -2.63693985103838e-24
+ uc = -2.32479618811687e-11 luc = -1.25407563961816e-16
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00451481860506789 lu0 = 2.00165886437757e-8
+ a0 = 1.29911774394725 la0 = -6.58785213852157e-7
+ keta = 0.0100612720038462 lketa = -2.73810483533195e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.225999022361107 lags = 4.70908816450275e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.302660162509807+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.4543785336408e-7
+ nfactor = {1.25753668288135+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.01234191539741e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.0345570080176767 lpclm = 2.90513436947359e-07 wpclm = 6.61744490042422e-24 ppclm = 3.78653234506086e-29
+ pdiblc1 = 0.39
+ pdiblc2 = 9.73517077413289e-05 lpdiblc2 = 3.76564938466757e-9
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 799970586.290556 lpscbe1 = 0.117684564487718
+ pscbe2 = 1.20422461789891e-08 lpscbe2 = -1.01669433691559e-14
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.35927238290888e-10 lagidl = 8.62858580323798e-17
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.630018700972499 lkt1 = 6.75584705460732e-7
+ kt2 = -0.0782500237215 lkt2 = 2.06224374338552e-7
+ at = -35310.746827625 lat = 0.362655119638908 pat = -1.05879118406788e-22
+ ute = -2.450110100875 lute = 9.52932535450658e-6
+ ua1 = -2.4337304253625e-09 lua1 = 1.74295726839279e-14 wua1 = 3.94430452610506e-31 pua1 = 4.51389830715758e-36
+ ub1 = 2.00558905818e-18 lub1 = -1.20956339581742e-23
+ uc1 = 9.6472508077075e-11 luc1 = -7.06548804180952e-16 wuc1 = -4.93038065763132e-32 puc1 = 2.35098870164458e-37
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.66 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1e-06 wmax = 1.26e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.01358213461837+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.82983594952644e-8
+ k1 = 0.438259517078265 lk1 = 4.6038977502179e-8
+ k2 = 0.01323300444793 lk2 = -1.29017230984511e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 32034.083885955 lvsat = 0.0428867311804437
+ ua = -6.34366705527208e-10 lua = -7.86498253019447e-16
+ ub = 9.9159484100627e-19 lub = 6.42521470050967e-25
+ uc = -6.41266971865545e-11 luc = 3.82599775786224e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0101366594698 lu0 = -2.49176114710077e-9
+ a0 = 1.188040607639 la0 = -2.14062017669315e-7
+ keta = 0.0112740092448839 lketa = -3.22365244655909e-08 wketa = 6.61744490042422e-24 pketa = 1.26217744835362e-29
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.263068487300985 lags = 3.22492576378146e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.264697760530965+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -6.55346819787902e-9
+ nfactor = {2.3242968912748+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.25868113403433e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.15964838675 leta0 = -3.18890874427738e-7
+ etab = -0.139629720257219 letab = 2.78778808774596e-7
+ dsub = 0.86055995 ldsub = -1.20336179029335e-6
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.276866772705234 lpclm = 1.26065703804917e-06 wpclm = -5.29395592033938e-23
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00186230851727895 lpdiblc2 = -3.3007664372529e-9
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 799999959.962669 lpscbe1 = 8.02241193014197e-5
+ pscbe2 = 9.63387073834225e-09 lpscbe2 = -5.24451141048652e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.0546779342355e-12 lalpha0 = 1.22301148496705e-17
+ alpha1 = 2.92931788562325e-15 lalpha1 = -1.172820668616e-20
+ beta0 = 57.0503955 lbeta0 = -0.000108302561126402 pbeta0 = 1.03397576569128e-25
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.6405047926645e-11 lagidl = 3.64634145825979e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.451571913615 lkt1 = -3.88685858264734e-8
+ kt2 = -0.00791993406450003 lkt2 = -7.53585265141372e-8
+ at = 103166.7354985 lat = -0.191771746107116
+ ute = 0.756589955825 lute = -3.30944548360509e-06 pute = -2.01948391736579e-28
+ ua1 = 3.996379086515e-09 lua1 = -8.31486896238996e-15
+ ub1 = -2.780979127635e-18 lub1 = 7.06850704412346e-24
+ uc1 = -2.22130792889e-10 luc1 = 5.69053745805855e-16 wuc1 = -9.86076131526265e-32 puc1 = -1.88079096131566e-37
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.67 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1e-06 wmax = 1.26e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0135817620874+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.82976130426718e-8
+ k1 = 0.46889012614082 lk1 = -1.53365846865645e-8
+ k2 = 0.004468587922708 lk2 = 4.65982751888154e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 78156.2910646471 lvsat = -0.0495298573763384
+ ua = -1.28367292089777e-09 lua = 5.14538037823651e-16
+ ub = 1.52974540449884e-18 lub = -4.35788572987695e-25
+ uc = -4.13713352669989e-11 luc = -7.33569202653429e-18
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00846149481000001 lu0 = 8.64821562174285e-10
+ a0 = 1.664236346647 la0 = -1.16823113437903e-6
+ keta = 0.0283355753681761 lketa = -6.64233475385135e-08 wketa = -1.32348898008484e-23 pketa = 1.89326617253043e-29
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.452034387421789 lags = 1.75536780485503e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.2627688523134+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.04184852473844e-8
+ nfactor = {1.6824868640504+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.73347972461008e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.0792967735 leta0 = 1.59891428355475e-07 weta0 = -2.56425989891439e-23 peta0 = -7.88860905221012e-30
+ etab = 0.00602426151443782 letab = -1.30728810826712e-08 wetab = -2.48154183765908e-24 petab = -3.15544362088405e-30
+ dsub = -0.0411199 ldsub = 6.033638805867e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.33312711053902 lpclm = 3.83921643945076e-8
+ pdiblc1 = 0.397789640581111 lpdiblc1 = -1.56083598905101e-8
+ pdiblc2 = 0.000215
+ pdiblcb = -0.4257466 lpdiblcb = 4.022425870578e-7
+ drout = 0.2074359732976 ldrout = 7.0644417491648e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0338000872575e-08 lpscbe2 = -1.93533992730523e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -9.4263944131529e-11 lalpha0 = 1.94989131434972e-16 walpha0 = 3.08148791101958e-32 palpha0 = 1.76324152623343e-38
+ alpha1 = -1.00379158635771e-10 lalpha1 = 2.01127174034959e-16 walpha1 = 1.08514115304068e-32 palpha1 = -3.1729163922586e-38
+ beta0 = -2.92305473080459 lbeta0 = 1.18682202249193e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.9731883172318e-10 lagidl = -2.98428722922003e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.42793321116691 lkt1 = -8.62342339988934e-8
+ kt2 = -0.0271141028514701 lkt2 = -3.68985371081153e-8
+ at = -8088.88726421299 lat = 0.0311548166580833 pat = -1.32348898008484e-23
+ ute = -0.595554641860501 lute = -6.00108732450936e-7
+ ua1 = -6.58322299788103e-11 lua1 = -1.75282094557869e-16
+ ub1 = 1.01445607323126e-18 lub1 = -5.36531717213893e-25
+ uc1 = 7.63492890397921e-11 luc1 = -2.90206441975695e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.68 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 1e-06 wmax = 1.26e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0292173636172+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.39915822729837e-8
+ k1 = 0.39769231810658 lk1 = 5.61270047650684e-8
+ k2 = 0.0233960636905084 lk2 = -1.43383045159601e-08 wk2 = 1.32348898008484e-23
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -31885.517316294 lvsat = 0.0609227370752887 pvsat = -2.64697796016969e-23
+ ua = -4.04712121209061e-10 lua = -3.67703922530296e-16
+ ub = 8.65580930285482e-19 lub = 2.30855227207905e-25
+ uc = -7.5763218738422e-11 luc = 2.71845763458875e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0113181849198 lu0 = -2.00253257180562e-9
+ a0 = -0.1393405367 la0 = 6.42078501473501e-7
+ keta = -0.042358236715718 lketa = 4.53436454588974e-9
+ a1 = 0.0
+ a2 = 0.8
+ ags = 1.2808267907332 lags = 1.6037855921993e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.26264494090254+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.05428592195409e-8
+ nfactor = {1.427577131768+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.8319610755911e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.33306106 leta0 = 4.1460301693698e-07 peta0 = 5.04870979341448e-29
+ etab = -0.0140459653375 letab = 7.07226792610489e-9
+ dsub = 0.80439263362832 ldsub = -2.45304951329654e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.11462330639098 lpclm = 2.57711643243433e-7
+ pdiblc1 = 0.61102244661888 lpdiblc1 = -2.29637163993218e-7
+ pdiblc2 = -0.000104560407338499 lpdiblc2 = 3.20753326339095e-10
+ pdiblcb = -0.025
+ drout = 0.8218430134048 ldrout = 8.97435533285599e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 7.49579255568821e-09 lpscbe2 = 9.17478353228516e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.76919111342539 lbeta0 = 1.32327226952781e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.804433234633e-10 lagidl = 2.81490218389788e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.51927367732618 lkt1 = 5.44720612054921e-9
+ kt2 = -0.0726276802030601 lkt2 = 8.78494242772801e-9
+ at = -19413.822844574 lat = 0.0425220282229658
+ ute = -2.153346615999 lute = 9.63498479127023e-7
+ ua1 = -1.04308281636238e-09 lua1 = 8.05616568264671e-16 wua1 = 3.94430452610506e-31
+ ub1 = 4.0779506741748e-19 lub1 = 7.23939541345907e-26
+ uc1 = 7.07257403564161e-11 luc1 = -2.33761028069585e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.69 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 1e-06 wmax = 1.26e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.961379729003999+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.80472923627924e-10
+ k1 = 0.436921098622959 lk1 = 3.63661734692107e-8
+ k2 = 0.00697647073255922 lk2 = -6.06721369647345e-09 pk2 = -1.57772181044202e-30
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 28540.8777037199 lvsat = 0.030483967832672
+ ua = -6.89954909723199e-10 lua = -2.24017716943703e-16
+ ub = 1.0404179671488e-18 lub = 1.42784042117633e-25
+ uc = -4.39756885037937e-11 luc = 1.11721483782075e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00920019660524 lu0 = -9.3563196414736e-10
+ a0 = 1.46331587308 la0 = -1.65232419794208e-7
+ keta = -0.0570929960904168 lketa = 1.1956749089985e-8
+ a1 = 0.0
+ a2 = 1.08040210428168 la2 = -1.41247793196124e-7
+ ags = 2.21682838003568 lags = -4.55457032662113e-07 pags = -4.03896783473158e-28
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.17421181309548+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -5.50895439891745e-8
+ nfactor = {1.454803372664+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 2.69481351553846e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = 5.08399250000001e-05 letab = -2.8758079190025e-11 wetab = 2.58493941422821e-26 petab = 9.24446373305873e-33
+ dsub = 0.00219906241307921 ldsub = 1.58786422879312e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.61513748818976 lpclm = 5.58613290338762e-9
+ pdiblc1 = -0.156228127591121 lpdiblc1 = 1.56852269505308e-07 ppdiblc1 = -5.04870979341448e-29
+ pdiblc2 = -0.010160361729811 lpdiblc2 = 5.38619229391214e-09 wpdiblc2 = 8.27180612553028e-25 ppdiblc2 = -5.91645678915759e-31
+ pdiblcb = 0.1779864 lpdiblcb = -1.022509482312e-07 ppdiblcb = 2.52435489670724e-29
+ drout = 1.57680657036212 ldrout = -2.90556504108222e-7
+ pscbe1 = 800072202.262479 lpscbe1 = -0.0363706622856625
+ pscbe2 = 9.42623497792119e-09 lpscbe2 = -5.49491994501789e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.76670428794479 lbeta0 = 1.33579923012603e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.608866469266e-10 lagidl = -1.42315451584627e-16
+ bgidl = 718501708.2624 lbgidl = 141.799978991857
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.50479609548 lkt1 = -1.84562961557289e-9
+ kt2 = -0.0933453834719999 lkt2 = 1.9221133248501e-8
+ at = 63420.7658079999 lat = 0.000795512377238711
+ ute = -0.29681663552 lute = 2.83030624703961e-8
+ ua1 = 7.12174600439999e-10 lua1 = -7.85645160734427e-17 wua1 = 7.88860905221012e-31
+ ub1 = 6.6569999932e-19 lub1 = -5.75212709274614e-26 wub1 = 7.3468396926393e-40
+ uc1 = 4.842226005912e-11 luc1 = -1.21411037663607e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.70 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1e-06 wmax = 1.26e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.809177898371427+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -3.8799100015522e-8
+ k1 = -0.859188811758427 lk1 = 3.65232029360011e-7
+ k2 = 0.497540891920585 lk2 = -1.30539595977775e-07 wk2 = 5.29395592033938e-23 pk2 = -1.26217744835362e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 340167.983973857 lvsat = -0.0485861127225686
+ ua = 4.6360367666286e-10 lua = -5.16713597743197e-16
+ ub = -3.74312666585699e-20 lub = 4.16269961759279e-25
+ uc = -4.00506840596299e-13 luc = 1.1568680925945e-19
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0115960246397143 lu0 = -1.54353259881863e-9
+ a0 = 0.0905905090000019 la0 = 1.83073305009902e-7
+ keta = -0.107328375378326 lketa = 2.47031225828439e-08 wketa = 2.64697796016969e-23 pketa = -1.26217744835362e-29
+ a1 = 0.0
+ a2 = 0.0957216198444293 la2 = 1.08598140161594e-7
+ ags = -1.75201096157886 lags = 5.51568480003769e-07 pags = 2.01948391736579e-28
+ b0 = 0.0
+ b1 = -5.53126201684571e-24 lb1 = 1.40346370532031e-30
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.146888130688428+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -6.20224638973629e-8
+ nfactor = {0.460556511571433+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 5.21754590359447e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 1.22133747383557 leta0 = -1.85564451248721e-07 peta0 = -2.01948391736579e-28
+ etab = 0.0825970448787428 letab = -2.0973454300718e-08 wetab = 9.51257704435982e-24 petab = -5.47272252997077e-30
+ dsub = 1.569009795062 ldsub = -2.38765164747896e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.676772125493857 lpclm = -1.00526085236927e-8
+ pdiblc1 = 1.274858227734 lpdiblc1 = -2.06261564690401e-7
+ pdiblc2 = 0.03404075974251 lpdiblc2 = -5.82909086062429e-9
+ pdiblcb = -0.618713571428571 lpdiblcb = 9.98981256192858e-8
+ drout = -1.060023465579 ldrout = 3.78494291401226e-7
+ pscbe1 = 799742134.776857 lpscbe1 = 0.0473783510442445
+ pscbe2 = 8.74071651536284e-09 lpscbe2 = 1.18989456610138e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 10.6076192291828 lbeta0 = -3.33520947772555e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1997599084.17429 lbgidl = -182.749235490394
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.18132435242857 lkt1 = -8.39210853952409e-8
+ kt2 = 0.251204129485714 lkt2 = -6.82024483227987e-08 wkt2 = -1.05879118406788e-22 pkt2 = -1.26217744835362e-29
+ at = 86010.699942857 lat = -0.00493629938060097
+ ute = -0.104191251857143 lute = -2.05723540025315e-8
+ ua1 = 1.06408379028571e-09 lua1 = -1.67855490540565e-16 pua1 = -1.88079096131566e-37
+ ub1 = 4.39e-19
+ uc1 = -3.96221633285712e-13 luc1 = 2.45756048898484e-19
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.71 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1e-06 wmax = 1.26e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.45474596731129+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.03919942004995e-07 wvth0 = -3.29901163110622e-07 pvth0 = 6.06137304018042e-14
+ k1 = 3.87262543122222 lk1 = -5.04158396945551e-07 wk1 = -4.77481090874912e-06 pk1 = 8.77290332697203e-13
+ k2 = -1.23821757446287 lk2 = 1.88376514326255e-07 wk2 = 1.79287706618172e-06 pk2 = -3.29410682000765e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -444299.081126228 lvsat = 0.0955463745494654 wvsat = 0.698665563810752 pvsat = -1.28367920035641e-7
+ ua = -1.40856932079402e-08 lua = 2.15647236675556e-15 wua = 1.58240049102342e-14 pua = -2.90739189417207e-21
+ ub = 1.34999204020476e-17 lub = -2.07098827238711e-24 wub = -1.55463171318762e-23 pub = 2.85637148559101e-30
+ uc = 2.0129128432757e-12 luc = -3.27738029517404e-19 wuc = -1.85348133553812e-18 puc = 3.40545686222426e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.0237963794061442 lu0 = 4.9592199737391e-09 wu0 = 3.51839538042294e-08 pu0 = -6.46445338431249e-15
+ a0 = -1.81630643727311 la0 = 5.33433201639502e-07 wa0 = 4.89812234461224e-06 pa0 = -8.9994671274264e-13
+ keta = 0.678955884962581 lketa = -1.19763243422372e-07 wketa = -5.26461530714046e-07 pketa = 9.67283564226838e-14
+ a1 = 0.0
+ a2 = 2.28472879813727 la2 = -2.93594715727683e-07 wa2 = -3.2978170890809e-06 pa2 = 6.05917827228101e-13
+ ags = 1.25
+ b0 = -1.01482832252494e-08 lb0 = 1.86457452182475e-15 wb0 = 1.30956714485817e-14 pb0 = -2.40610700226226e-21
+ b1 = 1.67516028991626e-09 lb1 = -3.07782225547183e-16 wb1 = -2.16168077826925e-15 pb1 = 3.97172094433745e-22
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.602175173640312+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 2.16287903653147e-08 wvoff = -4.89990236423409e-08 pvoff = 9.00273761087818e-15
+ nfactor = {-2.12235874457582+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 9.96321359117152e-07 wnfactor = 3.12449527861546e-06 pnfactor = -5.74072891025853e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 2.88894120920656 leta0 = -4.9195828835964e-07 weta0 = -3.45044695767136e-06 peta0 = 6.33960970873832e-13
+ etab = 0.181345053091477 letab = -3.91167220936683e-08 wetab = -3.86000006768583e-07 petab = 7.09209392436121e-14
+ dsub = 0.445819350865307 ldsub = -3.23980148643053e-08 wdsub = -1.64807488105155e-07 pdsub = 3.02805742120241e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.64983316297734 lpclm = 6.01154560942986e-07 wpclm = 4.26022694421274e-06 ppclm = -7.82744277141039e-13
+ pdiblc1 = -2.28698517554903 lpdiblc1 = 4.48166609325e-07 wpdiblc1 = 3.21438941442436e-06 ppdiblc1 = -5.90589410280431e-13
+ pdiblc2 = -0.0445117312871088 lpdiblc2 = 8.60359397372065e-09 wpdiblc2 = 5.82045397820781e-08 ppdiblc2 = -1.06940947077805e-14
+ pdiblcb = 3.4032208721455 lpdiblcb = -6.39063955501908e-07 wpdiblcb = -3.97997045332014e-06 ppdiblcb = 7.31251911299869e-13
+ drout = 1.0
+ pscbe1 = 800000000.0
+ pscbe2 = 1.44697279813175e-08 lpscbe2 = -9.33619007064111e-16 wpscbe2 = -5.17158598335559e-15 ppscbe2 = 9.50191007479866e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -0.780508729123767 lbeta0 = 1.758853966391e-06 wbeta0 = 1.80020130180728e-05 pbeta0 = -3.30756385784956e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.10115738502735e-09 lagidl = -1.65380964982323e-15 wagidl = -1.36044252722899e-14 pagidl = 2.49958186855363e-21
+ bgidl = 1018087901.40667 lbgidl = -2.78070734695029
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.270760618666667 lkt1 = -6.7488691890517e-8
+ kt2 = -0.12
+ at = -504708.512248689 lat = 0.103598313632988 wat = 0.781851080320874 pat = -1.43651844540595e-7
+ ute = -0.235274136333333 lute = 3.51189761093216e-9
+ ua1 = -1.54771143080642e-09 lua1 = 3.12017480816356e-16 wua1 = 1.97631448285446e-15 pua1 = -3.63114188878299e-22
+ ub1 = 7.98171532333336e-19 lub1 = -6.59916631502001e-26
+ uc1 = 3.44047199689403e-12 luc1 = -4.59171181855323e-19 wuc1 = -3.96416030601466e-17 puc1 = 7.28347065504992e-24
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.72 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.009332+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.49177002
+ k2 = -0.002490247
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 55237.817
+ ua = -1.4022531e-9
+ ub = 1.481232e-18
+ uc = -3.8916596e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0070157252
+ a0 = 1.216808
+ keta = 0.0066402373
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.28483517
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.28448891+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.6339038+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0017402344
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00056783834
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 799985290.0
+ pscbe2 = 1.0771971e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.4670794e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.54561
+ kt2 = -0.052484
+ at = 10000.0
+ ute = -1.2595
+ ua1 = -2.5605e-10
+ ub1 = 4.9434e-19
+ uc1 = 8.1951e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.73 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.009332+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.49177002
+ k2 = -0.002490247
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 55237.817
+ ua = -1.4022531e-9
+ ub = 1.481232e-18
+ uc = -3.8916596e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0070157252
+ a0 = 1.216808
+ keta = 0.0066402373
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.28483517
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.28448891+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.6339038+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0017402344
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00056783834
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 799985290.0
+ pscbe2 = 1.0771971e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.4670794e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.54561
+ kt2 = -0.052484
+ at = 10000.0
+ ute = -1.2595
+ ua1 = -2.5605e-10
+ ub1 = 4.9434e-19
+ uc1 = 8.1951e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.74 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.00965248881731+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.56510692328967e-9
+ k1 = 0.533820717223042 lk1 = -3.36562553037073e-7
+ k2 = -0.015002741397731 lk2 = 1.00146664323435e-07 wk2 = 3.30872245021211e-24 pk2 = -2.52435489670724e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 67741.5222028627 lvsat = -0.100076317954424
+ ua = -1.97423156119557e-09 lua = 4.5779628851602e-15
+ ub = 1.81069574535962e-18 lub = -2.6369398510384e-24
+ uc = -2.32479618811687e-11 luc = -1.25407563961816e-16
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00451481860506789 lu0 = 2.00165886437757e-8
+ a0 = 1.29911774394725 la0 = -6.58785213852143e-7
+ keta = 0.0100612720038463 lketa = -2.73810483533195e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.225999022361107 lags = 4.70908816450277e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.302660162509807+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.45437853364081e-7
+ nfactor = {1.25753668288135+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.01234191539741e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.0345570080176767 lpclm = 2.90513436947359e-07 wpclm = -6.61744490042422e-24 ppclm = -5.04870979341448e-29
+ pdiblc1 = 0.39
+ pdiblc2 = 9.73517077413289e-05 lpdiblc2 = 3.76564938466757e-9
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 799970586.290556 lpscbe1 = 0.117684564480442
+ pscbe2 = 1.20422461789891e-08 lpscbe2 = -1.01669433691559e-14
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.35927238290887e-10 lagidl = 8.62858580323798e-17
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.6300187009725 lkt1 = 6.75584705460732e-7
+ kt2 = -0.0782500237214999 lkt2 = 2.06224374338553e-7
+ at = -35310.746827625 lat = 0.362655119638908 wat = 1.38777878078145e-17 pat = 2.11758236813575e-22
+ ute = -2.450110100875 lute = 9.52932535450658e-06 pute = 6.46234853557053e-27
+ ua1 = -2.4337304253625e-09 lua1 = 1.74295726839279e-14
+ ub1 = 2.00558905818e-18 lub1 = -1.20956339581742e-23
+ uc1 = 9.64725080770751e-11 luc1 = -7.06548804180952e-16 wuc1 = -4.93038065763132e-32 puc1 = -3.76158192263132e-37
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.75 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.01358213461837+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.8298359495261e-8
+ k1 = 0.438259517078265 lk1 = 4.60389775021774e-8
+ k2 = 0.01323300444793 lk2 = -1.29017230984511e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 32034.083885955 lvsat = 0.0428867311804439
+ ua = -6.3436670552721e-10 lua = -7.86498253019447e-16
+ ub = 9.9159484100627e-19 lub = 6.42521470050961e-25
+ uc = -6.41266971865545e-11 luc = 3.82599775786226e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0101366594698 lu0 = -2.49176114710077e-9
+ a0 = 1.188040607639 la0 = -2.14062017669312e-7
+ keta = 0.0112740092448839 lketa = -3.22365244655909e-08 pketa = 1.26217744835362e-29
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.263068487300985 lags = 3.22492576378147e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.264697760530965+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -6.55346819787817e-9
+ nfactor = {2.3242968912748+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.25868113403433e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.15964838675 leta0 = -3.18890874427738e-7
+ etab = -0.139629720257219 letab = 2.78778808774596e-7
+ dsub = 0.86055995 ldsub = -1.20336179029335e-06 wdsub = -8.470329472543e-22
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.276866772705234 lpclm = 1.26065703804917e-06 ppclm = 2.01948391736579e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00186230851727895 lpdiblc2 = -3.3007664372529e-9
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 799999959.962669 lpscbe1 = 8.02241193014197e-5
+ pscbe2 = 9.63387073834223e-09 lpscbe2 = -5.24451141048627e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.0546779342355e-12 lalpha0 = 1.22301148496705e-17
+ alpha1 = 2.92931788562325e-15 lalpha1 = -1.172820668616e-20
+ beta0 = 57.0503955 lbeta0 = -0.000108302561126402
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.6405047926645e-11 lagidl = 3.64634145825981e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.451571913615 lkt1 = -3.88685858264768e-8
+ kt2 = -0.00791993406450003 lkt2 = -7.53585265141372e-8
+ at = 103166.7354985 lat = -0.191771746107116
+ ute = 0.756589955824999 lute = -3.30944548360509e-06 wute = -3.17637355220363e-22 pute = -1.21169035041947e-27
+ ua1 = 3.996379086515e-09 lua1 = -8.31486896238996e-15 pua1 = -6.01853107621011e-36
+ ub1 = -2.780979127635e-18 lub1 = 7.06850704412346e-24 wub1 = -1.46936793852786e-39 pub1 = 2.80259692864963e-45
+ uc1 = -2.22130792889e-10 luc1 = 5.69053745805855e-16 wuc1 = -1.97215226305253e-31
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.76 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0135817620874+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.82976130426718e-8
+ k1 = 0.468890126140821 lk1 = -1.53365846865628e-8
+ k2 = 0.004468587922708 lk2 = 4.65982751888153e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 78156.2910646471 lvsat = -0.0495298573763382
+ ua = -1.28367292089777e-09 lua = 5.14538037823651e-16
+ ub = 1.52974540449884e-18 lub = -4.35788572987695e-25
+ uc = -4.13713352669991e-11 luc = -7.33569202653429e-18
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00846149481000001 lu0 = 8.64821562174272e-10
+ a0 = 1.664236346647 la0 = -1.16823113437903e-6
+ keta = 0.0283355753681761 lketa = -6.64233475385135e-08 wketa = -1.32348898008484e-23 pketa = 6.31088724176809e-30
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.452034387421789 lags = 1.75536780485504e-06 pags = 8.07793566946316e-28
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.2627688523134+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.0418485247384e-8
+ nfactor = {1.6824868640504+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.73347972461008e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.0792967735 leta0 = 1.59891428355475e-07 weta0 = 1.48892510259545e-23 peta0 = -9.46633086265214e-30
+ etab = 0.00602426151443783 letab = -1.30728810826712e-08 wetab = 1.65436122510606e-24 petab = -1.57772181044202e-30
+ dsub = -0.0411199 ldsub = 6.03363880586701e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.333127110539021 lpclm = 3.83921643945084e-8
+ pdiblc1 = 0.39778964058111 lpdiblc1 = -1.56083598905093e-8
+ pdiblc2 = 0.000215
+ pdiblcb = -0.4257466 lpdiblcb = 4.022425870578e-7
+ drout = 0.2074359732976 ldrout = 7.0644417491648e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0338000872575e-08 lpscbe2 = -1.93533992730521e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -9.42639441315289e-11 lalpha0 = 1.94989131434972e-16 walpha0 = 2.46519032881566e-32 palpha0 = 8.22846045575601e-38
+ alpha1 = -1.00379158635771e-10 lalpha1 = 2.01127174034959e-16 walpha1 = -4.08658260074667e-32 palpha1 = 6.4187272095926e-38
+ beta0 = -2.92305473080459 lbeta0 = 1.18682202249193e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.9731883172318e-10 lagidl = -2.98428722922003e-16 wagidl = -3.94430452610506e-31
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.427933211166911 lkt1 = -8.62342339988934e-8
+ kt2 = -0.0271141028514701 lkt2 = -3.68985371081154e-8
+ at = -8088.88726421299 lat = 0.0311548166580833
+ ute = -0.595554641860502 lute = -6.00108732450933e-7
+ ua1 = -6.58322299788099e-11 lua1 = -1.75282094557869e-16
+ ub1 = 1.01445607323126e-18 lub1 = -5.36531717213891e-25
+ uc1 = 7.63492890397921e-11 luc1 = -2.90206441975695e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.77 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0292173636172+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.39915822729828e-8
+ k1 = 0.39769231810658 lk1 = 5.6127004765068e-8
+ k2 = 0.0233960636905084 lk2 = -1.43383045159601e-08 wk2 = -1.32348898008484e-23
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -31885.5173162939 lvsat = 0.0609227370752887 pvsat = 2.64697796016969e-23
+ ua = -4.04712121209062e-10 lua = -3.67703922530297e-16
+ ub = 8.6558093028548e-19 lub = 2.30855227207905e-25
+ uc = -7.57632187384221e-11 luc = 2.71845763458875e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0113181849198 lu0 = -2.00253257180561e-9
+ a0 = -0.139340536699999 la0 = 6.42078501473501e-7
+ keta = -0.042358236715718 lketa = 4.53436454588976e-9
+ a1 = 0.0
+ a2 = 0.8
+ ags = 1.2808267907332 lags = 1.6037855921993e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.262644940902541+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.05428592195407e-8
+ nfactor = {1.427577131768+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.8319610755911e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.33306106 leta0 = 4.1460301693698e-07 weta0 = -1.05879118406788e-22 peta0 = 1.51461293802434e-28
+ etab = -0.0140459653375 letab = 7.07226792610489e-9
+ dsub = 0.80439263362832 ldsub = -2.45304951329654e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.11462330639098 lpclm = 2.57711643243433e-7
+ pdiblc1 = 0.61102244661888 lpdiblc1 = -2.29637163993218e-7
+ pdiblc2 = -0.000104560407338499 lpdiblc2 = 3.20753326339095e-10 ppdiblc2 = -1.97215226305253e-31
+ pdiblcb = -0.025
+ drout = 0.8218430134048 ldrout = 8.97435533285599e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 7.49579255568821e-09 lpscbe2 = 9.17478353228516e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.76919111342541 lbeta0 = 1.32327226952781e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.804433234633e-10 lagidl = 2.81490218389789e-16 pagidl = -9.4039548065783e-38
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.51927367732618 lkt1 = 5.44720612054837e-9
+ kt2 = -0.0726276802030601 lkt2 = 8.78494242772796e-9
+ at = -19413.8228445739 lat = 0.0425220282229658
+ ute = -2.153346615999 lute = 9.63498479127025e-7
+ ua1 = -1.04308281636238e-09 lua1 = 8.05616568264671e-16
+ ub1 = 4.0779506741748e-19 lub1 = 7.23939541345903e-26
+ uc1 = 7.07257403564161e-11 luc1 = -2.33761028069585e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.78 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.961379729003999+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.80472923627924e-10
+ k1 = 0.436921098622959 lk1 = 3.63661734692105e-8
+ k2 = 0.00697647073255922 lk2 = -6.06721369647345e-09 pk2 = 3.15544362088405e-30
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 28540.8777037198 lvsat = 0.030483967832672
+ ua = -6.89954909723197e-10 lua = -2.24017716943704e-16
+ ub = 1.0404179671488e-18 lub = 1.42784042117634e-25
+ uc = -4.39756885037937e-11 luc = 1.11721483782075e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00920019660524 lu0 = -9.3563196414736e-10
+ a0 = 1.46331587308 la0 = -1.65232419794208e-7
+ keta = -0.0570929960904167 lketa = 1.19567490899849e-8
+ a1 = 0.0
+ a2 = 1.08040210428168 la2 = -1.41247793196124e-7
+ ags = 2.21682838003568 lags = -4.55457032662114e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.17421181309548+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -5.50895439891748e-8
+ nfactor = {1.454803372664+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 2.69481351553846e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = 5.08399250000001e-05 letab = -2.8758079190025e-11 wetab = 2.58493941422821e-26 petab = 6.16297582203915e-33
+ dsub = 0.0021990624130801 ldsub = 1.58786422879312e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.61513748818976 lpclm = 5.58613290338783e-9
+ pdiblc1 = -0.15622812759112 lpdiblc1 = 1.56852269505308e-7
+ pdiblc2 = -0.010160361729811 lpdiblc2 = 5.38619229391214e-09 wpdiblc2 = 1.65436122510606e-24 ppdiblc2 = 2.36658271566304e-30
+ pdiblcb = 0.1779864 lpdiblcb = -1.022509482312e-07 wpdiblcb = 5.29395592033938e-23 ppdiblcb = 3.78653234506086e-29
+ drout = 1.57680657036212 ldrout = -2.90556504108222e-7
+ pscbe1 = 800072202.26248 lpscbe1 = -0.0363706622856625
+ pscbe2 = 9.4262349779212e-09 lpscbe2 = -5.49491994501789e-17
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.76670428794479 lbeta0 = 1.335799230126e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 6.60886646926599e-10 lagidl = -1.42315451584627e-16
+ bgidl = 718501708.2624 lbgidl = 141.799978991856
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.50479609548 lkt1 = -1.84562961557331e-9
+ kt2 = -0.0933453834719999 lkt2 = 1.9221133248501e-8
+ at = 63420.765808 lat = 0.000795512377238738
+ ute = -0.296816635519999 lute = 2.83030624703963e-8
+ ua1 = 7.1217460044e-10 lua1 = -7.85645160734429e-17
+ ub1 = 6.6569999932e-19 lub1 = -5.75212709274614e-26
+ uc1 = 4.84222600591201e-11 luc1 = -1.21411037663607e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.79 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.809177898371427+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -3.87991000155228e-8
+ k1 = -0.859188811758429 lk1 = 3.65232029360011e-7
+ k2 = 0.497540891920585 lk2 = -1.30539595977775e-07 wk2 = 5.29395592033938e-23
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 340167.983973857 lvsat = -0.0485861127225687
+ ua = 4.63603676662857e-10 lua = -5.16713597743197e-16
+ ub = -3.74312666585638e-20 lub = 4.1626996175928e-25
+ uc = -4.00506840596299e-13 luc = 1.1568680925945e-19 wuc = 1.92592994438724e-34 puc = -4.59177480789956e-41
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0115960246397143 lu0 = -1.54353259881862e-09 wu0 = -1.32348898008484e-23
+ a0 = 0.0905905090000019 la0 = 1.83073305009903e-7
+ keta = -0.107328375378326 lketa = 2.47031225828439e-08 wketa = -2.64697796016969e-23 pketa = 1.26217744835362e-29
+ a1 = 0.0
+ a2 = 0.0957216198444275 la2 = 1.08598140161593e-7
+ ags = -1.75201096157886 lags = 5.51568480003768e-7
+ b0 = 0.0
+ b1 = -5.53126201684571e-24 lb1 = 1.40346370532031e-30
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.146888130688428+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -6.20224638973626e-8
+ nfactor = {0.460556511571433+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 5.21754590359447e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 1.22133747383557 leta0 = -1.85564451248721e-7
+ etab = 0.0825970448787428 letab = -2.09734543007181e-08 wetab = 8.89219158494505e-24 petab = -4.93038065763132e-30
+ dsub = 1.569009795062 ldsub = -2.38765164747897e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.67677212549386 lpclm = -1.00526085236927e-8
+ pdiblc1 = 1.274858227734 lpdiblc1 = -2.06261564690401e-7
+ pdiblc2 = 0.03404075974251 lpdiblc2 = -5.82909086062429e-9
+ pdiblcb = -0.618713571428571 lpdiblcb = 9.98981256192857e-08 ppdiblcb = -1.0097419586829e-28
+ drout = -1.060023465579 ldrout = 3.78494291401226e-07 pdrout = 2.01948391736579e-28
+ pscbe1 = 799742134.776859 lpscbe1 = 0.0473783510437897
+ pscbe2 = 8.74071651536286e-09 lpscbe2 = 1.18989456610131e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 10.6076192291829 lbeta0 = -3.33520947772548e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1997599084.17429 lbgidl = -182.749235490393
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.181324352428573 lkt1 = -8.39210853952416e-8
+ kt2 = 0.251204129485714 lkt2 = -6.82024483227987e-08 pkt2 = 1.26217744835362e-29
+ at = 86010.6999428573 lat = -0.00493629938060092
+ ute = -0.104191251857142 lute = -2.05723540025316e-8
+ ua1 = 1.06408379028571e-09 lua1 = -1.67855490540565e-16
+ ub1 = 4.39e-19
+ uc1 = -3.96221633285712e-13 luc1 = 2.45756048898484e-19
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.80 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.07478710999828+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 1.00020772643138e-08 wvth0 = 3.09009195638845e-07 pvth0 = -5.67751865423132e-14
+ k1 = -5.1286956204091 lk1 = 1.14968132383383e-06 wk1 = 4.50044014538965e-06 pk1 = -8.26879369232878e-13
+ k2 = 1.71253150513387 lk2 = -3.53773466315292e-07 wk2 = -1.24766979955512e-06 pk2 = 2.29238115281662e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 196599.062727445 lvsat = -0.0222077641152017 wvsat = 0.0382634794636934 pvsat = -7.03026387230283e-9
+ ua = 1.09499195020051e-08 lua = -2.44339586328081e-15 wua = -9.97349657282265e-15 pua = 1.83246044581443e-21
+ ub = -1.10176987810022e-17 lub = 2.43370745297217e-24 wub = 9.71742714167601e-24 pub = -1.78541204102156e-30
+ uc = -1.95046650906367e-12 luc = 4.00465549025965e-19 wuc = 2.23051236992751e-18 puc = -4.09818729263891e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0305045071030862 lu0 = -5.01764480726134e-09 wu0 = -2.07694281434273e-08 pu0 = 3.81602934107632e-15
+ a0 = 11.8945952872442 la0 = -1.98571190491125e-06 wa0 = -9.23003228336598e-06 pa0 = 1.69586152151968e-12
+ keta = 2.8725060656273 lketa = -5.22790798766443e-07 wketa = -2.78676626918679e-06 pketa = 5.12020926936497e-13
+ a1 = 0.0
+ a2 = -0.915692431984333 la2 = 2.94428278146248e-7
+ ags = -17.4584307788897 lags = 3.43735611229775e-06 wags = 1.92777694860391e-05 pags = -3.54196242097841e-12
+ b0 = 1.64909602410302e-08 lb0 = -3.02993359796521e-15 wb0 = -1.43542628027125e-14 pb0 = 2.63735176753078e-21
+ b1 = -2.72213547111387e-09 lb1 = 5.00146116514166e-16 wb1 = 2.3694343668197e-15 pb1 = -4.35343284518884e-22
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.671987908673984+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 3.44556936112566e-08 wvoff = 2.29382665064214e-08 pvoff = -4.21451652002409e-15
+ nfactor = {22.646881443356+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -3.55460544833213e-06 wnfactor = -2.23985273805635e-05 pnfactor = 4.11534863121308e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 1.19292230047207 leta0 = -1.80343646201125e-07 weta0 = -1.70281446230248e-06 peta0 = 3.12863209602221e-13
+ etab = -1.35054831533076 letab = 2.42342642166654e-07 wetab = 1.19251224702015e-06 petab = -2.19103852681754e-13
+ dsub = 0.110567598564005 ldsub = 2.919879534127e-08 wdsub = 1.80646712572534e-07 pdsub = -3.31907624410895e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -3.21037297476804 lpclm = 7.04144222182726e-07 wpclm = 4.83782521566382e-06 ppclm = -8.8886814034956e-13
+ pdiblc1 = 0.832472285528334 lpdiblc1 = -1.24980668371127e-07 wpdiblc1 = 8.470329472543e-22
+ pdiblc2 = 0.01197382863821 lpdiblc2 = -1.77466740803794e-9
+ pdiblcb = -0.459207391761761 lpdiblcb = 7.05915767105635e-8
+ drout = 1.0
+ pscbe1 = -62925658.37043 lpscbe1 = 158.547919989374 wpscbe1 = 889.186384591092 ppscbe1 = -0.000163372882000075
+ pscbe2 = -6.5697022353171e-09 lpscbe2 = 2.93201862492883e-15 wpscbe2 = 1.65081203815177e-14 ppscbe2 = -3.03308648205739e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 16.956339511641 lbeta0 = -1.49999037142943e-06 wbeta0 = -2.74606535724672e-07 pbeta0 = 5.04542826282924e-14
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -2.35747138643738e-08 lagidl = 4.349826202443e-15 wagidl = 2.00658446261473e-14 pagidl = -3.68675783069593e-21
+ bgidl = 1018087901.40667 lbgidl = -2.7807073469512
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.270760618666671 lkt1 = -6.74886918905166e-8
+ kt2 = -0.12
+ at = 254051.821833334 lat = -0.0358109988289039
+ ute = -0.235274136333333 lute = 3.51189761093237e-9
+ ua1 = 3.70235701333335e-10 lua1 = -4.03726996130774e-17
+ ub1 = 7.98171532333335e-19 lub1 = -6.59916631502001e-26
+ uc1 = -3.50303784483333e-11 luc1 = 6.60919358299763e-18 wuc1 = 1.23259516440783e-32 puc1 = -1.46936793852786e-39
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.81 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.9572343898185+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = -4.53474374450263e-8
+ k1 = 0.53569697239527 wk1 = -3.82354338127103e-8
+ k2 = 0.0019675153606175 wk2 = -3.88017989862948e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 158306.030778317 wvsat = -0.0897138920691308
+ ua = -3.04440037815081e-09 wua = 1.42937786804482e-15
+ ub = 2.17119171108135e-18 wub = -6.00563149227904e-25
+ uc = 5.8607676477916e-11 wuc = -8.48882670463519e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.0033462673844341 wu0 = 9.01941200165266e-9
+ a0 = 1.1024195284682 wa0 = 9.95674089300636e-8
+ keta = 0.0040678945416715 wketa = 2.23904996628595e-9
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.45201457917293 wags = -1.45518340921094e-7
+ b0 = 2.0495112354e-07 wb0 = -1.78396057355394e-13
+ b1 = -1.39285641711e-09 wb1 = 1.21238707542917e-15
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.13442087482445+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = -1.30624050007531e-7
+ nfactor = {0.824618722274099+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor = 7.04427790632126e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0017402344
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00033736812078709 wpdiblc2 = 7.8792085111712e-10
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 833131390.92478 wpscbe1 = -28.8514335493783
+ pscbe2 = 1.49760924337686e-08 wpscbe2 = -3.65940266866235e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.352161e-10 walpha0 = 2.9178288739842e-16
+ alpha1 = -3.352161e-10 walpha1 = 2.9178288739842e-16
+ beta0 = 120.508347 wbeta0 = -7.87813795975734e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.29414875946086e-09 wagidl = 2.99503246679646e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.61265322 wkt1 = 5.83565774796837e-8
+ kt2 = -0.052484
+ at = 10000.0
+ ute = -1.2595
+ ua1 = -2.5605e-10
+ ub1 = 4.9434e-19
+ uc1 = 8.1951e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.82 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.9572343898185+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = -4.53474374450254e-8
+ k1 = 0.53569697239527 wk1 = -3.82354338127099e-8
+ k2 = 0.0019675153606175 wk2 = -3.88017989862948e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 158306.030778317 wvsat = -0.0897138920691308
+ ua = -3.04440037815081e-09 wua = 1.42937786804482e-15
+ ub = 2.17119171108135e-18 wub = -6.00563149227903e-25
+ uc = 5.86076764779161e-11 wuc = -8.48882670463519e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.0033462673844341 wu0 = 9.01941200165266e-9
+ a0 = 1.1024195284682 wa0 = 9.95674089300636e-8
+ keta = 0.0040678945416715 wketa = 2.23904996628594e-9
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.45201457917293 wags = -1.45518340921094e-7
+ b0 = 2.0495112354e-07 wb0 = -1.78396057355394e-13
+ b1 = -1.39285641711e-09 wb1 = 1.21238707542917e-15
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.13442087482445+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = -1.30624050007531e-7
+ nfactor = {0.824618722274099+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor = 7.04427790632125e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0017402344
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00033736812078709 wpdiblc2 = 7.8792085111712e-10
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 833131390.924781 wpscbe1 = -28.8514335493783
+ pscbe2 = 1.49760924337686e-08 wpscbe2 = -3.65940266866235e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.352161e-10 walpha0 = 2.9178288739842e-16
+ alpha1 = -3.352161e-10 walpha1 = 2.9178288739842e-16
+ beta0 = 120.508347 wbeta0 = -7.87813795975734e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.29414875946086e-09 wagidl = 2.99503246679645e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.61265322 wkt1 = 5.83565774796837e-8
+ kt2 = -0.052484
+ at = 10000.0
+ ute = -1.2595
+ ua1 = -2.5605e-10
+ ub1 = 4.9434e-19
+ uc1 = 8.1951e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.83 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.803767503941558+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.22830797890052e-06 wvth0 = -1.79208920332374e-07 pvth0 = 1.07139156801441e-12
+ k1 = 0.664089130540597 lk1 = -1.02761655308897e-06 wk1 = -1.13389821594509e-07 pk1 = 6.01515653583976e-13
+ k2 = 0.00828562145384356 lk2 = -5.05684342358544e-08 wk2 = -2.02709409112943e-08 pk2 = 1.31187274812179e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 318291.572337945 lvsat = -1.28048155850367 wvsat = -0.21808683134919 pvsat = 1.02746273042281e-6
+ ua = -5.33075329062927e-09 lua = 1.829935825525e-14 wua = 2.92162459329878e-15 pua = -1.19435443590571e-20
+ ub = 1.25812904613413e-18 lub = 7.30790978250598e-24 wub = 4.80971847653579e-25 pub = -8.65631734519523e-30
+ uc = 1.11121790395146e-10 luc = -4.20308946525096e-16 wuc = -1.16959759087328e-16 puc = 2.56691659207598e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.0257110848295883 lu0 = 1.79002027424757e-07 wu0 = 2.63095996236154e-08 pu0 = -1.38386045246095e-13
+ a0 = 1.45067756329113 la0 = -2.78736432582746e-06 wa0 = -1.31922546983098e-07 pa0 = 1.85278379931071e-12
+ keta = 0.0297999939159457 lketa = -2.05952852921158e-07 wketa = -1.71812191391369e-08 pketa = 1.55434648707954e-13
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.192856447433508 lags = 2.07423249122116e-06 wags = 2.88483644078954e-08 pags = -1.3955845535429e-12
+ b0 = 7.05617342574457e-07 lb0 = -4.00719873927131e-12 wb0 = -6.14192055855239e-13 pb0 = 3.48799481446116e-18
+ b1 = -1.86011401954631e-09 lb1 = 3.73980509212036e-15 wb1 = 1.61910313828454e-15 pb1 = -3.25524677390553e-21
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.0463353984898642+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.4467249496828e-06 wvoff = -3.03776973951178e-07 pvoff = 1.38586977141426e-12
+ nfactor = {-1.14000080560518+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.57242901477318e-05 wnfactor = 2.08689383068581e-06 pnfactor = -1.1064889066157e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.17947409030897 lpclm = -9.42626732775589e-06 wpclm = -1.05673175978488e-06 ppclm = 8.45779885793833e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00375354045914309 lpdiblc2 = 2.73421312781871e-08 wpdiblc2 = 3.35194054078397e-09 ppdiblc2 = -2.05217290028364e-14
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 866293788.844594 lpscbe1 = -265.422978589948 wpscbe1 = -57.7298511101553 ppscbe1 = 0.000231135143618971
+ pscbe2 = 2.07109452206038e-08 lpscbe2 = -4.59002305001351e-14 wpscbe2 = -7.5455147779306e-15 ppscbe2 = 3.11034037306499e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -5.99336892238184e-10 lalpha0 = 2.11395230082289e-15 walpha0 = 5.21682129652045e-16 palpha0 = -1.84005215190033e-21
+ alpha1 = -6.70744927608712e-10 lalpha1 = 2.68548314998316e-15 walpha1 = 5.83837982977292e-16 palpha1 = -2.33753100630277e-21
+ beta0 = 189.848257890176 lbeta0 = -0.000554978133008765 wbeta0 = -0.000139137070781514 pbeta0 = 4.83070837266712e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -6.94185464414402e-09 lagidl = 2.91952639635328e-14 wagidl = 6.16072925504796e-15 pagidl = -2.53373918521226e-20
+ bgidl = 2079168106.13984 lbgidl = -8637.37338365895 wbgidl = -939.342668797136 pbgidl = 0.00751824791655971
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.534900784064941 lkt1 = -6.22309737323817e-07 wkt1 = -8.27936976732643e-08 pkt1 = 1.12972911520073e-12
+ kt2 = -0.184900132058433 lkt2 = 1.05982336588844e-06 wkt2 = 9.28316884299548e-08 pkt2 = -7.43000048132547e-13
+ at = -10036.9857713251 lat = 0.160370684238485 wat = -0.0219990954385094 pat = 1.76074886131347e-7
+ ute = -3.43606189231482 lute = 1.74206202440626e-05 wute = 8.58204186916902e-07 pute = -6.86883717156497e-12
+ ua1 = -7.6172834730993e-09 lua1 = 5.89173472693495e-14 wua1 = 4.51193148315825e-15 pua1 = -3.61122949054926e-20
+ ub1 = 6.83326414052414e-18 lub1 = -5.07350563280097e-23 wub1 = -4.20216384280999e-24 pub1 = 3.36329974201051e-29
+ uc1 = 2.15923921221768e-10 luc1 = -1.66260602146377e-15 wuc1 = -1.03974356336644e-16 puc1 = 8.3218298696536e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.84 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.28898644589216+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 7.14379111212181e-07 wvth0 = 2.39720780551531e-07 pvth0 = -6.05891100094613e-13
+ k1 = 0.313869860205983 lk1 = 3.74567896785643e-07 wk1 = 1.08272762688586e-07 pk1 = -2.85962149975529e-13
+ k2 = -0.0113967243124037 lk2 = 2.82344230258798e-08 wk2 = 2.14385089902605e-08 pk2 = -3.58062261705228e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -127615.224203281 lvsat = 0.504810197732726 wvsat = 0.138963898468592 pvsat = -4.02073059222729e-7
+ ua = 8.46782419676772e-10 lua = -6.43384532678076e-15 wua = -1.28923989157938e-15 pua = 4.91563273757763e-21
+ ub = 4.21132319453355e-18 lub = -4.51589108484764e-24 wub = -2.80255523416312e-24 pub = 4.49004838866801e-30
+ uc = -1.44139808872775e-11 luc = 8.23027636387965e-17 wuc = -4.32715490163555e-17 puc = -3.83362591644869e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0372827823004497 lu0 = -7.32085972013921e-08 wu0 = -2.36288594169527e-08 pu0 = 6.15542111837761e-14
+ a0 = 0.697811826347268 la0 = 2.26909069744023e-07 wa0 = 4.26710916603083e-07 pa0 = -3.8383543375358e-13
+ keta = -0.0401458857741497 lketa = 7.40917738081069e-08 wketa = 4.47575323451864e-08 pketa = -9.25515745886309e-14
+ a1 = 0.0
+ a2 = 0.8
+ ags = 1.49115277572598 lags = -3.12379936214226e-06 wags = -1.0689641089592e-06 pags = 2.99976347388858e-12
+ b0 = -7.94379697515045e-07 lb0 = 1.99838891003735e-12 wb0 = 6.91453667743355e-13 pb0 = -1.73946205541941e-18
+ b1 = 1.48459351569487e-08 lb1 = -6.31467552954354e-14 wb1 = -1.29223799997202e-14 pb1 = 5.49649691346675e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.434209696546482+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 4.7724930530236e-07 wvoff = 1.47548647392246e-07 pvoff = -4.21117512503914e-13
+ nfactor = {5.24464569723871+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -9.83812974903888e-06 wnfactor = -2.54196563594254e-06 pnfactor = 7.46782833274537e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.15964838675 leta0 = -3.18890874427738e-7
+ etab = -0.139629715253176 letab = 2.78778788739746e-07 wetab = -4.3556797369739e-15 petab = 1.74389787185995e-20
+ dsub = 0.86055995 ldsub = -1.20336179029335e-06 wdsub = -4.2351647362715e-22
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.8782865672848 lpclm = 6.81992292315401e-06 wpclm = 2.26435955491944e-06 ppclm = -4.83896403475676e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00618976065390853 lpdiblc2 = -1.24681915170744e-08 wpdiblc2 = -3.76675368368118e-09 ppdiblc2 = 7.9796219805642e-15
+ pdiblcb = 0.446683561701301 lpdiblcb = -2.68924164154103e-06 wpdiblcb = -5.84655000315499e-07 ppdiblcb = 2.34080251837817e-12
+ drout = 0.56
+ pscbe1 = 799999825.751094 lpscbe1 = 0.000349148282111855 wpscbe1 = 0.000116822077870893 ppscbe1 = -2.3408025170979e-10
+ pscbe2 = 9.64494290327994e-09 lpscbe2 = -1.59491184418896e-15 wpscbe2 = -9.63756888547083e-18 ppscbe2 = 9.31763464847991e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.43634373166531e-10 lalpha0 = 2.89441087032588e-16 walpha0 = 1.22365093396376e-16 palpha0 = -2.41293356381315e-22
+ alpha1 = 1.0816388134009e-14 lalpha1 = -4.37571965671298e-20 walpha1 = -6.86515990785695e-21 palpha1 = 2.78790641258702e-26
+ beta0 = 99.5562015493227 lbeta0 = -0.000193472847399029 wbeta0 = -3.69984222722852e-05 pbeta0 = 7.4134959654913e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.99964186932485e-10 lagidl = -1.80091157046962e-15 wagidl = -6.38513495194959e-16 pagidl = 1.88496072203575e-21
+ bgidl = -1158336212.27968 lbgidl = 4324.72949363981 wbgidl = 1878.68533759427 pbgidl = -0.00376438380755378
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.976517602574835 lkt1 = 1.14580609229925e-06 wkt1 = 4.56929630921825e-07 pkt1 = -1.03117898636527e-12
+ kt2 = 0.165175087925782 lkt2 = -3.41784344844624e-07 wkt2 = -1.5066748080005e-07 pkt2 = 2.31905611186206e-13
+ at = 161680.063572368 lat = -0.527138532881486 wat = -0.0509318848846585 pat = 2.91914050018946e-7
+ ute = 2.49214864685894 lute = -6.3143519225752e-06 wute = -1.51068616966579e-06 pute = 2.61556732246691e-12
+ ua1 = 1.48485670551999e-08 lua1 = -3.10299198638693e-14 wua1 = -9.44609384839589e-15 pua1 = 1.97719117292866e-20
+ ub1 = -1.32102875575673e-17 lub1 = 2.95139730428451e-23 wub1 = 9.07800588114452e-24 pub1 = -1.95372563492924e-29
+ uc1 = -5.13869094463099e-10 luc1 = 1.25929035860325e-15 wuc1 = 2.53938411663406e-16 puc1 = -6.00804173397788e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.85 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.853405309965567+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.58409185021411e-07 wvth0 = -1.39422741608603e-07 pvth0 = 1.53811286993877e-13
+ k1 = 0.653672335141335 lk1 = -3.06305535723996e-07 wk1 = -1.60840384701178e-07 pk1 = 2.53268744183204e-13
+ k2 = -0.0346845498984843 lk2 = 7.48970076509539e-08 wk2 = 3.40801518906036e-08 pk2 = -6.1136703224156e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 414226.002839943 lvsat = -0.580894949654276 wvsat = -0.292525898573937 pvsat = 4.62517286274688e-7
+ ua = -6.93410807565795e-09 lua = 9.15698172810778e-15 wua = 4.91832070271525e-15 pua = -7.52266127471013e-21
+ ub = 4.65797676531992e-18 lub = -5.41086558420014e-24 wub = -2.72291330550849e-24 pub = 4.33046722803907e-30
+ uc = 1.81806202337966e-10 luc = -3.10870092755669e-16 wuc = -1.94260915048072e-16 puc = 2.64206116202343e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.0180415821602378 lu0 = 3.76466575725148e-08 wu0 = 2.30691315939734e-08 pu0 = -3.20160944385199e-14
+ a0 = 3.54901848003353 la0 = -5.48614779206671e-06 wa0 = -1.64057505888433e-06 pa0 = 3.75845369576773e-12
+ keta = 0.160951848873145 lketa = -3.28854393329921e-07 wketa = -1.15433474702732e-07 pketa = 2.28428432536516e-13
+ a1 = 0.0
+ a2 = -0.545869846805198 la2 = 2.69676382574852e-06 wa2 = 1.17148845166831e-06 pa2 = -2.3473500697267e-12
+ ags = -4.28091834471354 lags = 8.44189002022939e-06 wags = 3.33278388649016e-06 pags = -5.82016424227718e-12
+ b0 = 3.36419783617054e-07 lb0 = -2.67431326689916e-13 wb0 = -2.92830612377317e-13 pb0 = 2.32780838039623e-19
+ b1 = -3.48964088427062e-08 lb1 = 3.65236208740251e-14 wb1 = 3.03749579210562e-14 pb1 = -3.17913356693436e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.259503986741162+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 1.27185709277017e-07 wvoff = -2.84184412274774e-09 pvoff = -1.19775121769102e-13
+ nfactor = {-0.319147594503196+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.31022647480301e-06 wnfactor = 1.74228708535462e-06 pnfactor = -1.11667022525755e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 1.30021981947533 leta0 = -2.60429149303676e-06 weta0 = -1.20077566296002e-06 peta0 = 2.40603382146987e-12
+ etab = -0.5255943379817 letab = 1.05214884013344e-06 wetab = 4.62737947120342e-07 petab = -9.27203286285926e-13
+ dsub = -1.0505222851039 ldsub = 2.62593674989809e-06 wdsub = 8.78616338751233e-07 pdsub = -1.76051255229503e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.71187071513153 lpclm = -2.37752669881392e-06 wpclm = -1.20010282898139e-06 ppclm = 2.10289357112401e-12
+ pdiblc1 = 0.425612538750144 lpdiblc1 = -7.13580191074433e-08 wpdiblc1 = -2.42179464636487e-08 ppdiblc1 = 4.8526298521446e-14
+ pdiblc2 = 0.000442038614921492 lpdiblc2 = -9.51291192728789e-10 wpdiblc2 = -1.97621721071068e-10 ppdiblc2 = 8.28034485727544e-16
+ pdiblcb = -2.4420486468052 lpdiblcb = 3.09900641280632e-06 wpdiblcb = 1.75505422646515e-06 ppdiblcb = -2.3473500697267e-12
+ drout = 0.130443268025862 ldrout = 8.60716999228736e-07 wdrout = 6.7016929833631e-08 pdrout = -1.34284033866331e-13
+ pscbe1 = 795949907.516755 lpscbe1 = 8.1153039617293 wpscbe1 = 3.52533091039368 ppscbe1 = -7.06382188107695e-6
+ pscbe2 = 1.13007831021364e-08 lpscbe2 = -4.91277349336426e-15 wpscbe2 = -8.38036654198051e-16 ppscbe2 = 2.59165404925861e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -9.87371464155049e-11 lalpha0 = 1.99479032183074e-16 walpha0 = 3.89361930508609e-18 palpha0 = -3.90815418595202e-24
+ alpha1 = -1.00395384042722e-10 lalpha1 = 2.01143460011354e-16 walpha1 = 1.41231166682103e-20 palpha1 = -1.41758382627833e-26
+ beta0 = -6.2085750409849 lbeta0 = 1.84515256925978e-05 wbeta0 = 2.85982267173492e-06 pbeta0 = -5.73032106150344e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.48486969965984e-09 lagidl = -3.17327934820334e-15 wagidl = -9.46639294590015e-16 pagidl = 2.50236255443501e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.311247690317049 lkt1 = -1.87217184798778e-07 wkt1 = -1.01566834621491e-07 pkt1 = 8.78988120272346e-14
+ kt2 = 0.067277764573018 lkt2 = -1.4562424743102e-07 wkt2 = -8.21617208244054e-08 pkt2 = 9.46383592329287e-14
+ at = -58472.4666282348 lat = -0.0860116430850422 wat = 0.0438554898297 pat = 1.0198545932042e-7
+ ute = 3.28580422869586 lute = -7.90462580253604e-06 wute = -3.37845974068789e-06 pute = 6.35808686325173e-12
+ ua1 = 3.14855775363349e-09 lua1 = -7.5862251260138e-15 wua1 = -2.79790854509362e-15 pua1 = 6.45072344694485e-21
+ ub1 = -6.89547190920106e-19 lub1 = 4.42575238576196e-24 wub1 = 1.48321931002245e-24 pub1 = -4.3193318687783e-30
+ uc1 = 1.36761881436912e-11 luc1 = 2.02230466849702e-16 wuc1 = 5.4552685093815e-17 puc1 = -2.01288413341321e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.86 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.06559072440258+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.45683175676997e-08 wvth0 = 3.16605444498152e-08 pvth0 = -1.79106529713978e-14
+ k1 = 0.279778588885957 lk1 = 6.89839558861536e-08 wk1 = 1.02635906735711e-07 pk1 = -1.11911042496189e-14
+ k2 = 0.0588673796765528 lk2 = -1.90041512771867e-08 wk2 = -3.08753756106278e-08 pk2 = 4.06130326123736e-15
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -417535.606324964 lvsat = 0.253971625597644 wvsat = 0.335682255406013 pvsat = -1.68035968744068e-7
+ ua = 3.27985481686099e-09 lua = -1.09510988788893e-15 wua = -3.20716570595157e-15 pua = 6.33157574720239e-22
+ ub = -1.2345664485046e-18 lub = 5.03674493441592e-25 wub = 1.82803590324448e-24 pub = -2.37470674110175e-31
+ uc = -2.05398107231978e-10 luc = 7.77796505018991e-17 wuc = 1.12838381188201e-16 puc = -4.40395817067802e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0252294278132964 lu0 = -5.78588308125063e-09 wu0 = -1.21087937565205e-08 pu0 = 3.29315010730734e-15
+ a0 = -5.09656835597266 la0 = 3.19171301959828e-06 wa0 = 4.3149307166307e-06 pa0 = -2.21928398280729e-12
+ keta = -0.219406486011187 lketa = 5.29238192185339e-08 wketa = 1.54108497140403e-07 pketa = -4.21197394875099e-14
+ a1 = 0.0
+ a2 = 3.4917396936104 la2 = -1.35591811108145e-06 wa2 = -2.34297690333663e-06 pa2 = 1.18023478444847e-12
+ ags = 5.34930966039938 lags = -1.22428762602661e-06 wags = -3.54133849490585e-06 pags = 1.07961923796858e-12
+ b0 = 3.36411426106461e-08 lb0 = 3.64775869833687e-14 wb0 = -2.92823337730985e-14 pb0 = -3.1751266288625e-20
+ b1 = 1.20971893018223e-09 lb1 = 2.82708926160482e-16 wb1 = -1.05297830978017e-15 pb1 = -2.46078952557506e-22
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0754758328357337+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -5.75294217269406e-08 wvoff = -1.62918018506628e-07 pvoff = 4.08986169737536e-14
+ nfactor = {0.469571439275535+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.18563152871185e-07 wnfactor = 8.33879002528737e-07 pnfactor = -2.04871055058488e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -3.09209424595066 leta0 = 1.80441908079547e-06 weta0 = 2.40155132592004e-06 peta0 = -1.20974065405968e-12
+ etab = 1.04919121363861 letab = -5.28515385951068e-07 wetab = -9.25475876817968e-07 petab = 4.66192739857146e-13
+ dsub = 2.75642785955825 ldsub = -1.19522473965408e-06 wdsub = -1.69911431618369e-06 pdsub = 8.26840771174766e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.93429263062313 lpclm = 1.28224777471044e-06 wpclm = 1.78344240667025e-06 ppclm = -8.91789238892313e-13
+ pdiblc1 = 0.693913943651026 lpdiblc1 = -3.4066099315282e-07 wpdiblc1 = -7.2151428122984e-08 ppdiblc1 = 9.66387158678163e-14
+ pdiblc2 = -0.000186043231205704 lpdiblc2 = -3.2086471707e-10 wpdiblc2 = 7.09252736409427e-11 ppdiblc2 = 5.58485005084273e-16
+ pdiblcb = 0.6454322 wpdiblcb = -5.8356577479684e-7
+ drout = 0.419898155164671 ldrout = 5.70181576996237e-07 wdrout = 3.49865747236643e-07 pdrout = -4.18188725904707e-13
+ pscbe1 = 808100184.96649 lpscbe1 = -4.08033047372464 wpscbe1 = -7.05066182078826 ppscbe1 = 3.55165103097096e-6
+ pscbe2 = -2.46149064829988e-08 lpscbe2 = 3.11369893609922e-14 wpscbe2 = 2.79501864077822e-14 ppscbe2 = -2.6304035449412e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 15.4316782236305 lbeta0 = -3.2695106374544e-06 wbeta0 = -5.79924331280747e-06 pbeta0 = 2.96106921635925e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.9155002283657e-09 lagidl = 2.24725016076352e-15 wagidl = 3.25111379885939e-15 pagidl = -1.71106075131224e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.490171920067543 lkt1 = -7.62503089862371e-09 wkt1 = -2.53311065945011e-08 pkt1 = 1.13784960275199e-14
+ kt2 = -0.169525802550641 lkt2 = 9.20633074087115e-08 wkt2 = 8.43432458108742e-08 pkt2 = -7.24881704428004e-14
+ at = -351850.595451777 lat = 0.208461666293399 wat = 0.289363671341388 pat = -1.4443920423285e-7
+ ute = -8.46880084627034 lute = 3.89385921317499e-06 wute = 5.49717471965438e-06 pute = -2.55068034053099e-12
+ ua1 = -1.02354812241228e-08 lua1 = 5.84777646924651e-15 wua1 = 8.00135956934344e-15 pua1 = -4.3888583353634e-21
+ ub1 = 6.65993281761436e-18 lub1 = -2.95116323164436e-24 wub1 = -5.44206201660692e-24 pub1 = 2.63180153304338e-30
+ uc1 = 4.07413843287467e-10 luc1 = -1.92977010960725e-16 wuc1 = -2.93064166148101e-16 puc1 = 1.47626091606281e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.87 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.952362636419151+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -2.46840687645923e-09 wvth0 = -7.84876773623398e-09 pvth0 = 1.99149138401781e-15
+ k1 = 0.250760756861332 lk1 = 8.36011954654138e-08 wk1 = 1.62039955832326e-07 pk1 = -4.11148841132035e-14
+ k2 = 0.059785373350045 lk2 = -1.9466574984316e-08 wk2 = -4.5966569284924e-08 pk2 = 1.16632355243716e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 23677.7266467225 lvsat = 0.0317179097398172 wvsat = 0.00423304327347462 pvsat = -1.07406276890852e-9
+ ua = 3.82457305850162e-09 lua = -1.36950244190529e-15 wua = -3.92959051134346e-15 pua = 9.97066789214711e-22
+ ub = -2.09995912615671e-18 lub = 9.39601343133321e-25 wub = 2.73348534215552e-24 pub = -6.93575436321147e-31
+ uc = -1.02800877021846e-10 luc = 2.60980399364586e-17 wuc = 5.12033382571833e-17 puc = -1.29919766260099e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0220970030333385 lu0 = -4.20797734956808e-09 wu0 = -1.12257955921839e-08 pu0 = 2.8483547929916e-15
+ a0 = 1.67337698123642 la0 = -2.1853185495006e-07 wa0 = -1.82843952507028e-07 pa0 = 4.63935446014657e-14
+ keta = -0.220275360449258 lketa = 5.33614999458468e-08 wketa = 1.42039184410068e-07 pketa = -3.60400283779197e-14
+ a1 = 0.0
+ a2 = 1.08040210428168 la2 = -1.41247793196123e-7
+ ags = 5.45324277778348 lags = -1.27664216704586e-06 wags = -2.81707930434329e-06 pags = 7.14785983128938e-13
+ b0 = 2.13694962696229e-07 lb0 = -5.42214639698024e-14 wb0 = -1.86006976508597e-13 pb0 = 4.71961081704558e-20
+ b1 = 3.56833708807187e-09 lb1 = -9.05404874367741e-16 wb1 = -3.10599550191199e-15 pb1 = 7.88093556686637e-22
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.0149749621301876+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -1.03092472027509e-07 wvoff = -1.64674260970583e-07 pvoff = 4.1783294258849e-14
+ nfactor = {0.465955227927072+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 5.2038475786238e-07 wnfactor = 8.60725266089283e-07 pnfactor = -2.18394403940632e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = 5.0839925e-05 letab = -2.8758079190025e-11 wetab = -6.46234853557053e-27 petab = 4.62223186652937e-33
+ dsub = 0.135738150968819 ldsub = 1.24903149322799e-07 wdsub = -1.16236722637567e-07 pdsub = 2.94930923449978e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.584855727258072 lpclm = 1.32696149498674e-08 wpclm = 2.63582197876433e-08 ppclm = -6.687950181378e-15
+ pdiblc1 = -0.433302714331551 lpdiblc1 = 2.27155235622718e-07 wpdiblc1 = 2.41174642100564e-07 ppdiblc1 = -6.11939654641024e-14
+ pdiblc2 = -0.0128910162527078 lpdiblc2 = 6.0790494579703e-09 wpdiblc2 = 2.37684962380499e-09 ppdiblc2 = -6.0308518559691e-16
+ pdiblcb = 1.5288616936104 lpdiblcb = -4.45012589104848e-07 wpdiblcb = -1.17584535374295e-06 ppdiblcb = 2.98350769141259e-13
+ drout = 2.68866710792933 ldrout = -5.72672213886763e-07 wdrout = -9.67799213807808e-07 pdrout = 2.45562597917097e-13
+ pscbe1 = 800072202.262481 lpscbe1 = -0.0363706622858899
+ pscbe2 = 6.56034039735564e-08 lpscbe2 = -1.43089508202197e-14 wpscbe2 = -4.88984167986425e-14 ppscbe2 = 1.240714198957e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.58381130825585 lbeta0 = 1.79985907428027e-07 wbeta0 = 1.5919593867522e-07 pbeta0 = -4.03932631078819e-14
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.98040736912706e-10 lagidl = -2.27862570299072e-16 wagidl = -2.93469776285604e-16 pagidl = 7.44629667462753e-23
+ bgidl = 718501708.2624 lbgidl = 141.799978991856
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.498446981600032 lkt1 = -3.45660932767902e-09 wkt1 = -5.52647316259135e-09 pkt1 = 1.40224861496388e-15
+ kt2 = 0.0445249489938775 lkt2 = -1.57611198190635e-08 wkt2 = -1.20006776803005e-07 pkt2 = 3.04496794985569e-14
+ at = 57341.8269867532 lat = 0.00233793976117014 wat = 0.00529130409184325 pat = -1.34257846113567e-9
+ ute = -1.30058452243721 lute = 2.8299209972156e-07 wute = 8.73711890098697e-07 pute = -2.21689539010413e-13
+ ua1 = 2.35875649582172e-09 lua1 = -4.96356680134332e-16 wua1 = -1.43323790167728e-15 pua1 = 3.63659752506281e-22
+ ub1 = 1.16910367748392e-18 lub1 = -1.85251396399027e-25 wub1 = -4.3817877107231e-25 pub1 = 1.1118041412049e-31
+ uc1 = 4.842226005912e-11 luc1 = -1.21411037663607e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.88 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.519906045771481+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.12196914991265e-07 wvth0 = -2.51791535056647e-07 pvth0 = 6.38878215645287e-14
+ k1 = -2.14640553063249 lk1 = 6.91841389090084e-07 wk1 = 1.12043488048633e-06 pk1 = -2.84291303530438e-13
+ k2 = 0.742351439930847 lk2 = -1.92656110756063e-07 wk2 = -2.13090983887778e-07 pk2 = 5.40682146147976e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 718646.288864315 lvsat = -0.144618548457339 wvsat = -0.329439703578072 pvsat = 8.35897243079749e-8
+ ua = -6.73429065317341e-10 lua = -2.28210869022336e-16 wua = 9.89709911073852e-16 pua = -2.51122064866502e-22
+ ub = 2.17252667570044e-18 lub = -1.444692968293e-25 wub = -1.92361855367503e-24 pub = 4.88085506479626e-31
+ uc = -1.75358786644502e-12 luc = 4.59008117191125e-19 wuc = 1.17776529410776e-18 puc = -2.98837921369845e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0114035110851051 lu0 = -1.49468555706697e-09 wu0 = 1.67569996868308e-10 pu0 = -4.25180380153854e-17
+ a0 = 1.9708531515954 la0 = -2.94011376083755e-07 wa0 = -1.63664114857212e-06 pa0 = 4.15269868550651e-13
+ keta = 0.185247310731128 lketa = -4.95329839807661e-08 wketa = -2.54667298126761e-07 pketa = 6.46174975555975e-14
+ a1 = 0.0
+ a2 = -0.0642388429300809 la2 = 1.49185388262758e-07 wa2 = 1.39234737525835e-07 pa2 = -3.53284476566427e-14
+ ags = -1.75201096157886 lags = 5.51568480003768e-07 pags = -1.0097419586829e-28
+ b0 = 4.84829725760104e-07 lb0 = -1.23017300806288e-13 wb0 = -4.22011404818764e-13 pb0 = 1.07078219778879e-19
+ b1 = 1.20004221723718e-07 lb1 = -3.04490311906242e-14 wb1 = -1.04455538724264e-13 pb1 = 2.65038172071237e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.202474522747349+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -1.50667298041583e-07 wvoff = -3.04096503027941e-07 pvoff = 7.71593180027886e-14
+ nfactor = {8.86283963789837+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -1.61018191413287e-06 wnfactor = -7.31361778667162e-06 pnfactor = 1.85570618186555e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.449680676841319 leta0 = 1.02303428230211e-08 weta0 = 6.71674923452659e-07 peta0 = -1.70426093352414e-13
+ etab = -0.509844467228317 letab = 1.29348507890743e-07 wetab = 5.15680168754675e-07 petab = -1.3084507625863e-13
+ dsub = 1.49522316817639 ldsub = -2.20043062548331e-07 wdsub = 6.42262559706178e-08 pdsub = -1.62963206061928e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.7113217975759 lpclm = -1.88190004700855e-08 wpclm = -3.00731470796508e-08 ppclm = 7.63054982796072e-15
+ pdiblc1 = 1.42365132059164 lpdiblc1 = -2.44015282520449e-07 wpdiblc1 = -1.2951429916088e-07 ppdiblc1 = 3.28620516689877e-14
+ pdiblc2 = 0.0434275473326668 lpdiblc2 = -8.21082863623756e-09 wpdiblc2 = -8.17056217303294e-09 ppdiblc2 = 2.07314125185017e-15
+ pdiblcb = 0.0411311718817835 lpdiblcb = -6.75262606350806e-08 wpdiblcb = -5.74350111578068e-07 ppdiblcb = 1.45731576861038e-13
+ drout = -1.060023465579 ldrout = 3.78494291401226e-07 pdrout = 1.0097419586829e-28
+ pscbe1 = 799742134.776855 lpscbe1 = 0.0473783510437897
+ pscbe2 = -6.50649866333954e-08 lpscbe2 = 1.8845931933654e-14 wpscbe2 = 6.42428605643206e-14 ppscbe2 = -1.63005337395668e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.94602021912431 lbeta0 = 5.95547553846634e-07 wbeta0 = 3.1871736818431e-06 pbeta0 = -8.08691139815094e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.98303042219644e-08 lagidl = -1.00808892811517e-14 wagidl = -3.45825361105938e-14 pagidl = 8.7747306349493e-21
+ bgidl = 1971613273.74545 lbgidl = -176.155777852855 wbgidl = 22.6188861403498 pbgidl = -5.73915783704968e-6
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.0451218924034116 lkt1 = -1.18480144184805e-07 wkt1 = -1.18555006925112e-07 pkt1 = 3.00813175721293e-14
+ kt2 = 0.251204129485714 lkt2 = -6.82024483227987e-08 wkt2 = -2.64697796016969e-23 pkt2 = -6.31088724176809e-30
+ at = 403130.148536321 lat = -0.0853999684305664 wat = -0.276030979301996 pat = 7.00381684712334e-8
+ ute = 0.635331794984893 lute = -2.08213755246902e-07 wute = -6.43704672613416e-07 pute = 1.6332911769622e-13
+ ua1 = 1.19632687647293e-09 lua1 = -2.01409925528107e-16 wua1 = -1.1510864044473e-16 pua1 = 2.92068606659631e-23
+ ub1 = -1.44875661968324e-19 lub1 = 1.48148523338208e-25 wub1 = 5.08224176973543e-25 pub1 = -1.28953245096028e-31
+ uc1 = 2.05303367647542e-10 luc1 = -5.19470178380938e-17 wuc1 = -1.79047546036807e-16 puc1 = 4.54302709985572e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.89 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.936922071118865+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -3.55773096061138e-08 wvth0 = 1.89007026543953e-07 pvth0 = -1.71014205540347e-14
+ k1 = 2.88672063246468 lk1 = -2.32909980234248e-07 wk1 = -2.47643625751504e-06 pk1 = 3.76572621267967e-13
+ k2 = -0.0980947878816334 lk2 = -3.82384039813927e-08 wk2 = 3.28357628052207e-07 pk2 = -4.54137632027716e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 68505.2416768007 lvsat = -0.0251661834344357 wvsat = 0.149760465927212 pvsat = -4.45516043573942e-9
+ ua = 2.43829787634319e-09 lua = -7.99937795194454e-16 wua = -2.56470703563015e-15 pua = 4.01941624002264e-22
+ ub = -4.08637341556229e-18 lub = 1.00549719363868e-24 wub = 3.68417835492037e-24 pub = -5.42251842927331e-31
+ uc = 3.5829983239602e-12 luc = -5.21498873330598e-19 wuc = -2.58599359830409e-18 puc = 3.92688791209661e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00826126749341798 lu0 = -9.17351715235518e-10 wu0 = -1.40819615485656e-09 pu0 = 2.47002204339477e-16
+ a0 = -2.91171647385821 la0 = 6.03077788909712e-07 wa0 = 3.65785823673631e-06 pa0 = -5.57504387010223e-13
+ keta = -2.67438764390233 lketa = 4.75876325138903e-07 wketa = 2.04142862556525e-06 pketa = -3.57251094792106e-13
+ a1 = 0.0
+ a2 = -0.542451352177139 la2 = 2.37048807224249e-07 wa2 = -3.2488105422695e-07 pa2 = 4.99449391094714e-14
+ ags = 16.2167446231118 lags = -2.7498848898382e-06 wags = -1.0034187524511e-05 pags = 1.84361137644098e-12
+ b0 = 7.09541097323297e-06 lb0 = -1.33759922514822e-12 wb0 = -6.17607418333531e-12 pb0 = 1.16428943626406e-18
+ b1 = -2.30638774816275e-07 lb1 = 3.39756584926584e-14 wb1 = 2.00755416168635e-13 pb1 = -2.95735071682133e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.37054951230353+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = 1.3834912699042e-07 wvoff = 6.30988779989219e-07 pvoff = -9.46467063018033e-14
+ nfactor = {-12.2125615188319+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 2.26206476659666e-06 wnfactor = 7.94425424778819e-06 pnfactor = -9.47668420641852e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.120015691344427 leta0 = 7.08006796033221e-08 weta0 = -7.68922002124965e-07 peta0 = 9.425910157474e-14
+ etab = 2.11494309327531 letab = -3.5291158496327e-07 wetab = -1.82396306385392e-06 petab = 2.99024593798246e-13
+ dsub = 0.572662647396033 ldsub = -5.05382503837928e-08 wdsub = -2.21575697391435e-07 pdsub = 3.62149296908775e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.19100937701794 lpclm = -1.06953438503709e-07 wpclm = 1.00672029215758e-06 ppclm = -1.82862619143413e-13
+ pdiblc1 = 0.317803627914611 lpdiblc1 = -4.08345684018201e-08 wpdiblc1 = 4.47984171917759e-07 ppdiblc1 = -7.3243474917704e-14
+ pdiblc2 = -0.0136219297357493 lpdiblc2 = 2.27104293397374e-09 wpdiblc2 = 2.22793722721138e-08 ppdiblc2 = -3.52151655355998e-15
+ pdiblcb = -2.1041531953047 lpdiblcb = 3.26633272001194e-07 wpdiblcb = 1.43181379465865e-06 ppdiblcb = -2.22866936123553e-13
+ drout = 1.0
+ pscbe1 = 1489778636.75105 lpscbe1 = -126.735098266179 wpscbe1 = -462.337430960944 ppscbe1 = 8.49466432027474e-5
+ pscbe2 = 1.88620777492216e-07 lpscbe2 = -2.77645145664369e-14 wpscbe2 = -1.53391958306774e-13 ppscbe2 = 2.36861644360761e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 32.8981065745096 lbeta0 = -4.17270712848737e-06 wbeta0 = -1.41508339121449e-05 pbeta0 = 2.37687300945109e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -6.74215300284889e-08 lagidl = 9.62481198118684e-15 wagidl = 5.82315252828736e-14 pagidl = -8.27827530705665e-21
+ bgidl = 1078721459.07394 lbgidl = -12.1020860678145 wbgidl = -52.7774009941531 pbgidl = 8.11362818703377e-6
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.588566358725377 lkt1 = -1.86314620540717e-08 wkt1 = 2.76628349491928e-07 pkt1 = -4.25269060524426e-14
+ kt2 = -0.12
+ at = -130379.210681383 lat = 0.0126233066665801 wat = 0.334621149380057 pat = -4.21587790879062e-8
+ ute = -1.43054535004171 lute = 1.71356050240271e-07 wute = 1.04040255214486e-06 pute = -1.46096955030291e-13
+ ua1 = 1.21327663024821e-09 lua1 = -2.04524154638499e-16 wua1 = -7.33809970445416e-16 pua1 = 1.42882712130979e-22
+ ub1 = 2.16054807692609e-18 lub1 = -2.75433896480079e-25 wub1 = -1.18585641293827e-24 pub1 = 1.8230526393024e-31
+ uc1 = -5.14996086770266e-10 luc1 = 8.03957618204534e-17 wuc1 = 4.17777607419219e-16 puc1 = -6.42262049213788e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.90 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0248735+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.47866595
+ k2 = -0.0038200645
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 24491.02
+ ua = -9.1237589e-10
+ ub = 1.27540665e-18
+ uc = -6.8009552e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0101068633
+ a0 = 1.2509318
+ keta = 0.0074076058
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.23496304
+ b0 = -6.114e-8
+ b1 = 4.1551e-10
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.32925646+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.8753257+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0017402344
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00083787503
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 790097310.0
+ pscbe2 = 9.5178184e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.1731672e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.52561
+ kt2 = -0.052484
+ at = 10000.0
+ ute = -1.2595
+ ua1 = -2.5605e-10
+ ub1 = 4.9434e-19
+ uc1 = 8.1951e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.91 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.0248735+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.47866595
+ k2 = -0.0038200645
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 24491.02
+ ua = -9.1237589e-10
+ ub = 1.27540665e-18
+ uc = -6.8009552e-11
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0101068633
+ a0 = 1.2509318
+ keta = 0.0074076058
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.23496304
+ b0 = -6.114e-8
+ b1 = 4.1551e-10
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.32925646+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.8753257+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0017402344
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00083787503
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 790097310.0
+ pscbe2 = 9.5178184e-9
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.1731672e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.52561
+ kt2 = -0.052484
+ at = 10000.0
+ ute = -1.2595
+ ua1 = -2.5605e-10
+ ub1 = 4.9434e-19
+ uc1 = 8.1951e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.92 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.07107107368712+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.6975304503957e-7
+ k1 = 0.494959691956788 lk1 = -1.30410760193024e-7
+ k2 = -0.0219500099959799 lk2 = 1.45107243054376e-07 wk2 = 6.61744490042422e-24
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -7001.32282608497 lvsat = 0.25205630352445 pvsat = -1.05879118406788e-22
+ ua = -9.72930690075804e-10 lua = 4.84664451675117e-16
+ ub = 1.97553469528639e-18 lub = -5.60363794028421e-24
+ uc = -6.33324781905928e-11 luc = -3.74340499917891e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0135316598112797 lu0 = -2.74111568556144e-8
+ a0 = 1.25390517231245 la0 = -2.37980780984495e-8
+ keta = 0.0041729146391196 lketa = 2.58896043891468e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.235885950503162 lags = -7.38672925020819e-9
+ b0 = -2.1049625676525e-07 lb0 = 1.19540760102851e-12 pb0 = 3.85185988877447e-34
+ b1 = 5.54899964395e-10 lb1 = -1.11564005789709e-15
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.406770782793162+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 6.20403943312289e-7
+ nfactor = {1.9727581440482+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.79823267699225e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.396720728175106 lpclm = 3.18917515537414e-06 wpclm = 7.94093388050907e-23 ppclm = -3.53409685539013e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00124613070937175 lpdiblc2 = -3.26756945342507e-9
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 780185378.314556 lpscbe1 = 79.3324547245211
+ pscbe2 = 9.45624298832649e-09 lpscbe2 = 4.92833154399738e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.78791201328988e-10 lalpha0 = -6.30623738186469e-16
+ alpha1 = 2.00093291345109e-10 lalpha1 = -8.01119979017463e-16
+ beta0 = -17.6851374054458 lbeta0 = 0.000165558316861501 wbeta0 = -3.3881317890172e-21 pbeta0 = -1.29246970711411e-26
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.2473359332894e-09 lagidl = -8.59735973819656e-15
+ bgidl = 678067937.029324 lbgidl = 2576.65827615647
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.658393804945 lkt1 = 1.06276612150386e-6
+ kt2 = -0.0464346937487055 lkt2 = -4.84170320705919e-8
+ at = -42850.2895453823 lat = 0.422999606493931
+ ute = -2.1559858653625 lute = 7.1752335046354e-6
+ ua1 = -8.8739865677e-10 lua1 = 5.05314607869572e-15 wua1 = -3.94430452610506e-31
+ ub1 = 5.65421034524769e-19 lub1 = -5.68913621700037e-25
+ uc1 = 6.08383565119522e-11 luc1 = -4.21342569372177e-16 wuc1 = -1.23259516440783e-32 puc1 = 9.4039548065783e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.93 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.931424890001001+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.89352988908622e-7
+ k1 = 0.475366820955461 lk1 = -5.19661360002648e-8
+ k2 = 0.020580422653778 lk2 = -2.51732536497375e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 79659.8715761156 lvsat = -0.0949119803230556
+ ua = -1.07621574714662e-09 lua = 8.98190243076449e-16
+ ub = 3.11014895451446e-20 lub = 2.18135345183782e-24
+ uc = -7.89567475031345e-11 luc = 2.51213526557224e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00203856309834001 lu0 = 1.86041337261739e-8
+ a0 = 1.3342832198798 la0 = -3.45610319619412e-7
+ keta = 0.0266133366277374 lketa = -6.39558536606079e-8
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.103287510643325 lags = 1.3505732498662e-6
+ b0 = 2.369754010965e-07 lb0 = -5.96149442117293e-13 wb0 = 1.0097419586829e-28 pb0 = 1.92592994438724e-34
+ b1 = -4.428765550625e-09 lb1 = 1.88376260255505e-14 wb1 = 1.18329135783152e-30 pb1 = 6.01853107621011e-36
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.2141298027224+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -1.50879105749367e-7
+ nfactor = {1.45311295769765+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.30069731318361e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.15964838675 leta0 = -3.18890874427738e-7
+ etab = -0.13962972175 letab = 2.78778814751293e-7
+ dsub = 0.860559949999999 ldsub = -1.20336179029335e-6
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.499175844155821 lpclm = -3.97755515854073e-07 wpclm = -4.2351647362715e-22
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000571364515296475 lpdiblc2 = -5.65985774921502e-10
+ pdiblcb = -0.4253733 lpdiblcb = 8.022411935289e-7
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 9.63056774515734e-09 lpscbe2 = -2.05116627240852e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.8882357677209e-11 lalpha0 = -7.04660838659988e-17 palpha0 = -4.70197740328915e-38
+ alpha1 = 5.76486309697828e-16 lalpha1 = -2.17347769761512e-21 walpha1 = -4.70197740328915e-38 palpha1 = -4.48415508583941e-43
+ beta0 = 44.3702748108915 lbeta0 = -8.28949848576519e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.52426666601935e-10 lagidl = 1.01064897515416e-15
+ bgidl = 1643864125.94135 lbgidl = -1290.13179666484
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.29497272611779 lkt1 = -3.92274844692243e-7
+ kt2 = -0.0595567802632005 lkt2 = 4.12029873634653e-9
+ at = 85711.3304407276 lat = -0.0917267939779163
+ ute = 0.238846717647019 lute = -2.41303673743506e-06 pute = 8.07793566946316e-28
+ ua1 = 7.5900833711339e-10 lua1 = -1.538627934146e-15
+ ub1 = 3.30240300647921e-19 lub1 = 3.72687243486922e-25
+ uc1 = -1.35100873510396e-10 luc1 = 3.63145791862891e-16 wuc1 = -4.93038065763132e-32 puc1 = 9.4039548065783e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.94 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.061364804764+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 7.10119063191853e-8
+ k1 = 0.413766816430901 lk1 = 7.14638258657435e-8
+ k2 = 0.016148557298043 lk2 = -1.62929787848946e-08 wk2 = 1.32348898008484e-23
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -22098.3541553459 lvsat = 0.108984334596523
+ ua = 4.019367961654e-10 lua = -2.06363278699178e-15 pua = 7.52316384526264e-37
+ ub = 5.9654698090848e-19 lub = 1.04835166109189e-24
+ uc = -1.07948548475125e-10 luc = 8.32131809927318e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0163677609381 lu0 = -1.01077528488819e-8
+ a0 = 1.1019775132 la0 = 1.19868290943225e-7
+ keta = -0.0112258518738237 lketa = 1.18637770331905e-8
+ a1 = 0.0
+ a2 = 1.2014932 la2 = -8.04485174115601e-7
+ ags = 0.69017923456467 lags = -2.3932225190965e-7
+ b0 = -1.00359076911e-07 lb0 = 7.97787835041088e-14
+ b1 = 1.04101231542e-08 lb1 = -1.08955449556346e-14
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.26374281077549+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -5.14678842841256e-8
+ nfactor = {2.2796045020617+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.55371068479592e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.4908273035 leta0 = 9.84488731823965e-07 weta0 = 1.81152554149113e-22 peta0 = -1.60138763759865e-28
+ etab = 0.1646140785 letab = -3.3084452785504e-07 wetab = 3.0605682664462e-23 petab = -4.18096279767136e-29
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -0.0781728254105092 lpclm = 7.59097065862075e-7
+ pdiblc1 = 0.389489651956151 lpdiblc1 = 1.0226012169478e-9
+ pdiblc2 = 0.00014727096940705 lpdiblc2 = 2.83784458064153e-10
+ pdiblcb = 0.1757466 lpdiblcb = -4.022425870578e-07 wpdiblcb = 5.29395592033938e-23 ppdiblcb = -1.0097419586829e-28
+ drout = 0.230404054267382 ldrout = 6.60422273130658e-7
+ pscbe1 = 801208203.44943 lpscbe1 = -2.42091712233741
+ pscbe2 = 1.00507884655452e-08 lpscbe2 = -1.04712675196577e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -9.29295206703718e-11 lalpha0 = 1.93649726571034e-16 palpha0 = -3.52648305246686e-38
+ alpha1 = -1.00374318353055e-10 lalpha1 = 2.01122315683467e-16 walpha1 = -2.37431050956489e-33 palpha1 = 1.51937523604514e-38
+ beta0 = -1.94293465000289 lbeta0 = 9.90432127505426e-06 pbeta0 = -3.23117426778526e-27
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.288606493881e-11 lagidl = 5.59182419645833e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.462742255496781 lkt1 = -5.61095022810914e-8
+ kt2 = -0.0552726153526562 lkt2 = -4.46402387235358e-9
+ at = 6941.291585795 lat = 0.0661073322869943
+ ute = -1.75342231902647 lute = 1.57893847622583e-6
+ ua1 = -1.02473306547338e-09 lua1 = 2.03551357768339e-15 wua1 = -3.45126646034193e-31 pua1 = 6.23012005935812e-37
+ ub1 = 1.52278585337946e-18 lub1 = -2.0168556345245e-24
+ uc1 = 9.50456168403066e-11 luc1 = -9.80063256869943e-17 puc1 = 4.70197740328915e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.95 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.018366643504+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.78532329232015e-8
+ k1 = 0.432867755450021 lk1 = 5.22915830412653e-8
+ k2 = 0.0128144370961878 lk2 = -1.29464123123259e-08 wk2 = -9.30578189122156e-25 pk2 = 1.4791141972894e-31
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 83159.69948823 lvsat = 0.0033333526386955
+ ua = -1.50387380767641e-09 lua = -1.50707792165844e-16
+ ub = 1.4920864527798e-18 lub = 1.49469140372073e-25
+ uc = -3.709118344729e-11 luc = 1.20913054212477e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0071682521172 lu0 = -8.73902261553511e-10
+ a0 = 1.3394750152 la0 = -1.18515789231741e-7
+ keta = 0.0104579165941823 lketa = -9.90093694250654e-09 wketa = 2.48154183765908e-24 pketa = -3.94430452610506e-31
+ a1 = 0.0
+ a2 = -0.00298640000000017 la2 = 4.044907482312e-7
+ ags = 0.0671372126770802 lags = 3.86045585845646e-7
+ b0 = -1.0035658374e-08 lb0 = -1.08818123542899e-14
+ b1 = -3.60877335600001e-10 lb1 = -8.43363210062051e-17
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.31848029847242+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 3.47393845437744e-9
+ nfactor = {1.713364626012+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.12982581027399e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = -0.3312255933375 letab = 1.66846113477429e-7
+ dsub = 0.22207119204782 ldsub = 3.80703961922649e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.72584571993678 lpclm = -4.7922880714994e-8
+ pdiblc1 = 0.58629466742446 lpdiblc1 = -1.96517087374106e-7
+ pdiblc2 = -8.02528565176401e-05 lpdiblc2 = 5.12157630431021e-10
+ pdiblcb = -0.225
+ drout = 0.94174920473634 ldrout = -5.35783287850013e-8
+ pscbe1 = 797583593.101141 lpscbe1 = 1.21722389638217
+ pscbe2 = 1.70748966138426e-08 lpscbe2 = -8.09745589598078e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.78167108971381 lbeta0 = 1.14714658211119e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 9.33780278834562e-10 lagidl = -3.04925512350389e-16 wagidl = -7.88860905221012e-31
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.527955168835281 lkt1 = 9.34685086290166e-9
+ kt2 = -0.043721514196242 lkt2 = -1.60582452893845e-8
+ at = 79757.062028558 lat = -0.00698025942683167
+ ute = -0.269351715315134 lute = 8.93278369508384e-8
+ ua1 = 1.6991477649732e-09 lua1 = -6.98535499903246e-16
+ ub1 = -1.45731157578876e-18 lub1 = 9.74366498346799e-25 pub1 = -3.50324616081204e-46
+ uc1 = -2.97133802380454e-11 luc1 = 2.72183967274513e-17 puc1 = 1.17549435082229e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.96 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.964069663223999+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = 5.02052155815168e-10
+ k1 = 0.49245552604504 lk1 = 2.22752565961242e-8
+ k2 = -0.00877721848985161 lk2 = -2.06998286900348e-9
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 29991.62874372 lvsat = 0.0301158644190397
+ ua = -2.03670644350239e-09 lua = 1.17697589976695e-16
+ ub = 1.977239645256e-18 lub = -9.49185327335398e-26
+ uc = -2.64272507891217e-11 luc = 6.71953063155065e-18
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00535288544443999 lu0 = 4.0557838615906e-11
+ a0 = 1.40065148788 la0 = -1.49332397344255e-7
+ keta = -0.00841324462297796 lketa = -3.94910289102723e-10
+ a1 = 0.0
+ a2 = 1.08040210428168 la2 = -1.41247793196124e-7
+ ags = 1.25135733083852 lags = -2.1048516693617e-7
+ b0 = -6.3748418616e-08 lb0 = 1.61750775006935e-14
+ b1 = -1.0644885756e-09 lb1 = 2.70095879752715e-16
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.2306490710988+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -4.07695492042182e-8
+ nfactor = {1.7497916338892+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 1.94633095068393e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = 5.08399250000001e-05 letab = -2.8758079190025e-11 wetab = 6.46234853557053e-27 petab = 4.62223186652937e-33
+ dsub = -0.0376376544259198 ldsub = 1.68894312553022e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.624170992526718 lpclm = 3.29403474745765e-9
+ pdiblc1 = -0.0735726147024405 lpdiblc1 = 1.35879838253524e-7
+ pdiblc2 = -0.00934576645145274 lpdiblc2 = 5.17950259014845e-09 ppdiblc2 = 1.57772181044202e-30
+ pdiblcb = -0.225
+ drout = 1.24512186381992 ldrout = -2.0639714846315e-7
+ pscbe1 = 800072202.26248 lpscbe1 = -0.0363706622856625
+ pscbe2 = -7.33225872081081e-09 lpscbe2 = 4.19723368221019e-15 wpscbe2 = 1.57772181044202e-30 ppscbe2 = -1.50463276905253e-36
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.82126401216118 lbeta0 = 1.19736320508008e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 5.6030851539112e-10 lagidl = -1.16795460535735e-16 pagidl = 9.4039548065783e-38
+ bgidl = 718501708.2624 lbgidl = 141.799978991856
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.506690131559999 lkt1 = -1.36505015888661e-9
+ kt2 = -0.134474175456 lkt2 = 2.96568650249773e-8
+ at = 65234.204608 lat = 0.000335383110198373
+ ute = 0.00262240899999999 lute = -4.76745046127971e-8
+ ua1 = 2.2097447748e-10 lua1 = 4.60691647255671e-17
+ ub1 = 5.15527117359999e-19 lub1 = -1.94174550691046e-26
+ uc1 = 4.842226005912e-11 luc1 = -1.21411037663607e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.97 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.895472038957145+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.69034288422878e-8
+ k1 = -0.475192721214421 lk1 = 2.67799549318011e-7
+ k2 = 0.424510226624299 lk2 = -1.12009306180152e-07 pk2 = -1.89326617253043e-29
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 227262.218143858 lvsat = -0.0199381940412253
+ ua = 8.02797630049988e-10 lua = -6.02778297117974e-16
+ ub = -6.96694930414279e-19 lub = 5.83546908955008e-25
+ uc = 3.13756247644326e-15 luc = 1.32689039345937e-20
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.011653454326 lu0 = -1.55810440540895e-9
+ a0 = -0.470320092428565 la0 = 3.25394834642178e-7
+ keta = -0.194608099147397 lketa = 4.68488687339417e-08 wketa = -2.64697796016969e-23 pketa = 6.31088724176809e-30
+ a1 = 0.0
+ a2 = 0.143440229653004 la2 = 9.64903541390352e-8
+ ags = -1.75201096157885 lags = 5.51568480003768e-07 pags = 2.01948391736579e-28
+ b0 = -1.44631992842857e-07 lb0 = 3.66979094399966e-14
+ b1 = -3.57990626714285e-08 lb1 = 9.08340356880958e-15
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.25110826016186+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -3.55783777856814e-8
+ nfactor = {-2.04597080806712+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 1.1577432867533e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 1.45153429224443 leta0 = -2.43972980574055e-7
+ etab = 0.259331250696142 letab = -6.58167545453843e-08 wetab = 1.6130021944784e-23 petab = -1.55306990715387e-30
+ dsub = 1.59102145467072 ldsub = -2.44350249175394e-07 pdsub = -2.01948391736579e-28
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.666465439125862 lpclm = -7.4374620714814e-9
+ pdiblc1 = 1.23047101218629 lpdiblc1 = -1.94999063327833e-7
+ pdiblc2 = 0.0312405399469343 lpdiblc2 = -5.11858269123347e-9
+ pdiblcb = -0.815555173997886 lpdiblcb = 1.49843335964005e-7
+ drout = -1.060023465579 ldrout = 3.78494291401226e-7
+ pscbe1 = 799742134.776859 lpscbe1 = 0.047378351043335
+ pscbe2 = 3.07580668600386e-08 lpscbe2 = -5.46753889839547e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 11.69992923758 lbeta0 = -6.10676043133179e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.17521467858986e-08 lagidl = 3.0072807604264e-15 wagidl = 7.88860905221012e-31 pagidl = -1.88079096131566e-37
+ bgidl = 2005351041.92001 lbgidl = -184.716162985087
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.221955593000001 lkt1 = -7.36115988313306e-8
+ kt2 = 0.251204129485713 lkt2 = -6.82024483227987e-08 wkt2 = -5.29395592033938e-23 pkt2 = -6.31088724176809e-30
+ at = -8590.79699999955 lat = 0.019067222243201
+ ute = -0.324802089714287 lute = 3.54038957194747e-8
+ ua1 = 1.02463369042857e-09 lua1 = -1.57845698353513e-16
+ ub1 = 6.13178884000001e-19 lub1 = -4.41949307739721e-26
+ uc1 = -6.17595002111428e-11 luc1 = 1.58156448122939e-17 wuc1 = -2.00296714216273e-32 puc1 = -5.51012976947947e-40
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.98 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.229468383140045+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.39270278536531e-07 wvth0 = -2.85292705885803e-07 pvth0 = 5.24176847305155e-14
+ k1 = -4.36452513875971 lk1 = 9.82398262390859e-07 wk1 = 2.38503239762763e-06 pk1 = -4.38209157513317e-13
+ k2 = 1.57213907098805 lk2 = -3.22866596641639e-07 wk2 = -7.91420932464288e-07 pk2 = 1.45410142184461e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 570385.915453225 lvsat = -0.0829813403189675 wvsat = -0.186716498330198 pvsat = 3.43059823877023e-8
+ ua = 3.10525826997244e-09 lua = -1.02581629787285e-15 wua = -3.01185875964387e-15 pua = 5.53377845485646e-22
+ ub = -1.57657227983769e-18 lub = 7.45209413996619e-25 wub = 2.00152685793402e-24 pub = -3.67746534188791e-31
+ uc = 2.00978530096759e-13 luc = -2.30810105691901e-20 wuc = -3.18578627460677e-19 puc = 5.85334069592327e-26
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0211474467981396 lu0 = -3.30246412429258e-09 wu0 = -1.00475056957155e-08 pu0 = 1.84605836399091e-15
+ a0 = -11.0879002943758 la0 = 2.27619469788656e-06 wa0 = 9.13943514313035e-06 pa0 = -1.67921583715277e-12
+ keta = -0.45033468060373 lketa = 9.38342807246583e-08 wketa = 5.50351904464447e-07 pketa = -1.01117806462966e-13
+ a1 = 0.0
+ a2 = -7.62025840628531 la2 = 1.52293799561589e-06 wa2 = 4.42030870023431e-06 pa2 = -8.12156578420152e-13
+ ags = 21.9054591209721 lags = -3.79508947067358e-06 wags = -1.38480849004834e-05 pags = 2.54435018302052e-12
+ b0 = -5.1915219842844e-06 lb0 = 9.63978148237526e-13 wb0 = 2.06148131062557e-12 pb0 = -3.78762145645168e-19
+ b1 = 3.22713135398827e-07 lb1 = -5.67871181192327e-14 wb1 = -1.70229522371079e-13 pb1 = 3.12767808338054e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.590138983148677+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 2.67127540408558e-08 wvoff = 1.07776432024766e-07 pvoff = -1.98020871852065e-14
+ nfactor = {-17.4790490535123+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 3.99330905202369e-06 wnfactor = 1.14750770719366e-05 pnfactor = -2.10835033565813e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -6.59726337903448 leta0 = 1.23485676196303e-06 weta0 = 3.73455818304312e-06 peta0 = -6.86161578645063e-13
+ etab = -1.34283219696216 letab = 2.28553542183219e-07 wetab = 4.94240831085623e-07 petab = -9.08083506178548e-14
+ dsub = 0.0836561835830043 ldsub = 3.26024941773637e-08 wdsub = 1.06269981956951e-07 pdsub = -1.95253025948966e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 15.7408700676124 lpclm = -2.7771030476772e-06 wpclm = -8.74797482033118e-06 ppclm = 1.60729165766391e-12
+ pdiblc1 = 6.54285626830813 lpdiblc1 = -1.17105954359087e-06 wpdiblc1 = -3.72549156489708e-06 ppdiblc1 = 6.84495741693236e-13
+ pdiblc2 = 0.132618981059993 lpdiblc2 = -2.37451478122592e-08 wpdiblc2 = -7.57652432826798e-08 ppdiblc2 = 1.39205754440566e-14
+ pdiblcb = -2.24374062827912 lpdiblcb = 4.1224813403546e-07 wpdiblcb = 1.52539770444004e-06 ppdiblcb = -2.80265896429882e-13
+ drout = 1.0
+ pscbe1 = 801248644.322891 lpscbe1 = -0.229417167377505 wpscbe1 = -0.724753371352563 ppscbe1 = 1.33161111178903e-7
+ pscbe2 = -2.80519894884281e-08 lpscbe2 = 5.33780918467735e-15 wpscbe2 = -8.12755845985368e-15 ppscbe2 = 1.4933006985043e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 13.4564961327463 lbeta0 = -9.33415348482759e-07 wbeta0 = -1.11655225213051e-06 pbeta0 = 2.05147494940691e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 1.24941972774721e-08 lagidl = -1.44757277336887e-15 wagidl = 4.65344841053808e-15 pagidl = -8.54992036813395e-22
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = 2.05119983359304 lkt1 = -4.91265264825549e-07 wkt1 = -1.49315590630972e-06 pkt1 = 2.74342014134005e-13
+ kt2 = -0.12
+ at = 925604.553668076 lat = -0.152575292121097 wat = -0.373344368917033 pat = 6.85956809342333e-8
+ ute = 6.12162148113926 lute = -1.14901684622416e-06 wute = -4.02281327125083e-06 pute = 7.3912355076673e-13
+ ua1 = -6.56909877244079e-10 lua1 = 1.51109345965687e-16 wua1 = 5.20023284182953e-16 pua1 = -9.55454380727867e-23
+ ub1 = 5.150259163673e-19 lub1 = -2.61609915719125e-26 wub1 = -8.26453706860854e-26 pub1 = 1.51846818922666e-32
+ uc1 = 6.58841669432414e-10 luc1 = -1.16582569889826e-16 wuc1 = -3.69201021914809e-16 puc1 = 6.78344113594736e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.99 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.12883844905462+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} wvth0 = 6.03446041026588e-8
+ k1 = 0.5505891619672 wk1 = -4.17465481531883e-8
+ k2 = -0.0742247222643192 wk2 = 4.08651303963909e-8
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -237702.895675431 wvsat = 0.152185791302105
+ ua = -1.2810064494546e-09 wua = 2.13965046611464e-16
+ ub = 3.64759366001001e-18 wub = -1.37689372503153e-24
+ uc = -7.46639522531846e-12 wuc = -3.51411976816733e-17
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0194897825025418 wu0 = -5.44614843515361e-9
+ a0 = 0.0592326835903076 wa0 = 6.91700539875733e-7
+ keta = -0.0524925631670172 wketa = 3.47679868538975e-8
+ a1 = 0.0
+ a2 = 0.108759816153846 wa2 = 4.01218060638227e-7
+ ags = 0.577783938340492 wags = -1.98984288229748e-7
+ b0 = -8.69913434169231e-08 wb0 = 1.50049521324402e-14
+ b1 = 3.57820029769231e-10 wb1 = 3.34851163389797e-17
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.378124576999246+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} wvoff = 2.83646286597299e-8
+ nfactor = {3.27957060511+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} wnfactor = -8.15068959611788e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.00728266104669468 wpclm = -3.21700289187961e-9
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00462803992120334 wpdiblc2 = 3.17259304013985e-9
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 1292305062.90435 wpscbe1 = -291.49755087533
+ pscbe2 = 8.19597902642107e-09 wpscbe2 = 7.67238135653037e-16
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.46486307692308e-10 walpha0 = -2.01111809843723e-16
+ alpha1 = 4.46486307692308e-10 walpha1 = -2.01111809843723e-16
+ beta0 = -90.551303076923 wbeta0 = 5.43001886578052e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.28415214603898e-09 wagidl = -1.22528363639629e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.17385123306154 wkt1 = 3.76260085036621e-7
+ kt2 = -0.0300782446267031 wkt2 = -1.30050218839845e-8
+ at = -249995.0962425 wat = 0.150909525701246
+ ute = -4.58147212363077 wute = 1.92817958805768e-6
+ ua1 = -3.28960529262205e-09 wua1 = 1.76077317231826e-15
+ ub1 = 1.35807361061972e-18 wub1 = -5.01338799825949e-25
+ uc1 = -2.03106574174729e-10 wuc1 = 1.22646295604921e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.100 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.10948925172375+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.87056177170956e-07 wvth0 = 4.91137069276693e-08 pvth0 = 2.24659868438929e-13
+ k1 = 0.574355740814426 lk1 = -4.75420297583363e-07 wk1 = -5.55414357999574e-08 pk1 = 2.75949249250966e-13
+ k2 = -0.0670095009372213 lk2 = -1.44331360963172e-07 wk2 = 3.66771836080165e-08 pk2 = 8.37745693728481e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -327296.44819703 lvsat = 1.79220550316356 wvsat = 0.204188774098032 pvsat = -1.04025378305333e-6
+ ua = -1.24500116300283e-09 lua = -7.20240136769779e-16 wua = 1.93066418984632e-16 pua = 4.18050567113583e-22
+ ub = 3.56520234338192e-18 lub = 1.64813389934676e-24 wub = -1.3290711518602e-24 pub = -9.56629985092422e-31
+ uc = 3.14482087977308e-12 luc = -2.12263933771552e-16 wuc = -4.1300289190227e-17 puc = 1.23204822059676e-22
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0194849088629452 lu0 = 9.74909852300865e-11 wu0 = -5.4433196178005e-09 pu0 = -5.65869070372145e-17
+ a0 = -0.697713175798624 la0 = 1.51417428666717e-05 wa0 = 1.13105629032174e-06 pa0 = -8.78875512393658e-12
+ keta = -0.0863636558239739 lketa = 6.77548293928021e-07 wketa = 5.44278596811787e-08 pketa = -3.93270846850888e-13
+ a1 = 0.0
+ a2 = -0.352282006377447 la2 = 9.22255751974938e-06 wa2 = 6.68821579982076e-07 pa2 = -5.35306935081468e-12
+ ags = 0.783913218218862 lags = -4.12335507816919e-06 wags = -3.18628359633966e-07 pags = 2.39332805940291e-12
+ b0 = 2.73404702607802e-07 lb0 = -7.20926627893431e-12 wb0 = -1.94180517732992e-13 pb0 = 4.18449028666766e-18
+ b1 = -1.58641297923116e-09 lb1 = 3.88919180018303e-14 wb1 = 1.16198055906569e-15 pb1 = -2.2574121528022e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.269132556912914+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -2.18024726893762e-06 wvoff = -3.48978493414242e-08 pvoff = 1.26548571885346e-12
+ nfactor = {3.44516134415316+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.31243293109206e-06 wnfactor = -9.11183156574235e-07 pnfactor = 1.92264273354621e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.55493289552115e-06 lcit = 2.31141792474922e-10 wcit = 6.7068551213997e-12 pcit = -1.34162139118162e-16
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.42345057948295 lpclm = -2.83286449235647e-05 wpclm = -8.25206463359257e-07 ppclm = 1.64428576960035e-11
+ pdiblc1 = 0.39
+ pdiblc2 = -0.00905765647069958 lpdiblc2 = 8.86088667485042e-08 wpdiblc2 = 5.74368511912036e-09 ppdiblc2 = -5.14314394663411e-14
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 1621356134.90286 lpscbe1 = -6582.24978762193 wpscbe1 = -482.489388507783 ppscbe1 = 0.00382054972517893
+ pscbe2 = 7.2406543815033e-09 lpscbe2 = 1.91100591252547e-14 wpscbe2 = 1.32173932101688e-15 ppscbe2 = -1.10920936602017e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 6.7758496560273e-10 lalpha0 = -4.62283584949844e-15 walpha0 = -3.35248912271717e-16 palpha0 = 2.68324278236325e-21
+ alpha1 = 6.7758496560273e-10 lalpha1 = -4.62283584949844e-15 walpha1 = -3.35248912271717e-16 palpha1 = 2.68324278236325e-21
+ beta0 = -148.728845080245 lbeta0 = 0.00116376801683074 wbeta0 = 8.80683073533859e-05 pbeta0 = -6.75488430298704e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 3.9323543701791e-09 lagidl = -1.29664642217051e-14 wagidl = -1.60152107939883e-15 pagidl = 7.5261533544256e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.28940056201675 lkt1 = 2.31141792474922e-06 wkt1 = 4.43328636250618e-07 pkt1 = -1.34162139118162e-12
+ kt2 = -0.0300782446267031 wkt2 = -1.30050218839845e-8
+ at = -249995.0962425 wat = 0.150909525701246
+ ute = -4.58147212363077 wute = 1.92817958805768e-6
+ ua1 = -3.28960529262205e-09 wua1 = 1.76077317231826e-15
+ ub1 = 1.35807361061972e-18 wub1 = -5.01338799825949e-25
+ uc1 = -2.18821282912638e-10 luc1 = 3.14352837765893e-16 wuc1 = 1.31767618570025e-16 puc1 = -1.824605092007e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.101 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.56202772763697+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.23494095626538e-06 wvth0 = 2.84967050756747e-07 pvth0 = -1.6630473227262e-12
+ k1 = 0.587705247905173 lk1 = -5.82266188019308e-07 wk1 = -5.38325070793442e-08 pk1 = 2.62271440055149e-13
+ k2 = -0.233856373756235 lk2 = 1.19106646096517e-06 wk2 = 1.22997276911365e-07 pk2 = -6.07108409962244e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -313363.519912931 lvsat = 1.68069006526947 wvsat = 0.177822484051951 pvsat = -8.2922503732394e-7
+ ua = -1.59757532470955e-09 lua = 2.1016693162297e-15 wua = 3.62563859498663e-16 pua = -9.38561690944112e-22
+ ub = 8.75656396131913e-18 lub = -3.99021383970707e-23 wub = -3.93592773514777e-24 pub = 1.99079540768336e-29
+ uc = -2.49330149931198e-12 luc = -1.67137907628029e-16 wuc = -3.53130171731087e-17 puc = 7.52842954362898e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0447887324855724 lu0 = -2.02427557169371e-07 wu0 = -1.81426114578996e-08 pu0 = 1.01585154270195e-13
+ a0 = 1.20739760524257 la0 = -1.06255160203468e-07 wa0 = 2.69944894710161e-08 pa0 = 4.78607455718019e-14
+ keta = -0.0161520739015416 lketa = 1.15593538713247e-07 wketa = 1.17972778136307e-08 pketa = -5.2067051948393e-14
+ a1 = 0.0
+ a2 = 0.8
+ ags = 0.272854897872505 lags = -3.29807346884838e-08 wags = -2.1457967453272e-08 pags = 1.48555848833495e-14
+ b0 = -1.90318281700636e-06 lb0 = 1.02115590791897e-11 wb0 = 9.82489784071182e-13 pb0 = -5.23326463800237e-18
+ b1 = 6.02145650419034e-09 lb1 = -2.19994380423233e-14 wb1 = -3.1729654388178e-15 pb1 = 1.2121628808456e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.07924646955952+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 4.30368818747113e-06 wvoff = 3.90326542316307e-07 pvoff = -2.13789677706245e-12
+ nfactor = {5.47057060858602+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.95232678993391e-05 wnfactor = -2.03024298397911e-06 pnfactor = 1.08792988031209e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.73243153846154e-05 wcit = -1.00555904921862e-11
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -3.89505208928862 lpclm = 1.42392303970704e-05 wpclm = 2.03054416826011e-06 ppclm = -6.4138078740593e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0038360916031534 lpdiblc2 = -1.45892502038793e-08 wpdiblc2 = -1.50329669949165e-09 ppdiblc2 = 6.57146806568382e-15
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 754703244.867284 lpscbe1 = 354.208547901191 wpscbe1 = 14.7906507774946 ppscbe1 = -0.000159546935489937
+ pscbe2 = 9.35337185609816e-09 lpscbe2 = 2.20043255416315e-15 wpscbe2 = 5.97097175957701e-17 ppscbe2 = -9.91145676323329e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.51791925600213e-10 lalpha0 = -2.81564864405997e-15 walpha0 = -1.5845841099034e-16 palpha0 = 1.26825881317095e-21
+ alpha1 = 5.4690284077448e-10 lalpha1 = -3.57689101450046e-15 walpha1 = -2.01299429756299e-16 palpha1 = 1.61114688882167e-21
+ beta0 = -95.6819979654929 lbeta0 = 0.000739195216032445 wbeta0 = 4.52718893679614e-05 pbeta0 = -3.32957327386969e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 7.10831861491262e-09 lagidl = -3.83860340540989e-14 wagidl = -2.82147087205647e-15 pagidl = 1.72903057682627e-20
+ bgidl = -437382581.235441 lbgidl = 11504.4263990593 wbgidl = 647.443398307559 pbgidl = -0.00518196409266635
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.65336777816859 lkt1 = 5.22451434358185e-06 wkt1 = 5.77514932220911e-07 pkt1 = -2.41561267638682e-12
+ kt2 = 0.0096260958744111 lkt2 = -3.17782940312004e-07 wkt2 = -3.25394874546827e-08 pkt2 = 1.56348646725561e-13
+ at = -559663.624232063 lat = 2.47850421653149 wat = 0.299975100841526 pat = -1.19308106291424e-6
+ ute = -9.79917174687212 lute = 4.17610746586244e-05 wute = 4.43635119621357e-06 pute = -2.00747358698604e-11
+ ua1 = -8.35599421874064e-09 lua1 = 4.055002423881e-14 wua1 = 4.33501335294486e-15 pua1 = -2.06035310836071e-20
+ ub1 = 3.32225859310738e-18 lub1 = -1.57208121624409e-23 wub1 = -1.60015728917074e-24 pub1 = 8.79464980417902e-30
+ uc1 = -8.85824387890296e-12 luc1 = -1.3661352665287e-15 wuc1 = 4.04541510973848e-17 puc1 = 5.48388103754494e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.102 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.525874946198378+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -9.13538127822098e-07 wvth0 = -2.35394246091233e-07 pvth0 = 4.20340373386851e-13
+ k1 = 0.422937600406743 lk1 = 7.74194796025288e-08 wk1 = 3.04316078273773e-08 pk1 = -7.50995775126844e-14
+ k2 = 0.123682702727529 lk2 = -2.40424538342397e-07 wk2 = -5.98438832482234e-08 pk2 = 1.24938776726987e-13
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 239998.020429625 lvsat = -0.534821794730849 wvsat = -0.0930654244829703 pvsat = 2.55337821378307e-7
+ ua = -1.86483270458357e-09 lua = 3.17169650752481e-15 wua = 4.5773867556243e-16 pua = -1.31961624278754e-21
+ ub = -3.36606649111377e-18 lub = 8.63363719213989e-24 wub = 1.97182568478341e-24 pub = -3.74511324640776e-30
+ uc = -5.49169724396132e-11 luc = 4.27524736967956e-17 wuc = -1.39534595276247e-17 puc = -1.02336703743364e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.0226468674732244 lu0 = 6.75665797604624e-08 wu0 = 1.43282187746004e-08 pu0 = -2.84193802690633e-14
+ a0 = 1.53979596918711 la0 = -1.43708945907424e-06 wa0 = -1.19286217208493e-07 pa0 = 6.33529638167875e-13
+ keta = 0.0570820188382189 lketa = -1.77616215113992e-07 wketa = -1.76850042465306e-08 pketa = 6.5972133651183e-14
+ a1 = 0.0
+ a2 = 0.8
+ ags = -0.747028384632029 lags = 4.05035961962324e-06 wags = 3.73647931719186e-07 pags = -1.56704294212809e-12
+ b0 = 1.36437424057204e-06 lb0 = -2.87086694161983e-12 wb0 = -6.54378588674234e-13 pb0 = 1.32031928261475e-18
+ b1 = -4.29912760458287e-09 lb1 = 1.93214251332476e-14 wb1 = -7.52460382247197e-17 pb1 = -2.80812580438687e-22
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.193789056491329+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -7.93206158351014e-07 wvoff = -2.36769240874915e-07 pvoff = 3.72827304261089e-13
+ nfactor = {-0.770757436219466+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.46534315747413e-06 wnfactor = 1.29080598525618e-06 pnfactor = -2.4172945496224e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.73243153846154e-05 wcit = -1.00555904921862e-11
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.15964838675 leta0 = -3.18890874427738e-7
+ etab = -0.13962972175 letab = 2.78778814751293e-7
+ dsub = 0.860559950000001 ldsub = -1.20336179029335e-6
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.0466107679763708 lpclm = -1.54213525943571e-06 wpclm = 2.62683342810006e-07 ppclm = 6.64234852202528e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00351522544686283 lpdiblc2 = -1.33045877853556e-08 wpdiblc2 = -1.70871167700311e-09 ppdiblc2 = 7.3938947898407e-15
+ pdiblcb = -1.11963934877123 lpdiblcb = 3.58189708377389e-06 wpdiblcb = 4.02974370073593e-07 ppdiblcb = -1.61340178361786e-12
+ drout = 0.56
+ pscbe1 = 886426217.291707 lpscbe1 = -173.175063652565 wpscbe1 = -50.1645594403035 ppscbe1 = 0.000100516383180997
+ pscbe2 = 1.00121335432869e-08 lpscbe2 = -4.37073351970058e-16 wpscbe2 = -2.21473075653097e-16 ppscbe2 = 1.34635152039333e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -5.20014928941236e-10 lalpha0 = 1.07520652909383e-15 walpha0 = 3.24401981645975e-16 palpha0 = -6.64985275220022e-22
+ alpha1 = -6.93616758145484e-10 lalpha1 = 1.38981824084217e-15 walpha1 = 4.02597835498468e-16 palpha1 = -8.06696520688593e-22
+ beta0 = 268.77533872015 lbeta0 = -0.000719994649947975 wbeta0 = -0.000130251924935992 pbeta0 = 3.69793160227639e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -4.07676848178068e-09 lagidl = 6.3960682628063e-15 wagidl = 2.2778143533362e-15 pagidl = -3.12587076505436e-21
+ bgidl = 3874765162.47088 lbgidl = -5760.26182329327 wbgidl = -1294.88679661512 pbgidl = 0.002594607405642
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.0845683999151641 lkt1 = -1.05653949751088e-06 wkt1 = -1.22125445947308e-07 pkt1 = 3.85560593817758e-13
+ kt2 = -0.0743404198762172 lkt2 = 1.83965696938064e-08 wkt2 = 8.58090046459047e-09 pkt2 = -8.28640735963452e-15
+ at = 197722.662773724 lat = -0.55386825450105 wat = -0.0650149840509721 pat = 2.68241784642656e-7
+ ute = 2.75729991293048 lute = -8.51168528929205e-06 wute = -1.46179132873541e-06 pute = 3.53985199598117e-12
+ ua1 = 3.48789929041716e-09 lua1 = -6.86976305229092e-15 wua1 = -1.5839361795862e-15 pua1 = 3.09436248512212e-21
+ ub1 = -1.01989151408656e-18 lub1 = 1.663997512685e-24 wub1 = 7.83659979516324e-25 pub1 = -7.4951806043323e-31
+ uc1 = -7.55044741369449e-10 luc1 = 1.62139623762862e-15 wuc1 = 3.59835383097939e-16 puc1 = -7.3032907438678e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.103 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.06928117724539+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.75302869732423e-07 wvth0 = 4.59491749538977e-09 pvth0 = -6.05338333340657e-14
+ k1 = 0.299818508810862 lk1 = 3.24117266363217e-07 wk1 = 6.61392668781756e-08 pk1 = -1.46648192305518e-13
+ k2 = 0.0449703132017618 lk2 = -8.27059259407634e-08 wk2 = -1.67290751870585e-08 pk2 = 3.85482130261647e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -270799.679102602 lvsat = 0.488680412145961 wvsat = 0.144354257182051 pvsat = -2.20387829623391e-7
+ ua = 2.69782732993461e-09 lua = -5.97065597142042e-15 wua = -1.33260879347484e-15 pua = 2.26776206238892e-21
+ ub = -6.09102342914811e-19 lub = 3.10941714857674e-24 wub = 6.99797689455266e-25 pub = -1.19630877524491e-30
+ uc = -1.09813714348657e-10 luc = 1.5275088705243e-16 wuc = 1.08260233133935e-18 puc = -4.03619237111843e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.0245015227487024 lu0 = -2.69062056240897e-08 wu0 = -4.72109726200391e-09 pu0 = 9.75036290090995e-15
+ a0 = -0.599729273655665 la0 = 2.84994787434285e-06 wa0 = 9.87725414049565e-07 pa0 = -1.58462609876773e-12
+ keta = -0.0934386501621791 lketa = 1.23987016544182e-07 wketa = 4.77189553786664e-08 pketa = -6.50799385804919e-14
+ a1 = 0.0
+ a2 = 2.59261216431569 la2 = -3.59191614984077e-06 wa2 = -8.07450240919478e-07 pa2 = 1.61791469358831e-12
+ ags = 2.73907773928819 lags = -2.93486626237779e-06 wags = -1.18924666667338e-06 pags = 1.56458054019284e-12
+ b0 = -1.36669311658798e-07 lb0 = 1.36823558422324e-13 wb0 = 2.10756294371806e-14 pb0 = -3.31106242042848e-20
+ b1 = -4.18341012226084e-10 lb1 = 1.15453649721848e-14 wb1 = 6.28518927873986e-15 pb1 = -1.30254267194061e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.199409588222231+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -5.34105838317848e-09 wvoff = -3.7341073899678e-08 pvoff = -2.67734950367036e-14
+ nfactor = {2.51966398386984+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.12778282586567e-06 wnfactor = -1.39338253156758e-07 pnfactor = 4.48332655645464e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.73243153846154e-05 wcit = -1.00555904921862e-11
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -0.490827303499999 leta0 = 9.84488731823965e-07 weta0 = -4.4254162771587e-23 peta0 = -9.62410304369634e-29
+ etab = -0.122304207890111 letab = 2.44063110888277e-07 wetab = 1.66536612189642e-07 petab = -3.33694905552588e-13
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.29025759379565 lpclm = 3.14032499370281e-06 wpclm = 1.28396522870028e-06 ppclm = -1.38214136485804e-12
+ pdiblc1 = 0.375960985250206 lpdiblc1 = 2.81304371416497e-08 wpdiblc1 = 7.85247377919792e-09 ppdiblc1 = -1.57342608430137e-14
+ pdiblc2 = -0.00669261974503682 lpdiblc2 = 7.14920848454504e-09 wpdiblc2 = 3.97009281514423e-09 ppdiblc2 = -3.98491317162316e-15
+ pdiblcb = 1.56427869754246 lpdiblcb = -1.79595807492039e-06 wpdiblcb = -8.05948740147185e-07 ppdiblcb = 8.08957346794154e-13
+ drout = -0.28031738154589 ldrout = 1.68377166787709e-06 wdrout = 2.96439166576256e-07 pdrout = -5.93984940561341e-13
+ pscbe1 = 723307141.234561 lpscbe1 = 153.672011972651 wpscbe1 = 45.2162849237138 ppscbe1 = -9.06013622390474e-5
+ pscbe2 = 1.07196033089474e-08 lpscbe2 = -1.85465386792629e-15 wpscbe2 = -3.88201670948611e-16 ppscbe2 = 4.6871474047662e-22
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.71378445183803e-11 lalpha0 = 1.67761770091967e-16 walpha0 = -1.4970319330588e-17 palpha0 = 1.50262035326491e-23
+ alpha1 = -1.00377846806954e-10 lalpha1 = 2.01125857309084e-16 walpha1 = 2.04802825915812e-21 palpha1 = -2.05567354864956e-27
+ beta0 = -194.855803547109 lbeta0 = 0.000208998369640627 wbeta0 = 0.000111972840902259 pbeta0 = -1.15560596499736e-10
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 4.90202955629876e-10 lagidl = -2.75492311639068e-15 wagidl = -2.42224160960975e-16 pagidl = 1.92361356731385e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.60675497261295 lkt1 = -1.02170296394287e-08 wkt1 = 8.3589618223716e-08 pkt1 = -2.66374688588396e-14
+ kt2 = -0.0813584684536592 lkt2 = 3.24588652240297e-08 wkt2 = 1.5141069104292e-08 pkt2 = -2.14312337485697e-14
+ at = -275740.891632723 lat = 0.394826293760443 wat = 0.164077841506328 pat = -1.90799069989749e-7
+ ute = -4.71174433763247 lute = 6.4542851540212e-06 wute = 1.71710535756792e-06 pute = -2.82980819795546e-12
+ ua1 = -4.81737567659755e-09 lua1 = 9.77179047319037e-15 wua1 = 2.20137189458855e-15 pua1 = -4.49038421826829e-21
+ ub1 = 4.66382505497671e-18 lub1 = -9.72465293939386e-24 wub1 = -1.82316029406934e-24 pub1 = 4.47385374681939e-30
+ uc1 = 2.16356236445235e-10 luc1 = -3.25031957850934e-16 wuc1 = -7.04125898206517e-17 puc1 = 1.31772987133306e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.104 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.881378171726709+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.33015777058567e-08 wvth0 = -7.95125200483304e-08 pvth0 = 2.38875772740068e-14
+ k1 = 0.622458808473364 lk1 = 2.72550462075082e-10 wk1 = -1.10044752006656e-07 pk1 = 3.01935215218109e-14
+ k2 = -0.0415441063801841 lk2 = 4.13145196948195e-09 wk2 = 3.15514489787862e-08 pk2 = -9.91254233639113e-15
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 301738.72991216 lvsat = -0.0859952827496531 wvsat = -0.126870307502828 pvsat = 5.1849216361457e-8
+ ua = -4.12867780064813e-09 lua = 8.81332502814796e-16 wua = 1.52352075620937e-15 pua = -5.99029418904262e-22
+ ub = 2.97129458894317e-18 lub = -4.84345405027861e-25 wub = -8.58580032731202e-25 pub = 3.67886370978483e-31
+ uc = 6.65176850621943e-11 luc = -2.4238757472422e-17 wuc = -6.01379234884707e-17 puc = 2.10871383315111e-23
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.00625117325150133 lu0 = 3.96129019028279e-09 wu0 = 7.78906658949114e-09 pu0 = -2.80650139224273e-15
+ a0 = 3.80991448227088 la0 = -1.57615708172457e-06 wa0 = -1.43392261483878e-06 pa0 = 8.46061942212456e-13
+ keta = -0.0135478117091812 lketa = 4.37979455912393e-08 wketa = 1.39336976917236e-08 pketa = -3.11685605266037e-14
+ a1 = 0.0
+ a2 = -2.78522432863138 la2 = 1.80599580673447e-06 wa2 = 1.61490048183896e-06 pa2 = -8.13478664418184e-13
+ ags = 0.208204726885906 lags = -3.94545501020205e-07 wags = -8.18801276207598e-08 pags = 4.53080201849937e-13
+ b0 = 9.78806855898077e-08 lb0 = -9.86020139660098e-14 wb0 = -6.26381209428696e-14 pb0 = 5.09156296059341e-20
+ b1 = 3.92510449523064e-08 lb1 = -2.82721068101533e-14 wb1 = -2.29920351997986e-14 pb1 = 1.63610896381107e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.294954741440977+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = 9.0560764892533e-08 wvoff = -1.36549908239862e-08 pvoff = -5.05479982605169e-14
+ nfactor = {1.71982162248329+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.2495465294406e-07 wnfactor = -3.74784866721928e-09 pnfactor = 3.12236092175968e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 4.47779741078923e-05 lcit = -1.75188132312909e-11 wcit = -2.0186256022987e-11 pcit = 1.01684833052273e-17
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = 0.242621887979425 letab = -1.22225254097141e-07 wetab = -3.33079556045242e-07 petab = 1.67786329838316e-13
+ dsub = 0.359016089122396 ldsub = -9.93857161830895e-08 wdsub = -7.94872278877695e-08 pdsub = 7.97839537094744e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.13587742734056 lpclm = -2.98599789467295e-07 wpclm = -2.37995605998134e-07 ppclm = 1.45500949636297e-13
+ pdiblc1 = 1.1541126351864 lpdiblc1 = -7.52926052903759e-07 wpdiblc1 = -3.29579832227593e-07 ppdiblc1 = 3.22957679962101e-13
+ pdiblc2 = 0.00304289178008881 lpdiblc2 = -2.62264570510388e-09 wpdiblc2 = -1.81277371234368e-09 ppdiblc2 = 1.81954079661186e-15
+ pdiblcb = 0.473146348931077 lpdiblcb = -7.00752529251637e-07 wpdiblcb = -4.05226621232033e-07 ppdiblcb = 4.06739332209092e-13
+ drout = 2.0438083268447 ldrout = -6.49030001782921e-07 wdrout = -6.39670600775425e-07 pdrout = 3.45619324551863e-13
+ pscbe1 = 953385717.53088 lpscbe1 = -77.2654476489829 wpscbe1 = -90.4325698474272 ppscbe1 = 4.55538697069541e-5
+ pscbe2 = 4.5742548364341e-08 lpscbe2 = -3.70083395772117e-14 wpscbe2 = -1.66396281743756e-14 ppscbe2 = 1.67808078190409e-20
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 18.5556099011584 lbeta0 = -5.20970861404288e-06 wbeta0 = -6.83397320699219e-06 pbeta0 = 3.68972344658515e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -3.68749353895651e-09 lagidl = 1.43836871921e-15 wagidl = 2.68233612886287e-15 pagidl = -1.01186410607191e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.725270856730285 lkt1 = 1.08741274273316e-07 wkt1 = 1.14528378819411e-07 pkt1 = -5.76917238478383e-14
+ kt2 = -0.0987730019545587 lkt2 = 4.9938407178488e-08 wkt2 = 3.19536561528327e-08 pkt2 = -3.83065821845626e-14
+ at = 124204.462139948 lat = -0.00661205601786169 wat = -0.0257987022309343 pat = -2.13717114715959e-10
+ ute = 3.3633267884672 lute = -1.6509302125922e-06 wute = -2.10852357584309e-06 pute = 1.01010180826397e-12
+ ua1 = 9.84165260362252e-09 lua1 = -4.94195995959976e-15 wua1 = -4.72617199700787e-15 pua1 = 2.46302019467546e-21
+ ub1 = -1.06180622085862e-17 lub1 = 5.61428160932397e-24 wub1 = 5.31719464344604e-24 pub1 = -2.69315613567772e-30
+ uc1 = -2.40237700270098e-10 luc1 = 1.33266444030158e-16 wuc1 = 1.22195094229709e-16 puc1 = -6.15537014016138e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.105 pmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.852666450325067+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -2.77646192626696e-08 wvth0 = -6.46620119499948e-08 pvth0 = 1.64068862781082e-14
+ k1 = 0.666392475378712 lk1 = -2.18582873691568e-08 wk1 = -1.00958606163032e-07 pk1 = 2.56165300175646e-14
+ k2 = -0.0499945300865534 lk2 = 8.38820925436245e-09 wk2 = 2.39238548481591e-08 pk2 = -6.07027146218796e-15
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 113098.970120475 lvsat = 0.00902878936949142 wvsat = -0.0482381769914611 pvsat = 1.22396173625744e-8
+ ua = -3.19734682274636e-09 lua = 4.12190355323402e-16 wua = 6.73673048733405e-16 pua = -1.70933083674273e-22
+ ub = 2.42248527187219e-18 lub = -2.07892041311746e-25 wub = -2.58434898597213e-25 pub = 6.55734621257669e-32
+ uc = 3.70173222797515e-11 luc = -9.37845122693377e-18 wuc = -3.68252731244269e-17 puc = 9.3437870256802e-24
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = -0.00234557434522299 lu0 = 1.99391113642646e-09 wu0 = 4.46843395232563e-09 pu0 = -1.13378915202544e-15
+ a0 = 0.547853854172759 la0 = 6.70505046491832e-08 wa0 = 4.94991206687488e-07 pa0 = -1.25595603846436e-13
+ keta = 0.158012375370252 lketa = -4.2622582126845e-08 wketa = -9.65987887490347e-08 pketa = 2.45103004656588e-14
+ a1 = 0.0
+ a2 = 1.08040210428168 la2 = -1.41247793196124e-7
+ ags = -1.58676556808507 lags = 5.09640270576409e-07 wags = 1.6473379180926e-06 pags = -4.17983991971389e-13
+ b0 = -1.97185130287197e-07 lb0 = 5.00323746631613e-14 wb0 = 7.74509641160783e-14 pb0 = -1.96518654780649e-20
+ b1 = -3.40002407327725e-08 lb1 = 8.62698308184855e-15 wb1 = 1.91169710832424e-14 pb1 = -4.85060642386433e-21
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0.165100632334302+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -1.4118430870541e-07 wvoff = -2.29705871013023e-07 pvoff = 5.82839597697474e-14
+ nfactor = {-0.388946893182752+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 7.37301637757938e-07 wnfactor = 1.24139270849313e-06 pnfactor = -3.14982296104088e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 0.49
+ etab = 2.90228515959039e-05 letab = -2.32223677039835e-11 wetab = 1.2663331913501e-11 petab = -3.21310519640836e-18
+ dsub = -0.311527448575071 ldsub = 2.38389191691868e-07 wdsub = 1.58974455775539e-07 pdsub = -4.03370655872948e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.447649365780035 lpclm = 4.80833966667745e-08 wpclm = 1.02458836160157e-07 ppclm = -2.59971878754252e-14
+ pdiblc1 = -1.15509388340255 lpdiblc1 = 4.10297474324608e-07 wpdiblc1 = 6.27749769338394e-07 ppdiblc1 = -1.59280832223539e-13
+ pdiblc2 = -0.0155920557246656 lpdiblc2 = 6.76439230630858e-09 wpdiblc2 = 3.62554742468736e-09 ppdiblc2 = -9.19921024708198e-16
+ pdiblcb = -1.62129269786215 lpdiblcb = 3.54285535106658e-07 wpdiblcb = 8.10453242464065e-07 ppdiblcb = -2.05638732570135e-13
+ drout = 1.08388936285629 ldrout = -1.65487142296144e-07 wdrout = 9.3584535245824e-08 pdrout = -2.37454848815288e-14
+ pscbe1 = 800072202.262479 lpscbe1 = -0.0363706622861173
+ pscbe2 = -6.5212424568799e-08 lpscbe2 = 1.88833418033178e-14 wpscbe2 = 3.35955119995127e-14 ppscbe2 = -8.52429004617235e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.11752930476661 lbeta0 = 5.52030039019352e-07 wbeta0 = 9.88902484429397e-07 pbeta0 = -2.50917194081725e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.77806705459672e-09 lagidl = 4.7652758796399e-16 wagidl = 1.3572684765143e-15 pagidl = -3.44383802351402e-22
+ bgidl = 718501708.262399 lbgidl = 141.799978991857
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.506690131559999 lkt1 = -1.3650501588864e-9
+ kt2 = 0.0185874300836493 lkt2 = -9.17991533341455e-09 wkt2 = -8.88418844389108e-08 pkt2 = 2.25421178643381e-14
+ at = 156265.507045123 lat = -0.0227622623510802 wat = -0.0528374991424447 pat = 1.34066171699099e-8
+ ute = 0.361190373811001 lute = -1.38655030028187e-07 wute = -2.08124392664772e-07 pute = 5.28080265240106e-14
+ ua1 = -3.46129801756714e-10 lua1 = 1.89962234809136e-16 wua1 = 3.2916558442678e-16 pua1 = -8.35201712333602e-23
+ ub1 = 6.16897967224791e-19 lub1 = -4.51385849178483e-26 wub1 = -5.88389054028908e-26 pub1 = 1.49293719845917e-32
+ uc1 = 4.842226005912e-11 luc1 = -1.21411037663607e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.24e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.106 pmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.895472038957143+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.69034288422874e-8
+ k1 = -0.475192721214427 lk1 = 2.6779954931801e-7
+ k2 = 0.424510226624299 lk2 = -1.12009306180152e-07 wk2 = -5.29395592033938e-23 pk2 = 9.46633086265214e-30
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 227262.218143857 lvsat = -0.0199381940412253
+ ua = 8.02797630049995e-10 lua = -6.02778297117977e-16
+ ub = -6.96694930414282e-19 lub = 5.83546908955007e-25
+ uc = 3.13756247644295e-15 luc = 1.32689039345937e-20
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.011653454326 lu0 = -1.55810440540896e-9
+ a0 = -0.470320092428571 la0 = 3.25394834642178e-7
+ keta = -0.194608099147397 lketa = 4.68488687339417e-08 wketa = -1.32348898008484e-23 pketa = -4.73316543132607e-30
+ a1 = 0.0
+ a2 = 0.143440229652999 la2 = 9.64903541390354e-8
+ ags = -1.75201096157886 lags = 5.51568480003768e-7
+ b0 = -1.44631992842857e-07 lb0 = 3.66979094399967e-14
+ b1 = -3.57990626714285e-08 lb1 = 9.08340356880958e-15
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.251108260161858+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope/sqrt(l*w*mult))} lvoff = -3.55783777856817e-8
+ nfactor = {-2.04597080806715+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = 1.1577432867533e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = 1.45153429224443 leta0 = -2.43972980574055e-7
+ etab = 0.259331250696142 letab = -6.58167545453844e-08 wetab = 4.66840058209615e-23 petab = -1.91052250483214e-30
+ dsub = 1.59102145467071 ldsub = -2.44350249175394e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.666465439125856 lpclm = -7.43746207148098e-9
+ pdiblc1 = 1.23047101218629 lpdiblc1 = -1.94999063327833e-7
+ pdiblc2 = 0.0312405399469343 lpdiblc2 = -5.11858269123347e-9
+ pdiblcb = -0.815555173997886 lpdiblcb = 1.49843335964006e-7
+ drout = -1.060023465579 ldrout = 3.78494291401226e-7
+ pscbe1 = 799742134.776859 lpscbe1 = 0.047378351043335
+ pscbe2 = 3.07580668600386e-08 lpscbe2 = -5.46753889839546e-15
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 11.69992923758 lbeta0 = -6.10676043133186e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = -1.17521467858986e-08 lagidl = 3.0072807604264e-15 wagidl = -2.95822839457879e-31 pagidl = 3.29138418230241e-37
+ bgidl = 2005351041.92 lbgidl = -184.716162985088
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.221955593000001 lkt1 = -7.3611598831331e-8
+ kt2 = 0.251204129485714 lkt2 = -6.82024483227987e-08 wkt2 = 5.29395592033938e-23 pkt2 = 6.31088724176809e-30
+ at = -8590.79699999979 lat = 0.019067222243201
+ ute = -0.324802089714286 lute = 3.54038957194749e-8
+ ua1 = 1.02463369042857e-09 lua1 = -1.57845698353513e-16
+ ub1 = 6.13178883999999e-19 lub1 = -4.41949307739717e-26
+ uc1 = -6.17595002111428e-11 luc1 = 1.58156448122939e-17 wuc1 = 1.07852076885685e-32 puc1 = 8.26519465421921e-40
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8__model.107 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = -1.8665e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.52161e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -2.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25.0e+6
+ tnoib = .0e-6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+sky130_fd_pr__pfet_01v8__toxe_slope_spectre*(4.075605e-09*(sky130_fd_pr__pfet_01v8__toxe_slope1/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.233669742410836+sky130_fd_pr__pfet_01v8__vth0_slope_spectre*(sky130_fd_pr__pfet_01v8__vth0_slope1/sqrt(l*w*mult))} lvth0 = -1.3849835019363e-07 wvth0 = -2.82854101681267e-07 pvth0 = 5.19696326642044e-14
+ k1 = -3.73744999519629 lk1 = 8.67183865038519e-07 wk1 = 2.0210577924838e-06 pk1 = -3.71335011386425e-13
+ k2 = 1.02672245256729 lk2 = -2.22655565089337e-07 wk2 = -4.74843564717764e-07 pk2 = 8.7244432676289e-14
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ w0 = 0.0
+ k3b = 2.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 783459.568999875 lvsat = -0.122130001906054 wvsat = -0.310391307820318 pvsat = 5.70291261597504e-8
+ ua = -1.12852673699409e-09 lua = -2.47930277187866e-16 wua = -5.54433613723269e-16 pua = 1.01867751150217e-22
+ ub = 1.5267370666053e-18 lub = 1.75029077846608e-25 wub = 2.00266186697553e-25 pub = -3.67955072805007e-32
+ uc = 8.54868350516763e-13 luc = -1.43222148944418e-19 wuc = -6.98117334484663e-19 puc = 1.28267192216871e-25
+ rdsw = 547.88
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1.0
+ u0 = 0.00679387706662439 lu0 = -6.65239696812094e-10 wu0 = -1.71623163859876e-09 pu0 = 3.15328387654667e-16
+ a0 = 8.65828800305226 la0 = -1.3518317165648e-06 wa0 = -2.3218883719601e-06 pa0 = 4.26607516245345e-13
+ keta = 1.16054493462406 lketa = -2.0213746361999e-07 wketa = -3.84654494537373e-07 pketa = 7.06737242448352e-14
+ a1 = 0.0
+ a2 = -4.57882396553973 la2 = 9.64126121514382e-07 wa2 = 2.65496221663659e-06 pa2 = -4.8780417294929e-13
+ ags = -13.0499332375962 lags = 2.62736963354326e-06 wags = 6.44115038806357e-06 pags = -1.18345188425008e-12
+ b0 = -6.0977537441079e-06 lb0 = 1.13048282816518e-12 wb0 = 2.58748740468979e-12 pb0 = -4.7540682332587e-19
+ b1 = -5.0222040431473e-08 lb1 = 1.17333805415958e-14 wb1 = 4.62340621934893e-14 pb1 = -8.49472294899636e-21
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.420632381326312+sky130_fd_pr__pfet_01v8__voff_slope_spectre*(sky130_fd_pr__pfet_01v8__voff_slope1/sqrt(l*w*mult))} lvoff = -4.43120243177315e-09 wvoff = 9.38934221448478e-09 pvoff = -1.72513201309396e-15
+ nfactor = {7.71690314501171+sky130_fd_pr__pfet_01v8__nfactor_slope_spectre*(sky130_fd_pr__pfet_01v8__nfactor_slope1/sqrt(l*w*mult))} lnfactor = -6.36018833267731e-07 wnfactor = -3.14946489374756e-06 pnfactor = 5.78660633322921e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0.0
+ eta0 = -1.98586831984566 leta0 = 3.87591313553092e-07 weta0 = 1.05795600376902e-06 peta0 = -1.94381430440494e-13
+ etab = -0.922404099585086 letab = 1.51307026567837e-07 wetab = 2.50210825583231e-07 petab = -4.59719856168837e-14
+ dsub = 0.266743858520667 ldsub = -1.03675360195782e-9
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.68745274242588 lpclm = -5.62492522268703e-07 wpclm = -1.75178328475506e-06 ppclm = 3.21860398257902e-13
+ pdiblc1 = 2.61300083018655 lpdiblc1 = -4.49015414378475e-07 wpdiblc1 = -1.44447692726621e-06 ppdiblc1 = 2.65398079277402e-13
+ pdiblc2 = 0.0598055254345681 lpdiblc2 = -1.03669131698329e-08 wpdiblc2 = -3.35019690444118e-08 ppdiblc2 = 6.15541727843691e-15
+ pdiblcb = 1.713355663646 lpdiblcb = -3.14801038968818e-07 wpdiblcb = -7.71428401893897e-07 ppdiblcb = 1.41736854565171e-13
+ drout = -0.60355488200225 ldrout = 2.94625949134919e-07 wdrout = 9.30754887981309e-07 pdrout = -1.7101038783347e-13
+ pscbe1 = 747355239.108776 lpscbe1 = 9.67257985282731 wpscbe1 = 30.5567143825683 ppscbe1 = -5.61427680365219e-6
+ pscbe2 = -6.52517064117004e-08 lpscbe2 = 1.2172624774141e-14 wpscbe2 = 1.34643550732985e-14 ppscbe2 = -2.47384635068235e-21
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 28.7068524242102 lbeta0 = -3.7354090609823e-06 wbeta0 = -9.96835010516876e-06 pbeta0 = 1.83151486987297e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 2.6872205821541e-08 lagidl = -4.08928741719629e-15 wagidl = -3.69201072031463e-15 pagidl = 6.78344205675566e-22
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.170264511828361 lkt1 = -8.31089562482399e-08 wkt1 = -2.03746469075227e-07 pkt1 = 3.74349500025985e-14
+ kt2 = -0.12
+ at = 382882.576833005 lat = -0.0528593551512584 wat = -0.0583310579143037 pat = 1.07173402637688e-8
+ ute = -3.68743648343475 lute = 6.53230800780916e-07 wute = 1.67067982305438e-06 pute = -3.0695901592925e-13
+ ua1 = -1.31186963806207e-10 lua1 = 5.45166979110061e-17 wua1 = 2.14876776945801e-16 pua1 = -3.94799548585828e-23
+ ub1 = 3.7264e-19
+ uc1 = 2.60259203177738e-10 luc1 = -4.33498176174554e-17 wuc1 = -1.37850924145181e-16 puc1 = 2.53277638459666e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.0
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 8.04e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 4.86838e-11
+ cgso = 4.86838e-11
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 8.8560258e-12
+ cgdl = 8.8560258e-12
+ cf = 1.2e-11
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 9.1275e-9
+ dwc = -2.252e-8
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0006889421079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.2317732e-11
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.ends sky130_fd_pr__pfet_01v8
