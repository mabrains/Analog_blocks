magic
tech sky130A
magscale 1 2
timestamp 1624884095
<< checkpaint >>
rect -1260 -1394 8305 2381
<< nwell >>
rect 0 953 7045 1121
rect 2042 417 2199 953
<< pwell >>
rect 66 10 6979 96
<< mvpsubdiff >>
rect 92 36 116 70
rect 150 36 185 70
rect 219 36 254 70
rect 288 36 323 70
rect 357 36 392 70
rect 426 36 461 70
rect 495 36 530 70
rect 564 36 599 70
rect 633 36 668 70
rect 702 36 737 70
rect 771 36 806 70
rect 840 36 875 70
rect 909 36 944 70
rect 978 36 1013 70
rect 1047 36 1082 70
rect 1116 36 1151 70
rect 1185 36 1220 70
rect 1254 36 1289 70
rect 1323 36 1358 70
rect 1392 36 1427 70
rect 1461 36 1496 70
rect 1530 36 1565 70
rect 1599 36 1634 70
rect 1668 36 1703 70
rect 1737 36 1772 70
rect 1806 36 1841 70
rect 1875 36 1910 70
rect 1944 36 1979 70
rect 2013 36 2048 70
rect 2082 36 2117 70
rect 2151 36 2186 70
rect 2220 36 2255 70
rect 2289 36 2324 70
rect 2358 36 2393 70
rect 2427 36 2462 70
rect 2496 36 2531 70
rect 2565 36 2600 70
rect 2634 36 2669 70
rect 2703 36 2738 70
rect 2772 36 2807 70
rect 2841 36 2876 70
rect 2910 36 2945 70
rect 2979 36 3014 70
rect 3048 36 3083 70
rect 3117 36 3152 70
rect 3186 36 3221 70
rect 3255 36 3290 70
rect 3324 36 3359 70
rect 3393 36 3427 70
rect 3461 36 3495 70
rect 3529 36 3563 70
rect 3597 36 3631 70
rect 3665 36 3699 70
rect 3733 36 3767 70
rect 3801 36 3835 70
rect 3869 36 3903 70
rect 3937 36 3971 70
rect 4005 36 4039 70
rect 4073 36 4107 70
rect 4141 36 4175 70
rect 4209 36 4243 70
rect 4277 36 4311 70
rect 4345 36 4379 70
rect 4413 36 4447 70
rect 4481 36 4515 70
rect 4549 36 4583 70
rect 4617 36 4651 70
rect 4685 36 4719 70
rect 4753 36 4787 70
rect 4821 36 4855 70
rect 4889 36 4923 70
rect 4957 36 4991 70
rect 5025 36 5059 70
rect 5093 36 5127 70
rect 5161 36 5195 70
rect 5229 36 5263 70
rect 5297 36 5331 70
rect 5365 36 5399 70
rect 5433 36 5467 70
rect 5501 36 5535 70
rect 5569 36 5603 70
rect 5637 36 5671 70
rect 5705 36 5739 70
rect 5773 36 5807 70
rect 5841 36 5875 70
rect 5909 36 5943 70
rect 5977 36 6011 70
rect 6045 36 6079 70
rect 6113 36 6147 70
rect 6181 36 6215 70
rect 6249 36 6283 70
rect 6317 36 6351 70
rect 6385 36 6419 70
rect 6453 36 6487 70
rect 6521 36 6555 70
rect 6589 36 6623 70
rect 6657 36 6691 70
rect 6725 36 6759 70
rect 6793 36 6827 70
rect 6861 36 6895 70
rect 6929 36 6953 70
<< mvnsubdiff >>
rect 67 1020 110 1054
rect 144 1020 178 1054
rect 212 1020 246 1054
rect 280 1020 314 1054
rect 348 1020 382 1054
rect 416 1020 450 1054
rect 484 1020 518 1054
rect 552 1020 586 1054
rect 620 1020 654 1054
rect 688 1020 722 1054
rect 756 1020 790 1054
rect 824 1020 858 1054
rect 892 1020 926 1054
rect 960 1020 994 1054
rect 1028 1020 1062 1054
rect 1096 1020 1130 1054
rect 1164 1020 1198 1054
rect 1232 1020 1266 1054
rect 1300 1020 1334 1054
rect 1368 1020 1402 1054
rect 1436 1020 1470 1054
rect 1504 1020 1538 1054
rect 1572 1020 1606 1054
rect 1640 1020 1674 1054
rect 1708 1020 1742 1054
rect 1776 1020 1810 1054
rect 1844 1020 1878 1054
rect 1912 1020 1946 1054
rect 1980 1020 2014 1054
rect 2048 1020 2082 1054
rect 2116 1020 2150 1054
rect 2184 1020 2218 1054
rect 2252 1020 2286 1054
rect 2320 1020 2354 1054
rect 2388 1020 2422 1054
rect 2456 1020 2490 1054
rect 2524 1020 2558 1054
rect 2592 1020 2626 1054
rect 2660 1020 2694 1054
rect 2728 1020 2762 1054
rect 2796 1020 2830 1054
rect 2864 1020 2898 1054
rect 2932 1020 2966 1054
rect 3000 1020 3034 1054
rect 3068 1020 3102 1054
rect 3136 1020 3170 1054
rect 3204 1020 3238 1054
rect 3272 1020 3306 1054
rect 3340 1020 3374 1054
rect 3408 1020 3442 1054
rect 3476 1020 3510 1054
rect 3544 1020 3578 1054
rect 3612 1020 3646 1054
rect 3680 1020 3714 1054
rect 3748 1020 3782 1054
rect 3816 1020 3850 1054
rect 3884 1020 3918 1054
rect 3952 1020 3986 1054
rect 4020 1020 4054 1054
rect 4088 1020 4122 1054
rect 4156 1020 4190 1054
rect 4224 1020 4258 1054
rect 4292 1020 4326 1054
rect 4360 1020 4394 1054
rect 4428 1020 4462 1054
rect 4496 1020 4530 1054
rect 4564 1020 4598 1054
rect 4632 1020 4666 1054
rect 4700 1020 4734 1054
rect 4768 1020 4802 1054
rect 4836 1020 4870 1054
rect 4904 1020 4938 1054
rect 4972 1020 5006 1054
rect 5040 1020 5074 1054
rect 5108 1020 5142 1054
rect 5176 1020 5210 1054
rect 5244 1020 5278 1054
rect 5312 1020 5346 1054
rect 5380 1020 5414 1054
rect 5448 1020 5482 1054
rect 5516 1020 5550 1054
rect 5584 1020 5618 1054
rect 5652 1020 5686 1054
rect 5720 1020 5754 1054
rect 5788 1020 5822 1054
rect 5856 1020 5890 1054
rect 5924 1020 5958 1054
rect 5992 1020 6026 1054
rect 6060 1020 6094 1054
rect 6128 1020 6162 1054
rect 6196 1020 6230 1054
rect 6264 1020 6298 1054
rect 6332 1020 6366 1054
rect 6400 1020 6434 1054
rect 6468 1020 6502 1054
rect 6536 1020 6570 1054
rect 6604 1020 6638 1054
rect 6672 1020 6706 1054
rect 6740 1020 6774 1054
rect 6808 1020 6842 1054
rect 6876 1020 6910 1054
rect 6944 1020 6978 1054
<< mvpsubdiffcont >>
rect 116 36 150 70
rect 185 36 219 70
rect 254 36 288 70
rect 323 36 357 70
rect 392 36 426 70
rect 461 36 495 70
rect 530 36 564 70
rect 599 36 633 70
rect 668 36 702 70
rect 737 36 771 70
rect 806 36 840 70
rect 875 36 909 70
rect 944 36 978 70
rect 1013 36 1047 70
rect 1082 36 1116 70
rect 1151 36 1185 70
rect 1220 36 1254 70
rect 1289 36 1323 70
rect 1358 36 1392 70
rect 1427 36 1461 70
rect 1496 36 1530 70
rect 1565 36 1599 70
rect 1634 36 1668 70
rect 1703 36 1737 70
rect 1772 36 1806 70
rect 1841 36 1875 70
rect 1910 36 1944 70
rect 1979 36 2013 70
rect 2048 36 2082 70
rect 2117 36 2151 70
rect 2186 36 2220 70
rect 2255 36 2289 70
rect 2324 36 2358 70
rect 2393 36 2427 70
rect 2462 36 2496 70
rect 2531 36 2565 70
rect 2600 36 2634 70
rect 2669 36 2703 70
rect 2738 36 2772 70
rect 2807 36 2841 70
rect 2876 36 2910 70
rect 2945 36 2979 70
rect 3014 36 3048 70
rect 3083 36 3117 70
rect 3152 36 3186 70
rect 3221 36 3255 70
rect 3290 36 3324 70
rect 3359 36 3393 70
rect 3427 36 3461 70
rect 3495 36 3529 70
rect 3563 36 3597 70
rect 3631 36 3665 70
rect 3699 36 3733 70
rect 3767 36 3801 70
rect 3835 36 3869 70
rect 3903 36 3937 70
rect 3971 36 4005 70
rect 4039 36 4073 70
rect 4107 36 4141 70
rect 4175 36 4209 70
rect 4243 36 4277 70
rect 4311 36 4345 70
rect 4379 36 4413 70
rect 4447 36 4481 70
rect 4515 36 4549 70
rect 4583 36 4617 70
rect 4651 36 4685 70
rect 4719 36 4753 70
rect 4787 36 4821 70
rect 4855 36 4889 70
rect 4923 36 4957 70
rect 4991 36 5025 70
rect 5059 36 5093 70
rect 5127 36 5161 70
rect 5195 36 5229 70
rect 5263 36 5297 70
rect 5331 36 5365 70
rect 5399 36 5433 70
rect 5467 36 5501 70
rect 5535 36 5569 70
rect 5603 36 5637 70
rect 5671 36 5705 70
rect 5739 36 5773 70
rect 5807 36 5841 70
rect 5875 36 5909 70
rect 5943 36 5977 70
rect 6011 36 6045 70
rect 6079 36 6113 70
rect 6147 36 6181 70
rect 6215 36 6249 70
rect 6283 36 6317 70
rect 6351 36 6385 70
rect 6419 36 6453 70
rect 6487 36 6521 70
rect 6555 36 6589 70
rect 6623 36 6657 70
rect 6691 36 6725 70
rect 6759 36 6793 70
rect 6827 36 6861 70
rect 6895 36 6929 70
<< mvnsubdiffcont >>
rect 110 1020 144 1054
rect 178 1020 212 1054
rect 246 1020 280 1054
rect 314 1020 348 1054
rect 382 1020 416 1054
rect 450 1020 484 1054
rect 518 1020 552 1054
rect 586 1020 620 1054
rect 654 1020 688 1054
rect 722 1020 756 1054
rect 790 1020 824 1054
rect 858 1020 892 1054
rect 926 1020 960 1054
rect 994 1020 1028 1054
rect 1062 1020 1096 1054
rect 1130 1020 1164 1054
rect 1198 1020 1232 1054
rect 1266 1020 1300 1054
rect 1334 1020 1368 1054
rect 1402 1020 1436 1054
rect 1470 1020 1504 1054
rect 1538 1020 1572 1054
rect 1606 1020 1640 1054
rect 1674 1020 1708 1054
rect 1742 1020 1776 1054
rect 1810 1020 1844 1054
rect 1878 1020 1912 1054
rect 1946 1020 1980 1054
rect 2014 1020 2048 1054
rect 2082 1020 2116 1054
rect 2150 1020 2184 1054
rect 2218 1020 2252 1054
rect 2286 1020 2320 1054
rect 2354 1020 2388 1054
rect 2422 1020 2456 1054
rect 2490 1020 2524 1054
rect 2558 1020 2592 1054
rect 2626 1020 2660 1054
rect 2694 1020 2728 1054
rect 2762 1020 2796 1054
rect 2830 1020 2864 1054
rect 2898 1020 2932 1054
rect 2966 1020 3000 1054
rect 3034 1020 3068 1054
rect 3102 1020 3136 1054
rect 3170 1020 3204 1054
rect 3238 1020 3272 1054
rect 3306 1020 3340 1054
rect 3374 1020 3408 1054
rect 3442 1020 3476 1054
rect 3510 1020 3544 1054
rect 3578 1020 3612 1054
rect 3646 1020 3680 1054
rect 3714 1020 3748 1054
rect 3782 1020 3816 1054
rect 3850 1020 3884 1054
rect 3918 1020 3952 1054
rect 3986 1020 4020 1054
rect 4054 1020 4088 1054
rect 4122 1020 4156 1054
rect 4190 1020 4224 1054
rect 4258 1020 4292 1054
rect 4326 1020 4360 1054
rect 4394 1020 4428 1054
rect 4462 1020 4496 1054
rect 4530 1020 4564 1054
rect 4598 1020 4632 1054
rect 4666 1020 4700 1054
rect 4734 1020 4768 1054
rect 4802 1020 4836 1054
rect 4870 1020 4904 1054
rect 4938 1020 4972 1054
rect 5006 1020 5040 1054
rect 5074 1020 5108 1054
rect 5142 1020 5176 1054
rect 5210 1020 5244 1054
rect 5278 1020 5312 1054
rect 5346 1020 5380 1054
rect 5414 1020 5448 1054
rect 5482 1020 5516 1054
rect 5550 1020 5584 1054
rect 5618 1020 5652 1054
rect 5686 1020 5720 1054
rect 5754 1020 5788 1054
rect 5822 1020 5856 1054
rect 5890 1020 5924 1054
rect 5958 1020 5992 1054
rect 6026 1020 6060 1054
rect 6094 1020 6128 1054
rect 6162 1020 6196 1054
rect 6230 1020 6264 1054
rect 6298 1020 6332 1054
rect 6366 1020 6400 1054
rect 6434 1020 6468 1054
rect 6502 1020 6536 1054
rect 6570 1020 6604 1054
rect 6638 1020 6672 1054
rect 6706 1020 6740 1054
rect 6774 1020 6808 1054
rect 6842 1020 6876 1054
rect 6910 1020 6944 1054
<< locali >>
rect 67 1020 79 1054
rect 144 1020 152 1054
rect 212 1020 225 1054
rect 280 1020 298 1054
rect 348 1020 371 1054
rect 416 1020 444 1054
rect 484 1020 517 1054
rect 552 1020 586 1054
rect 624 1020 654 1054
rect 697 1020 722 1054
rect 770 1020 790 1054
rect 843 1020 858 1054
rect 916 1020 926 1054
rect 989 1020 994 1054
rect 1096 1020 1101 1054
rect 1164 1020 1173 1054
rect 1232 1020 1245 1054
rect 1300 1020 1317 1054
rect 1368 1020 1389 1054
rect 1436 1020 1461 1054
rect 1504 1020 1533 1054
rect 1572 1020 1605 1054
rect 1640 1020 1674 1054
rect 1711 1020 1742 1054
rect 1783 1020 1810 1054
rect 1855 1020 1878 1054
rect 1927 1020 1946 1054
rect 1999 1020 2014 1054
rect 2071 1020 2082 1054
rect 2143 1020 2150 1054
rect 2215 1020 2218 1054
rect 2252 1020 2253 1054
rect 2320 1020 2325 1054
rect 2388 1020 2397 1054
rect 2456 1020 2469 1054
rect 2524 1020 2541 1054
rect 2592 1020 2613 1054
rect 2660 1020 2685 1054
rect 2728 1020 2757 1054
rect 2796 1020 2829 1054
rect 2864 1020 2898 1054
rect 2935 1020 2966 1054
rect 3007 1020 3034 1054
rect 3079 1020 3102 1054
rect 3151 1020 3170 1054
rect 3223 1020 3238 1054
rect 3295 1020 3306 1054
rect 3367 1020 3374 1054
rect 3439 1020 3442 1054
rect 3476 1020 3477 1054
rect 3544 1020 3549 1054
rect 3612 1020 3621 1054
rect 3680 1020 3693 1054
rect 3748 1020 3765 1054
rect 3816 1020 3837 1054
rect 3884 1020 3909 1054
rect 3952 1020 3981 1054
rect 4020 1020 4053 1054
rect 4088 1020 4122 1054
rect 4159 1020 4190 1054
rect 4231 1020 4258 1054
rect 4303 1020 4326 1054
rect 4375 1020 4394 1054
rect 4447 1020 4462 1054
rect 4519 1020 4530 1054
rect 4591 1020 4598 1054
rect 4663 1020 4666 1054
rect 4700 1020 4701 1054
rect 4768 1020 4773 1054
rect 4836 1020 4845 1054
rect 4904 1020 4917 1054
rect 4972 1020 4989 1054
rect 5040 1020 5061 1054
rect 5108 1020 5133 1054
rect 5176 1020 5205 1054
rect 5244 1020 5277 1054
rect 5312 1020 5346 1054
rect 5383 1020 5414 1054
rect 5455 1020 5482 1054
rect 5527 1020 5550 1054
rect 5599 1020 5618 1054
rect 5671 1020 5686 1054
rect 5743 1020 5754 1054
rect 5815 1020 5822 1054
rect 5887 1020 5890 1054
rect 5924 1020 5925 1054
rect 5992 1020 5997 1054
rect 6060 1020 6069 1054
rect 6128 1020 6141 1054
rect 6196 1020 6213 1054
rect 6264 1020 6285 1054
rect 6332 1020 6357 1054
rect 6400 1020 6429 1054
rect 6468 1020 6501 1054
rect 6536 1020 6570 1054
rect 6607 1020 6638 1054
rect 6679 1020 6706 1054
rect 6751 1020 6774 1054
rect 6823 1020 6842 1054
rect 6895 1020 6910 1054
rect 6967 1020 6978 1054
rect 173 402 211 436
rect 408 402 446 436
rect 292 315 326 353
rect 657 368 691 406
rect 775 334 949 436
rect 1155 396 1193 430
rect 1040 315 1074 353
rect 1405 368 1439 406
rect 1618 402 1656 436
rect 1502 315 1536 353
rect 1867 368 1901 406
rect 1964 376 1998 414
rect 2706 368 2740 406
rect 2801 315 2835 353
rect 2983 368 3017 406
rect 3207 396 3245 430
rect 3087 315 3121 353
rect 3448 368 3482 406
rect 3552 368 3586 406
rect 3734 380 3768 418
rect 3958 371 3996 405
rect 3838 315 3872 353
rect 4199 368 4233 406
rect 4303 368 4337 406
rect 4390 368 4424 406
rect 4667 380 4701 418
rect 4885 396 4923 430
rect 4765 315 4799 353
rect 5128 368 5162 406
rect 5230 368 5264 406
rect 5312 368 5346 406
rect 5516 429 5550 467
rect 5613 380 5647 418
rect 5893 368 5927 406
rect 6094 402 6132 436
rect 5978 315 6012 353
rect 6336 368 6370 406
rect 6458 334 6630 436
rect 6726 368 6760 406
rect 6828 368 6862 406
rect 112 36 116 70
rect 150 36 151 70
rect 219 36 224 70
rect 288 36 297 70
rect 357 36 370 70
rect 426 36 443 70
rect 495 36 516 70
rect 564 36 589 70
rect 633 36 662 70
rect 702 36 735 70
rect 771 36 806 70
rect 842 36 875 70
rect 915 36 944 70
rect 988 36 1013 70
rect 1061 36 1082 70
rect 1134 36 1151 70
rect 1207 36 1220 70
rect 1279 36 1289 70
rect 1351 36 1358 70
rect 1423 36 1427 70
rect 1495 36 1496 70
rect 1530 36 1533 70
rect 1599 36 1605 70
rect 1668 36 1677 70
rect 1737 36 1749 70
rect 1806 36 1821 70
rect 1875 36 1893 70
rect 1944 36 1965 70
rect 2013 36 2037 70
rect 2082 36 2109 70
rect 2151 36 2181 70
rect 2220 36 2253 70
rect 2289 36 2324 70
rect 2359 36 2393 70
rect 2431 36 2462 70
rect 2503 36 2531 70
rect 2575 36 2600 70
rect 2647 36 2669 70
rect 2719 36 2738 70
rect 2791 36 2807 70
rect 2863 36 2876 70
rect 2935 36 2945 70
rect 3007 36 3014 70
rect 3079 36 3083 70
rect 3151 36 3152 70
rect 3186 36 3189 70
rect 3255 36 3261 70
rect 3324 36 3333 70
rect 3393 36 3405 70
rect 3461 36 3477 70
rect 3529 36 3549 70
rect 3597 36 3621 70
rect 3665 36 3693 70
rect 3733 36 3765 70
rect 3801 36 3835 70
rect 3871 36 3903 70
rect 3943 36 3971 70
rect 4015 36 4039 70
rect 4087 36 4107 70
rect 4159 36 4175 70
rect 4231 36 4243 70
rect 4303 36 4311 70
rect 4375 36 4379 70
rect 4481 36 4485 70
rect 4549 36 4557 70
rect 4617 36 4629 70
rect 4685 36 4701 70
rect 4753 36 4773 70
rect 4821 36 4845 70
rect 4889 36 4917 70
rect 4957 36 4989 70
rect 5025 36 5059 70
rect 5095 36 5127 70
rect 5167 36 5195 70
rect 5239 36 5263 70
rect 5311 36 5331 70
rect 5383 36 5399 70
rect 5455 36 5467 70
rect 5527 36 5535 70
rect 5599 36 5603 70
rect 5705 36 5709 70
rect 5773 36 5781 70
rect 5841 36 5853 70
rect 5909 36 5925 70
rect 5977 36 5997 70
rect 6045 36 6069 70
rect 6113 36 6141 70
rect 6181 36 6213 70
rect 6249 36 6283 70
rect 6319 36 6351 70
rect 6391 36 6419 70
rect 6463 36 6487 70
rect 6535 36 6555 70
rect 6607 36 6623 70
rect 6679 36 6691 70
rect 6751 36 6759 70
rect 6823 36 6827 70
rect 6929 36 6933 70
<< viali >>
rect 79 1020 110 1054
rect 110 1020 113 1054
rect 152 1020 178 1054
rect 178 1020 186 1054
rect 225 1020 246 1054
rect 246 1020 259 1054
rect 298 1020 314 1054
rect 314 1020 332 1054
rect 371 1020 382 1054
rect 382 1020 405 1054
rect 444 1020 450 1054
rect 450 1020 478 1054
rect 517 1020 518 1054
rect 518 1020 551 1054
rect 590 1020 620 1054
rect 620 1020 624 1054
rect 663 1020 688 1054
rect 688 1020 697 1054
rect 736 1020 756 1054
rect 756 1020 770 1054
rect 809 1020 824 1054
rect 824 1020 843 1054
rect 882 1020 892 1054
rect 892 1020 916 1054
rect 955 1020 960 1054
rect 960 1020 989 1054
rect 1028 1020 1062 1054
rect 1101 1020 1130 1054
rect 1130 1020 1135 1054
rect 1173 1020 1198 1054
rect 1198 1020 1207 1054
rect 1245 1020 1266 1054
rect 1266 1020 1279 1054
rect 1317 1020 1334 1054
rect 1334 1020 1351 1054
rect 1389 1020 1402 1054
rect 1402 1020 1423 1054
rect 1461 1020 1470 1054
rect 1470 1020 1495 1054
rect 1533 1020 1538 1054
rect 1538 1020 1567 1054
rect 1605 1020 1606 1054
rect 1606 1020 1639 1054
rect 1677 1020 1708 1054
rect 1708 1020 1711 1054
rect 1749 1020 1776 1054
rect 1776 1020 1783 1054
rect 1821 1020 1844 1054
rect 1844 1020 1855 1054
rect 1893 1020 1912 1054
rect 1912 1020 1927 1054
rect 1965 1020 1980 1054
rect 1980 1020 1999 1054
rect 2037 1020 2048 1054
rect 2048 1020 2071 1054
rect 2109 1020 2116 1054
rect 2116 1020 2143 1054
rect 2181 1020 2184 1054
rect 2184 1020 2215 1054
rect 2253 1020 2286 1054
rect 2286 1020 2287 1054
rect 2325 1020 2354 1054
rect 2354 1020 2359 1054
rect 2397 1020 2422 1054
rect 2422 1020 2431 1054
rect 2469 1020 2490 1054
rect 2490 1020 2503 1054
rect 2541 1020 2558 1054
rect 2558 1020 2575 1054
rect 2613 1020 2626 1054
rect 2626 1020 2647 1054
rect 2685 1020 2694 1054
rect 2694 1020 2719 1054
rect 2757 1020 2762 1054
rect 2762 1020 2791 1054
rect 2829 1020 2830 1054
rect 2830 1020 2863 1054
rect 2901 1020 2932 1054
rect 2932 1020 2935 1054
rect 2973 1020 3000 1054
rect 3000 1020 3007 1054
rect 3045 1020 3068 1054
rect 3068 1020 3079 1054
rect 3117 1020 3136 1054
rect 3136 1020 3151 1054
rect 3189 1020 3204 1054
rect 3204 1020 3223 1054
rect 3261 1020 3272 1054
rect 3272 1020 3295 1054
rect 3333 1020 3340 1054
rect 3340 1020 3367 1054
rect 3405 1020 3408 1054
rect 3408 1020 3439 1054
rect 3477 1020 3510 1054
rect 3510 1020 3511 1054
rect 3549 1020 3578 1054
rect 3578 1020 3583 1054
rect 3621 1020 3646 1054
rect 3646 1020 3655 1054
rect 3693 1020 3714 1054
rect 3714 1020 3727 1054
rect 3765 1020 3782 1054
rect 3782 1020 3799 1054
rect 3837 1020 3850 1054
rect 3850 1020 3871 1054
rect 3909 1020 3918 1054
rect 3918 1020 3943 1054
rect 3981 1020 3986 1054
rect 3986 1020 4015 1054
rect 4053 1020 4054 1054
rect 4054 1020 4087 1054
rect 4125 1020 4156 1054
rect 4156 1020 4159 1054
rect 4197 1020 4224 1054
rect 4224 1020 4231 1054
rect 4269 1020 4292 1054
rect 4292 1020 4303 1054
rect 4341 1020 4360 1054
rect 4360 1020 4375 1054
rect 4413 1020 4428 1054
rect 4428 1020 4447 1054
rect 4485 1020 4496 1054
rect 4496 1020 4519 1054
rect 4557 1020 4564 1054
rect 4564 1020 4591 1054
rect 4629 1020 4632 1054
rect 4632 1020 4663 1054
rect 4701 1020 4734 1054
rect 4734 1020 4735 1054
rect 4773 1020 4802 1054
rect 4802 1020 4807 1054
rect 4845 1020 4870 1054
rect 4870 1020 4879 1054
rect 4917 1020 4938 1054
rect 4938 1020 4951 1054
rect 4989 1020 5006 1054
rect 5006 1020 5023 1054
rect 5061 1020 5074 1054
rect 5074 1020 5095 1054
rect 5133 1020 5142 1054
rect 5142 1020 5167 1054
rect 5205 1020 5210 1054
rect 5210 1020 5239 1054
rect 5277 1020 5278 1054
rect 5278 1020 5311 1054
rect 5349 1020 5380 1054
rect 5380 1020 5383 1054
rect 5421 1020 5448 1054
rect 5448 1020 5455 1054
rect 5493 1020 5516 1054
rect 5516 1020 5527 1054
rect 5565 1020 5584 1054
rect 5584 1020 5599 1054
rect 5637 1020 5652 1054
rect 5652 1020 5671 1054
rect 5709 1020 5720 1054
rect 5720 1020 5743 1054
rect 5781 1020 5788 1054
rect 5788 1020 5815 1054
rect 5853 1020 5856 1054
rect 5856 1020 5887 1054
rect 5925 1020 5958 1054
rect 5958 1020 5959 1054
rect 5997 1020 6026 1054
rect 6026 1020 6031 1054
rect 6069 1020 6094 1054
rect 6094 1020 6103 1054
rect 6141 1020 6162 1054
rect 6162 1020 6175 1054
rect 6213 1020 6230 1054
rect 6230 1020 6247 1054
rect 6285 1020 6298 1054
rect 6298 1020 6319 1054
rect 6357 1020 6366 1054
rect 6366 1020 6391 1054
rect 6429 1020 6434 1054
rect 6434 1020 6463 1054
rect 6501 1020 6502 1054
rect 6502 1020 6535 1054
rect 6573 1020 6604 1054
rect 6604 1020 6607 1054
rect 6645 1020 6672 1054
rect 6672 1020 6679 1054
rect 6717 1020 6740 1054
rect 6740 1020 6751 1054
rect 6789 1020 6808 1054
rect 6808 1020 6823 1054
rect 6861 1020 6876 1054
rect 6876 1020 6895 1054
rect 6933 1020 6944 1054
rect 6944 1020 6967 1054
rect 5516 467 5550 501
rect 139 402 173 436
rect 211 402 245 436
rect 374 402 408 436
rect 446 402 480 436
rect 657 406 691 440
rect 292 353 326 387
rect 657 334 691 368
rect 1121 396 1155 430
rect 1193 396 1227 430
rect 1405 406 1439 440
rect 1040 353 1074 387
rect 292 281 326 315
rect 1584 402 1618 436
rect 1656 402 1690 436
rect 1867 406 1901 440
rect 1405 334 1439 368
rect 1502 353 1536 387
rect 1040 281 1074 315
rect 1867 334 1901 368
rect 1964 414 1998 448
rect 1964 342 1998 376
rect 2706 406 2740 440
rect 2983 406 3017 440
rect 2706 334 2740 368
rect 2801 353 2835 387
rect 1502 281 1536 315
rect 3173 396 3207 430
rect 3245 396 3279 430
rect 3448 406 3482 440
rect 2983 334 3017 368
rect 3087 353 3121 387
rect 2801 281 2835 315
rect 3448 334 3482 368
rect 3552 406 3586 440
rect 3552 334 3586 368
rect 3734 418 3768 452
rect 4199 406 4233 440
rect 3734 346 3768 380
rect 3838 353 3872 387
rect 3924 371 3958 405
rect 3996 371 4030 405
rect 3087 281 3121 315
rect 4199 334 4233 368
rect 4303 406 4337 440
rect 4303 334 4337 368
rect 4390 406 4424 440
rect 4390 334 4424 368
rect 4667 418 4701 452
rect 4851 396 4885 430
rect 4923 396 4957 430
rect 5128 406 5162 440
rect 4667 346 4701 380
rect 4765 353 4799 387
rect 3838 281 3872 315
rect 5128 334 5162 368
rect 5230 406 5264 440
rect 5230 334 5264 368
rect 5312 406 5346 440
rect 5516 395 5550 429
rect 5613 418 5647 452
rect 5312 334 5346 368
rect 5613 346 5647 380
rect 5893 406 5927 440
rect 6060 402 6094 436
rect 6132 402 6166 436
rect 6336 406 6370 440
rect 5893 334 5927 368
rect 5978 353 6012 387
rect 4765 281 4799 315
rect 6336 334 6370 368
rect 6726 406 6760 440
rect 6726 334 6760 368
rect 6828 406 6862 440
rect 6828 334 6862 368
rect 5978 281 6012 315
rect 78 36 112 70
rect 151 36 185 70
rect 224 36 254 70
rect 254 36 258 70
rect 297 36 323 70
rect 323 36 331 70
rect 370 36 392 70
rect 392 36 404 70
rect 443 36 461 70
rect 461 36 477 70
rect 516 36 530 70
rect 530 36 550 70
rect 589 36 599 70
rect 599 36 623 70
rect 662 36 668 70
rect 668 36 696 70
rect 735 36 737 70
rect 737 36 769 70
rect 808 36 840 70
rect 840 36 842 70
rect 881 36 909 70
rect 909 36 915 70
rect 954 36 978 70
rect 978 36 988 70
rect 1027 36 1047 70
rect 1047 36 1061 70
rect 1100 36 1116 70
rect 1116 36 1134 70
rect 1173 36 1185 70
rect 1185 36 1207 70
rect 1245 36 1254 70
rect 1254 36 1279 70
rect 1317 36 1323 70
rect 1323 36 1351 70
rect 1389 36 1392 70
rect 1392 36 1423 70
rect 1461 36 1495 70
rect 1533 36 1565 70
rect 1565 36 1567 70
rect 1605 36 1634 70
rect 1634 36 1639 70
rect 1677 36 1703 70
rect 1703 36 1711 70
rect 1749 36 1772 70
rect 1772 36 1783 70
rect 1821 36 1841 70
rect 1841 36 1855 70
rect 1893 36 1910 70
rect 1910 36 1927 70
rect 1965 36 1979 70
rect 1979 36 1999 70
rect 2037 36 2048 70
rect 2048 36 2071 70
rect 2109 36 2117 70
rect 2117 36 2143 70
rect 2181 36 2186 70
rect 2186 36 2215 70
rect 2253 36 2255 70
rect 2255 36 2287 70
rect 2325 36 2358 70
rect 2358 36 2359 70
rect 2397 36 2427 70
rect 2427 36 2431 70
rect 2469 36 2496 70
rect 2496 36 2503 70
rect 2541 36 2565 70
rect 2565 36 2575 70
rect 2613 36 2634 70
rect 2634 36 2647 70
rect 2685 36 2703 70
rect 2703 36 2719 70
rect 2757 36 2772 70
rect 2772 36 2791 70
rect 2829 36 2841 70
rect 2841 36 2863 70
rect 2901 36 2910 70
rect 2910 36 2935 70
rect 2973 36 2979 70
rect 2979 36 3007 70
rect 3045 36 3048 70
rect 3048 36 3079 70
rect 3117 36 3151 70
rect 3189 36 3221 70
rect 3221 36 3223 70
rect 3261 36 3290 70
rect 3290 36 3295 70
rect 3333 36 3359 70
rect 3359 36 3367 70
rect 3405 36 3427 70
rect 3427 36 3439 70
rect 3477 36 3495 70
rect 3495 36 3511 70
rect 3549 36 3563 70
rect 3563 36 3583 70
rect 3621 36 3631 70
rect 3631 36 3655 70
rect 3693 36 3699 70
rect 3699 36 3727 70
rect 3765 36 3767 70
rect 3767 36 3799 70
rect 3837 36 3869 70
rect 3869 36 3871 70
rect 3909 36 3937 70
rect 3937 36 3943 70
rect 3981 36 4005 70
rect 4005 36 4015 70
rect 4053 36 4073 70
rect 4073 36 4087 70
rect 4125 36 4141 70
rect 4141 36 4159 70
rect 4197 36 4209 70
rect 4209 36 4231 70
rect 4269 36 4277 70
rect 4277 36 4303 70
rect 4341 36 4345 70
rect 4345 36 4375 70
rect 4413 36 4447 70
rect 4485 36 4515 70
rect 4515 36 4519 70
rect 4557 36 4583 70
rect 4583 36 4591 70
rect 4629 36 4651 70
rect 4651 36 4663 70
rect 4701 36 4719 70
rect 4719 36 4735 70
rect 4773 36 4787 70
rect 4787 36 4807 70
rect 4845 36 4855 70
rect 4855 36 4879 70
rect 4917 36 4923 70
rect 4923 36 4951 70
rect 4989 36 4991 70
rect 4991 36 5023 70
rect 5061 36 5093 70
rect 5093 36 5095 70
rect 5133 36 5161 70
rect 5161 36 5167 70
rect 5205 36 5229 70
rect 5229 36 5239 70
rect 5277 36 5297 70
rect 5297 36 5311 70
rect 5349 36 5365 70
rect 5365 36 5383 70
rect 5421 36 5433 70
rect 5433 36 5455 70
rect 5493 36 5501 70
rect 5501 36 5527 70
rect 5565 36 5569 70
rect 5569 36 5599 70
rect 5637 36 5671 70
rect 5709 36 5739 70
rect 5739 36 5743 70
rect 5781 36 5807 70
rect 5807 36 5815 70
rect 5853 36 5875 70
rect 5875 36 5887 70
rect 5925 36 5943 70
rect 5943 36 5959 70
rect 5997 36 6011 70
rect 6011 36 6031 70
rect 6069 36 6079 70
rect 6079 36 6103 70
rect 6141 36 6147 70
rect 6147 36 6175 70
rect 6213 36 6215 70
rect 6215 36 6247 70
rect 6285 36 6317 70
rect 6317 36 6319 70
rect 6357 36 6385 70
rect 6385 36 6391 70
rect 6429 36 6453 70
rect 6453 36 6463 70
rect 6501 36 6521 70
rect 6521 36 6535 70
rect 6573 36 6589 70
rect 6589 36 6607 70
rect 6645 36 6657 70
rect 6657 36 6679 70
rect 6717 36 6725 70
rect 6725 36 6751 70
rect 6789 36 6793 70
rect 6793 36 6823 70
rect 6861 36 6895 70
rect 6933 36 6967 70
<< metal1 >>
rect 67 1054 6979 1064
rect 67 1020 79 1054
rect 113 1020 152 1054
rect 186 1020 225 1054
rect 259 1020 298 1054
rect 332 1020 371 1054
rect 405 1020 444 1054
rect 478 1020 517 1054
rect 551 1020 590 1054
rect 624 1020 663 1054
rect 697 1020 736 1054
rect 770 1020 809 1054
rect 843 1020 882 1054
rect 916 1020 955 1054
rect 989 1020 1028 1054
rect 1062 1020 1101 1054
rect 1135 1020 1173 1054
rect 1207 1020 1245 1054
rect 1279 1020 1317 1054
rect 1351 1020 1389 1054
rect 1423 1020 1461 1054
rect 1495 1020 1533 1054
rect 1567 1020 1605 1054
rect 1639 1020 1677 1054
rect 1711 1020 1749 1054
rect 1783 1020 1821 1054
rect 1855 1020 1893 1054
rect 1927 1020 1965 1054
rect 1999 1020 2037 1054
rect 2071 1020 2109 1054
rect 2143 1020 2181 1054
rect 2215 1020 2253 1054
rect 2287 1020 2325 1054
rect 2359 1020 2397 1054
rect 2431 1020 2469 1054
rect 2503 1020 2541 1054
rect 2575 1020 2613 1054
rect 2647 1020 2685 1054
rect 2719 1020 2757 1054
rect 2791 1020 2829 1054
rect 2863 1020 2901 1054
rect 2935 1020 2973 1054
rect 3007 1020 3045 1054
rect 3079 1020 3117 1054
rect 3151 1020 3189 1054
rect 3223 1020 3261 1054
rect 3295 1020 3333 1054
rect 3367 1020 3405 1054
rect 3439 1020 3477 1054
rect 3511 1020 3549 1054
rect 3583 1020 3621 1054
rect 3655 1020 3693 1054
rect 3727 1020 3765 1054
rect 3799 1020 3837 1054
rect 3871 1020 3909 1054
rect 3943 1020 3981 1054
rect 4015 1020 4053 1054
rect 4087 1020 4125 1054
rect 4159 1020 4197 1054
rect 4231 1020 4269 1054
rect 4303 1020 4341 1054
rect 4375 1020 4413 1054
rect 4447 1020 4485 1054
rect 4519 1020 4557 1054
rect 4591 1020 4629 1054
rect 4663 1020 4701 1054
rect 4735 1020 4773 1054
rect 4807 1020 4845 1054
rect 4879 1020 4917 1054
rect 4951 1020 4989 1054
rect 5023 1020 5061 1054
rect 5095 1020 5133 1054
rect 5167 1020 5205 1054
rect 5239 1020 5277 1054
rect 5311 1020 5349 1054
rect 5383 1020 5421 1054
rect 5455 1020 5493 1054
rect 5527 1020 5565 1054
rect 5599 1020 5637 1054
rect 5671 1020 5709 1054
rect 5743 1020 5781 1054
rect 5815 1020 5853 1054
rect 5887 1020 5925 1054
rect 5959 1020 5997 1054
rect 6031 1020 6069 1054
rect 6103 1020 6141 1054
rect 6175 1020 6213 1054
rect 6247 1020 6285 1054
rect 6319 1020 6357 1054
rect 6391 1020 6429 1054
rect 6463 1020 6501 1054
rect 6535 1020 6573 1054
rect 6607 1020 6645 1054
rect 6679 1020 6717 1054
rect 6751 1020 6789 1054
rect 6823 1020 6861 1054
rect 6895 1020 6933 1054
rect 6967 1020 6979 1054
rect 67 861 6979 1020
rect 1958 701 4508 753
tri 4508 701 4514 707 sw
rect 4658 701 4664 753
rect 4716 701 4728 753
rect 4780 701 5583 753
rect 1958 673 2010 701
tri 2010 673 2038 701 nw
tri 4399 673 4427 701 ne
rect 4427 673 4514 701
tri 4514 673 4542 701 sw
rect 127 436 257 442
rect 127 402 139 436
rect 173 402 211 436
rect 245 402 257 436
rect 127 396 257 402
rect 362 436 492 442
rect 362 402 374 436
rect 408 402 446 436
rect 480 402 492 436
rect 286 387 332 399
rect 362 396 492 402
rect 651 440 697 452
rect 651 406 657 440
rect 691 406 697 440
rect 1399 440 1445 452
rect 1861 451 1907 452
rect 286 353 292 387
rect 326 353 332 387
rect 651 368 697 406
rect 1109 430 1239 436
rect 286 334 332 353
tri 332 334 353 355 sw
tri 630 334 651 355 se
rect 651 334 657 368
rect 691 334 697 368
rect 286 321 353 334
tri 353 321 366 334 sw
tri 617 321 630 334 se
rect 630 321 697 334
rect 286 315 697 321
rect 286 281 292 315
rect 326 281 697 315
rect 286 269 697 281
rect 1034 387 1080 399
rect 1109 396 1121 430
rect 1155 396 1193 430
rect 1227 396 1239 430
rect 1109 390 1239 396
rect 1399 406 1405 440
rect 1439 406 1445 440
rect 1034 353 1040 387
rect 1074 353 1080 387
rect 1399 368 1445 406
rect 1572 436 1702 442
rect 1572 402 1584 436
rect 1618 402 1656 436
rect 1690 402 1702 436
rect 1034 334 1080 353
tri 1080 334 1101 355 sw
tri 1378 334 1399 355 se
rect 1399 334 1405 368
rect 1439 334 1445 368
rect 1034 321 1101 334
tri 1101 321 1114 334 sw
tri 1365 321 1378 334 se
rect 1378 321 1445 334
rect 1034 315 1445 321
rect 1034 281 1040 315
rect 1074 281 1445 315
rect 1034 269 1445 281
rect 1496 387 1542 399
rect 1572 396 1702 402
rect 1861 440 1913 451
rect 1861 406 1867 440
rect 1901 406 1913 440
rect 1496 353 1502 387
rect 1536 353 1542 387
rect 1861 368 1913 406
rect 1496 334 1542 353
tri 1542 334 1563 355 sw
tri 1840 334 1861 355 se
rect 1861 334 1867 368
rect 1901 334 1913 368
rect 1496 322 1563 334
tri 1563 322 1575 334 sw
tri 1828 322 1840 334 se
rect 1840 322 1913 334
rect 1958 448 2004 673
tri 2004 667 2010 673 nw
rect 3161 621 4224 673
rect 4276 621 4288 673
rect 4340 621 4346 673
tri 4427 667 4433 673 ne
rect 4433 621 4439 673
rect 4491 621 4503 673
rect 4555 621 5309 673
rect 5361 621 5373 673
rect 5425 621 5856 673
rect 5908 621 5920 673
rect 5972 621 5978 673
rect 3161 593 3233 621
tri 3233 593 3261 621 nw
rect 3161 467 3227 593
tri 3227 587 3233 593 nw
rect 3912 541 3918 593
rect 3970 541 3982 593
rect 4034 569 4040 593
tri 4040 569 4064 593 sw
rect 4034 541 5653 569
tri 5573 513 5601 541 ne
rect 5601 513 5653 541
rect 3728 485 4710 513
tri 5041 501 5053 513 se
rect 5053 501 5556 513
tri 5601 507 5607 513 ne
tri 5025 485 5041 501 se
rect 5041 485 5516 501
tri 3227 467 3230 470 sw
rect 3728 467 3790 485
tri 3790 467 3808 485 nw
tri 4624 467 4642 485 ne
rect 4642 467 4710 485
tri 5007 467 5025 485 se
rect 5025 467 5070 485
tri 5070 467 5088 485 nw
tri 5476 467 5494 485 ne
rect 5494 467 5516 485
rect 5550 467 5556 501
rect 3161 452 3230 467
tri 3230 452 3245 467 sw
rect 3728 452 3775 467
tri 3775 452 3790 467 nw
tri 4642 452 4657 467 ne
rect 4657 456 4710 467
tri 5000 460 5007 467 se
rect 5007 460 5063 467
tri 5063 460 5070 467 nw
tri 5494 460 5501 467 ne
rect 5501 460 5556 467
rect 4657 452 4658 456
tri 4992 452 5000 460 se
rect 5000 452 5055 460
tri 5055 452 5063 460 nw
tri 5501 452 5509 460 ne
rect 5509 452 5556 460
rect 1958 414 1964 448
rect 1998 414 2004 448
rect 1958 376 2004 414
rect 1958 342 1964 376
rect 1998 342 2004 376
rect 1958 330 2004 342
rect 2700 440 2746 452
rect 2700 406 2706 440
rect 2740 406 2746 440
rect 2700 368 2746 406
rect 2977 440 3023 452
rect 2977 406 2983 440
rect 3017 406 3023 440
rect 2700 334 2706 368
rect 2740 334 2746 368
rect 1496 321 1575 322
tri 1575 321 1576 322 sw
tri 1827 321 1828 322 se
rect 1828 321 1913 322
rect 1496 315 1913 321
rect 1496 281 1502 315
rect 1536 281 1913 315
rect 2700 306 2746 334
rect 2795 387 2841 399
rect 2795 353 2801 387
rect 2835 353 2841 387
rect 2977 368 3023 406
rect 3161 440 3245 452
tri 3245 440 3257 452 sw
rect 3442 440 3488 452
rect 3161 436 3257 440
tri 3257 436 3261 440 sw
rect 3161 430 3291 436
rect 2795 334 2841 353
tri 2841 334 2862 355 sw
tri 2956 334 2977 355 se
rect 2977 334 2983 368
rect 3017 334 3023 368
rect 2795 321 2862 334
tri 2862 321 2875 334 sw
tri 2943 321 2956 334 se
rect 2956 321 3023 334
rect 2795 315 3023 321
rect 1496 269 1913 281
rect 2795 281 2801 315
rect 2835 281 3023 315
rect 2795 269 3023 281
rect 3081 387 3127 399
rect 3161 396 3173 430
rect 3207 396 3245 430
rect 3279 396 3291 430
rect 3161 390 3291 396
rect 3442 406 3448 440
rect 3482 406 3488 440
rect 3081 353 3087 387
rect 3121 353 3127 387
rect 3442 368 3488 406
rect 3081 334 3127 353
tri 3127 334 3148 355 sw
tri 3421 334 3442 355 se
rect 3442 334 3448 368
rect 3482 334 3488 368
rect 3081 321 3148 334
tri 3148 321 3161 334 sw
tri 3408 321 3421 334 se
rect 3421 321 3488 334
rect 3546 440 3592 452
rect 3546 406 3552 440
rect 3586 406 3592 440
rect 3546 368 3592 406
rect 3546 334 3552 368
rect 3586 334 3592 368
rect 3728 418 3734 452
rect 3768 418 3774 452
tri 3774 451 3775 452 nw
rect 3728 380 3774 418
rect 4193 440 4239 452
rect 3728 346 3734 380
rect 3768 346 3774 380
rect 3728 334 3774 346
rect 3832 387 3878 399
rect 3832 353 3838 387
rect 3872 353 3878 387
rect 3912 362 3918 414
rect 3970 362 3982 414
rect 4034 362 4042 414
rect 4193 406 4199 440
rect 4233 406 4239 440
rect 4193 368 4239 406
rect 3832 334 3878 353
tri 3878 334 3899 355 sw
tri 4172 334 4193 355 se
rect 4193 334 4199 368
rect 4233 334 4239 368
rect 3546 322 3592 334
rect 3081 315 3488 321
rect 3081 281 3087 315
rect 3121 281 3488 315
rect 3081 269 3488 281
rect 3832 321 3899 334
tri 3899 321 3912 334 sw
tri 4159 321 4172 334 se
rect 4172 321 4239 334
rect 4294 445 4346 452
rect 4294 381 4346 393
rect 4294 322 4346 329
rect 4381 444 4433 452
tri 4657 451 4658 452 ne
rect 4381 380 4433 392
tri 4990 450 4992 452 se
rect 4992 450 5053 452
tri 5053 450 5055 452 nw
tri 4980 440 4990 450 se
rect 4990 440 5043 450
tri 5043 440 5053 450 nw
rect 5122 440 5168 452
tri 4976 436 4980 440 se
rect 4980 436 5039 440
tri 5039 436 5043 440 nw
rect 4658 392 4710 404
rect 4839 430 5009 436
rect 4658 334 4710 340
rect 4759 387 4805 399
rect 4839 396 4851 430
rect 4885 396 4923 430
rect 4957 406 5009 430
tri 5009 406 5039 436 nw
rect 5122 406 5128 440
rect 5162 406 5168 440
rect 4957 396 4998 406
rect 4839 395 4998 396
tri 4998 395 5009 406 nw
rect 4839 390 4993 395
tri 4993 390 4998 395 nw
rect 4759 353 4765 387
rect 4799 353 4805 387
rect 5122 368 5168 406
rect 4759 334 4805 353
tri 4805 334 4826 355 sw
tri 5101 334 5122 355 se
rect 5122 334 5128 368
rect 5162 334 5168 368
rect 4381 322 4433 328
rect 4759 330 4826 334
tri 4826 330 4830 334 sw
tri 5097 330 5101 334 se
rect 5101 330 5168 334
rect 4759 322 4830 330
tri 4830 322 4838 330 sw
tri 5089 322 5097 330 se
rect 5097 322 5168 330
rect 5221 444 5273 452
rect 5221 380 5273 392
rect 5221 322 5273 328
rect 5303 444 5355 452
tri 5509 451 5510 452 ne
rect 5303 380 5355 392
rect 5510 429 5556 452
rect 5510 395 5516 429
rect 5550 395 5556 429
rect 5510 383 5556 395
rect 5607 462 5653 513
tri 5653 462 5659 468 sw
rect 5607 456 5659 462
rect 5607 392 5659 404
rect 5607 334 5659 340
rect 5884 444 5936 452
rect 6050 442 6056 445
rect 5884 380 5936 392
rect 5303 322 5355 328
rect 5884 322 5936 328
rect 5972 387 6018 399
rect 6048 396 6056 442
rect 6050 393 6056 396
rect 6108 393 6120 445
rect 6172 393 6178 445
rect 6330 440 6376 452
rect 6330 406 6336 440
rect 6370 406 6376 440
rect 5972 353 5978 387
rect 6012 353 6018 387
rect 6330 368 6376 406
rect 5972 334 6018 353
tri 6018 334 6039 355 sw
tri 6309 334 6330 355 se
rect 6330 334 6336 368
rect 6370 334 6376 368
rect 3832 315 4239 321
rect 3832 281 3838 315
rect 3872 281 4239 315
rect 3832 269 4239 281
rect 4759 321 4838 322
tri 4838 321 4839 322 sw
tri 5088 321 5089 322 se
rect 5089 321 5168 322
rect 4759 315 5168 321
rect 4759 281 4765 315
rect 4799 281 5168 315
rect 4759 269 5168 281
rect 5972 321 6039 334
tri 6039 321 6052 334 sw
tri 6296 321 6309 334 se
rect 6309 321 6376 334
rect 6720 440 6766 452
rect 6720 406 6726 440
rect 6760 406 6766 440
rect 6720 368 6766 406
rect 6720 334 6726 368
rect 6760 334 6766 368
rect 6720 322 6766 334
rect 6822 440 6868 452
rect 6822 406 6828 440
rect 6862 406 6868 440
rect 6822 368 6868 406
rect 6822 334 6828 368
rect 6862 334 6868 368
rect 6822 322 6868 334
rect 5972 315 6376 321
rect 5972 281 5978 315
rect 6012 281 6376 315
rect 5972 269 6376 281
rect 66 70 6979 241
rect 66 36 78 70
rect 112 36 151 70
rect 185 36 224 70
rect 258 36 297 70
rect 331 36 370 70
rect 404 36 443 70
rect 477 36 516 70
rect 550 36 589 70
rect 623 36 662 70
rect 696 36 735 70
rect 769 36 808 70
rect 842 36 881 70
rect 915 36 954 70
rect 988 36 1027 70
rect 1061 36 1100 70
rect 1134 36 1173 70
rect 1207 36 1245 70
rect 1279 36 1317 70
rect 1351 36 1389 70
rect 1423 36 1461 70
rect 1495 36 1533 70
rect 1567 36 1605 70
rect 1639 36 1677 70
rect 1711 36 1749 70
rect 1783 36 1821 70
rect 1855 36 1893 70
rect 1927 36 1965 70
rect 1999 36 2037 70
rect 2071 36 2109 70
rect 2143 36 2181 70
rect 2215 36 2253 70
rect 2287 36 2325 70
rect 2359 36 2397 70
rect 2431 36 2469 70
rect 2503 36 2541 70
rect 2575 36 2613 70
rect 2647 36 2685 70
rect 2719 36 2757 70
rect 2791 36 2829 70
rect 2863 36 2901 70
rect 2935 36 2973 70
rect 3007 36 3045 70
rect 3079 36 3117 70
rect 3151 36 3189 70
rect 3223 36 3261 70
rect 3295 36 3333 70
rect 3367 36 3405 70
rect 3439 36 3477 70
rect 3511 36 3549 70
rect 3583 36 3621 70
rect 3655 36 3693 70
rect 3727 36 3765 70
rect 3799 36 3837 70
rect 3871 36 3909 70
rect 3943 36 3981 70
rect 4015 36 4053 70
rect 4087 36 4125 70
rect 4159 36 4197 70
rect 4231 36 4269 70
rect 4303 36 4341 70
rect 4375 36 4413 70
rect 4447 36 4485 70
rect 4519 36 4557 70
rect 4591 36 4629 70
rect 4663 36 4701 70
rect 4735 36 4773 70
rect 4807 36 4845 70
rect 4879 36 4917 70
rect 4951 36 4989 70
rect 5023 36 5061 70
rect 5095 36 5133 70
rect 5167 36 5205 70
rect 5239 36 5277 70
rect 5311 36 5349 70
rect 5383 36 5421 70
rect 5455 36 5493 70
rect 5527 36 5565 70
rect 5599 36 5637 70
rect 5671 36 5709 70
rect 5743 36 5781 70
rect 5815 36 5853 70
rect 5887 36 5925 70
rect 5959 36 5997 70
rect 6031 36 6069 70
rect 6103 36 6141 70
rect 6175 36 6213 70
rect 6247 36 6285 70
rect 6319 36 6357 70
rect 6391 36 6429 70
rect 6463 36 6501 70
rect 6535 36 6573 70
rect 6607 36 6645 70
rect 6679 36 6717 70
rect 6751 36 6789 70
rect 6823 36 6861 70
rect 6895 36 6933 70
rect 6967 36 6979 70
rect 66 26 6979 36
rect 6048 -134 6054 -82
rect 6106 -134 6118 -82
rect 6170 -134 6176 -82
<< via1 >>
rect 4664 701 4716 753
rect 4728 701 4780 753
rect 4224 621 4276 673
rect 4288 621 4340 673
rect 4439 621 4491 673
rect 4503 621 4555 673
rect 5309 621 5361 673
rect 5373 621 5425 673
rect 5856 621 5908 673
rect 5920 621 5972 673
rect 3918 541 3970 593
rect 3982 541 4034 593
rect 4658 452 4710 456
rect 3918 405 3970 414
rect 3918 371 3924 405
rect 3924 371 3958 405
rect 3958 371 3970 405
rect 3918 362 3970 371
rect 3982 405 4034 414
rect 3982 371 3996 405
rect 3996 371 4030 405
rect 4030 371 4034 405
rect 3982 362 4034 371
rect 4294 440 4346 445
rect 4294 406 4303 440
rect 4303 406 4337 440
rect 4337 406 4346 440
rect 4294 393 4346 406
rect 4294 368 4346 381
rect 4294 334 4303 368
rect 4303 334 4337 368
rect 4337 334 4346 368
rect 4294 329 4346 334
rect 4381 440 4433 444
rect 4381 406 4390 440
rect 4390 406 4424 440
rect 4424 406 4433 440
rect 4381 392 4433 406
rect 4381 368 4433 380
rect 4381 334 4390 368
rect 4390 334 4424 368
rect 4424 334 4433 368
rect 4658 418 4667 452
rect 4667 418 4701 452
rect 4701 418 4710 452
rect 4658 404 4710 418
rect 4658 380 4710 392
rect 4658 346 4667 380
rect 4667 346 4701 380
rect 4701 346 4710 380
rect 4658 340 4710 346
rect 4381 328 4433 334
rect 5221 440 5273 444
rect 5221 406 5230 440
rect 5230 406 5264 440
rect 5264 406 5273 440
rect 5221 392 5273 406
rect 5221 368 5273 380
rect 5221 334 5230 368
rect 5230 334 5264 368
rect 5264 334 5273 368
rect 5221 328 5273 334
rect 5303 440 5355 444
rect 5303 406 5312 440
rect 5312 406 5346 440
rect 5346 406 5355 440
rect 5303 392 5355 406
rect 5607 452 5659 456
rect 5607 418 5613 452
rect 5613 418 5647 452
rect 5647 418 5659 452
rect 5607 404 5659 418
rect 5303 368 5355 380
rect 5303 334 5312 368
rect 5312 334 5346 368
rect 5346 334 5355 368
rect 5607 380 5659 392
rect 5607 346 5613 380
rect 5613 346 5647 380
rect 5647 346 5659 380
rect 5607 340 5659 346
rect 5884 440 5936 444
rect 5884 406 5893 440
rect 5893 406 5927 440
rect 5927 406 5936 440
rect 5884 392 5936 406
rect 5884 368 5936 380
rect 5884 334 5893 368
rect 5893 334 5927 368
rect 5927 334 5936 368
rect 5303 328 5355 334
rect 5884 328 5936 334
rect 6056 436 6108 445
rect 6056 402 6060 436
rect 6060 402 6094 436
rect 6094 402 6108 436
rect 6056 393 6108 402
rect 6120 436 6172 445
rect 6120 402 6132 436
rect 6132 402 6166 436
rect 6166 402 6172 436
rect 6120 393 6172 402
rect 6054 -134 6106 -82
rect 6118 -134 6170 -82
<< metal2 >>
rect 4658 701 4664 753
rect 4716 701 4728 753
rect 4780 701 4786 753
rect 4658 673 4716 701
tri 4716 673 4744 701 nw
rect 4218 621 4224 673
rect 4276 621 4288 673
rect 4340 621 4346 673
tri 4260 593 4288 621 ne
rect 4288 593 4346 621
rect 3912 541 3918 593
rect 3970 541 3982 593
rect 4034 541 4040 593
tri 4288 587 4294 593 ne
rect 3912 445 3964 541
tri 3964 507 3998 541 nw
tri 3964 445 3967 448 sw
rect 4294 445 4346 593
rect 3912 414 3967 445
tri 3967 414 3998 445 sw
rect 3912 362 3918 414
rect 3970 362 3982 414
rect 4034 362 4040 414
rect 4294 381 4346 393
rect 4294 323 4346 329
rect 4381 621 4439 673
rect 4491 621 4503 673
rect 4555 621 4561 673
rect 4381 444 4433 621
tri 4433 587 4467 621 nw
rect 4381 380 4433 392
rect 4658 456 4710 673
tri 4710 667 4716 673 nw
rect 5303 621 5309 673
rect 5361 621 5373 673
rect 5425 621 5431 673
rect 5850 621 5856 673
rect 5908 621 5920 673
rect 5972 621 5978 673
rect 4658 392 4710 404
rect 4658 334 4710 340
rect 5221 444 5273 450
rect 5221 380 5273 392
rect 4381 322 4433 328
rect 5221 322 5273 328
rect 5303 444 5355 621
tri 5355 587 5389 621 nw
tri 5850 587 5884 621 ne
rect 5303 380 5355 392
rect 5607 456 5659 462
rect 5607 392 5659 404
rect 5607 334 5659 340
rect 5884 444 5936 621
tri 5936 587 5970 621 nw
rect 5884 380 5936 392
rect 5303 322 5355 328
rect 5884 322 5936 328
rect 6048 393 6056 445
rect 6108 393 6120 445
rect 6172 393 6178 445
rect 6048 -82 6100 393
tri 6100 359 6134 393 nw
tri 6100 -82 6143 -39 sw
rect 6048 -134 6054 -82
rect 6106 -134 6118 -82
rect 6170 -134 6176 -82
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_0
timestamp 1624884095
transform -1 0 5800 0 1 2
box -46 24 399 1116
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_1
timestamp 1624884095
transform 1 0 2551 0 1 2
box -46 24 399 1116
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_2
timestamp 1624884095
transform 1 0 6190 0 1 2
box -46 24 399 1116
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_3
timestamp 1624884095
transform 1 0 504 0 1 2
box -46 24 399 1116
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_4
timestamp 1624884095
transform 1 0 1714 0 1 2
box -46 24 399 1116
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_5
timestamp 1624884095
transform 1 0 3302 0 1 2
box -46 24 399 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_0
timestamp 1624884095
transform 1 0 6476 0 1 2
box -42 24 569 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_1
timestamp 1624884095
transform 1 0 1252 0 1 2
box -42 24 569 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_2
timestamp 1624884095
transform 1 0 42 0 1 2
box -42 24 569 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_3
timestamp 1624884095
transform -1 0 5514 0 1 2
box -42 24 569 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_4
timestamp 1624884095
transform -1 0 4587 0 1 2
box -42 24 569 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_5
timestamp 1624884095
transform -1 0 1324 0 1 2
box -42 24 569 1116
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_6
timestamp 1624884095
transform 1 0 5728 0 1 2
box -42 24 569 1116
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_0
timestamp 1624884095
transform 1 0 3588 0 1 2
box 0 24 534 1116
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_1
timestamp 1624884095
transform 1 0 4515 0 1 2
box 0 24 534 1116
use sky130_fd_io__hvsbt_nor  sky130_fd_io__hvsbt_nor_2
timestamp 1624884095
transform 1 0 2837 0 1 2
box 0 24 534 1116
<< labels >>
flabel metal1 s 370 401 484 436 3 FreeSans 200 0 0 0 DM_H_N[0]
port 1 nsew
flabel metal1 s 137 405 237 435 3 FreeSans 100 0 0 0 DM_H_N[1]
port 2 nsew
flabel metal1 s 1592 403 1689 435 3 FreeSans 100 0 0 0 INP_DIS_H_N
port 3 nsew
flabel metal1 s 1871 366 1900 434 3 FreeSans 100 90 0 0 INP_DIS_I_H
port 4 nsew
flabel metal1 s 1968 381 1992 460 3 FreeSans 100 0 0 0 INP_DIS_I_H_N
port 5 nsew
flabel metal1 s 2710 350 2734 419 3 FreeSans 100 90 0 0 VTRIP_SEL_H
port 6 nsew
flabel metal1 s 3449 350 3476 443 3 FreeSans 100 0 0 0 TRIPSEL_I_H
port 7 nsew
flabel metal1 s 3561 350 3588 444 3 FreeSans 100 0 0 0 TRIPSEL_I_H_N
port 8 nsew
flabel metal1 s 3741 364 3768 472 3 FreeSans 100 0 0 0 IBUF_MODE_SEL[1]
port 9 nsew
flabel metal1 s 3941 376 4023 407 3 FreeSans 100 0 0 0 IBUF_MODE_SEL[0]
port 10 nsew
flabel metal1 s 5232 347 5266 432 3 FreeSans 100 0 0 0 MODE_VCCD_N
port 11 nsew
flabel metal1 s 6334 359 6365 436 3 FreeSans 100 0 0 0 MODE_REF_N
port 12 nsew
flabel metal1 s 6831 342 6858 433 3 FreeSans 100 0 0 0 HYS_TRIM
port 13 nsew
flabel metal1 s 6724 344 6759 442 3 FreeSans 100 0 0 0 MODE_REF_3V_N
port 14 nsew
flabel metal1 s 1137 405 1215 431 3 FreeSans 100 0 0 0 DM_H_N[2]
port 15 nsew
flabel metal1 s 4309 345 4337 439 3 FreeSans 100 0 0 0 MODE_NORMAL_N
port 16 nsew
flabel metal1 s 102 885 445 1044 3 FreeSans 100 0 0 0 VDDIO_Q
port 17 nsew
flabel metal1 s 106 46 259 205 3 FreeSans 100 0 0 0 VSSD
port 18 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 36563994
string GDS_START 36516372
<< end >>
