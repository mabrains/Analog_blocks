**.subckt untitled-11
XM12 inn mir VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM2 inp mir VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM3 bg_out mir VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XQ2 GND GND net3 sky130_fd_pr__pnp_05v5_W0p68L0p68
XQ3 GND GND net1 sky130_fd_pr__pnp_05v5_W0p68L0p68
XQ4 GND GND net1 sky130_fd_pr__pnp_05v5_W0p68L0p68
XQ8 GND GND net1 sky130_fd_pr__pnp_05v5_W0p68L0p68
XQ10 GND GND net1 sky130_fd_pr__pnp_05v5_W0p68L0p68
XQ12 GND GND net1 sky130_fd_pr__pnp_05v5_W0p68L0p68
XQ14 GND GND net1 sky130_fd_pr__pnp_05v5_W0p68L0p68
XQ16 GND GND net1 sky130_fd_pr__pnp_05v5_W0p68L0p68
XQ18 GND GND net1 sky130_fd_pr__pnp_05v5_W0p68L0p68
XM15 net2 bg_out GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=8 m=8 
XM16 VDD net2 inn GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM17 net2 bg_out VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=5 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2 
XM4 net5 net5 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM19 net5 inp net4 GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM1 mir inn net4 GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM7 mir net5 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM22 net4 net6 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM8 net6 mir VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM6 net6 net6 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XC1 mir GND sky130_fd_pr__cap_mim_m3_1 W=14 L=14 MF=1 m=1
XR7 GND bg_out GND sky130_fd_pr__res_xhigh_po_0p35 L=14.5 mult=1 m=1
XR6 GND net7 GND sky130_fd_pr__res_xhigh_po_0p35 L=15.2 mult=1 m=1
XR4 GND net3 GND sky130_fd_pr__res_xhigh_po_0p35 L=15.2 mult=1 m=1
XR2 net1 net7 GND sky130_fd_pr__res_xhigh_po_0p35 L=2.3 mult=1 m=1
XR1 net7 inp GND sky130_fd_pr__res_xhigh_po_0p35 L=5 mult=1 m=1
XR3 net3 inn GND sky130_fd_pr__res_xhigh_po_0p35 L=5 mult=1 m=1
XM5 net9 net9 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1.2 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM9 net9 bg_out net10 GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=8 m=8 
XM10 net8 pos net10 GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM11 net8 net9 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1.2 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM13 net10 vb GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
Vs VDD GND 2.2
XM14 out net8 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1.2 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=12 m=12 
XM18 out vb GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=12 m=12 
XM20 vb vb GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM21 bp vb GND GND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM23 bp bp VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=1.2 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM24 ldo_out out VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=800 m=800 
C2 net8 net11 8p m=1
R9 out net11 10k m=1
XM26 vb mir VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XR10 pos ldo_out GND sky130_fd_pr__res_xhigh_po_0p35 L=5.5 mult=1 m=1
XR11 GND pos GND sky130_fd_pr__res_xhigh_po_0p35 L=9 mult=1 m=1
**** begin user architecture code


.lib /home/mustafa/mabrains/pdks/share/pdk/sky130A/libs.tech/ngspice/sky130.lib_mod.spice fs_hh

.nodeset v(inn)=1.1
.nodeset v(inp)=1.1
.nodeset v(mir)=0.9
.nodeset v(bg_out)=1.2
.nodeset v(ldo_out)=1.8
.nodeset v(pos)=1.2

.control
op
print all
.endc

.control

dc Vs 2.5 0 -0.02
plot vdd ldo_out
meas DC Vref_Sup_pos10per FIND bg_out AT=2
meas DC Vref_Sup_neg10per FIND bg_out AT=2.4
.endc

*Temprature Variation
.control
let i=16
dc temp 85 0 -1
set appendwrite
write temp_var_ldo.raw
load temp_var_ldo.raw
plot v (ldo_out)
.endc




.control
alter Vs AC =1
ac dec 10 1 1G
plot vdb (ldo_out)
let psrr = vdb(ldo_out)
meas ac PSRR_1k FIND vdb(ldo_out) AT=1k
meas ac PSRR_1M FIND vdb(ldo_out) AT=100k
set appendwrite
write psrr_ldo.raw
load psrr_ldo.raw
quit
.endc







**Transient
*.control
*alter @Vs[pulse] = [ 0 2 15u 1u 5u 100u 200u ]
*tran 0.1u 100u
*plot vdd ldo_out
*.endc
*.control
*alter @Vs[pulse] = [ 0 2.2 15u 1u 5u 100u 200u ]
*tran 0.1u 100u
*plot vdd ldo_out
*.endc
*.control
*alter @Vs[pulse] = [ 0 2.4 15u 1u 5u 100u 200u ]
*tran 0.1u 100u
*plot vdd ldo_out
*.endc





**** end user architecture code
**.ends
.GLOBAL VDD
.GLOBAL GND
** flattened .save nodes
.end
