magic
tech sky130A
magscale 1 2
timestamp 1624884095
<< checkpaint >>
rect -69 -220 3205 4407
<< nwell >>
rect 1191 2415 1685 3147
<< pwell >>
rect 1240 1958 1508 1968
rect 1240 1306 1945 1958
rect 1240 1159 1508 1306
<< mvnmos >>
rect 1610 1332 1710 1932
rect 1766 1332 1866 1932
<< mvpmos >>
rect 1310 2481 1410 3081
rect 1466 2481 1566 3081
<< mvndiff >>
rect 1557 1854 1610 1932
rect 1557 1820 1565 1854
rect 1599 1820 1610 1854
rect 1557 1786 1610 1820
rect 1557 1752 1565 1786
rect 1599 1752 1610 1786
rect 1557 1718 1610 1752
rect 1557 1684 1565 1718
rect 1599 1684 1610 1718
rect 1557 1650 1610 1684
rect 1557 1616 1565 1650
rect 1599 1616 1610 1650
rect 1557 1582 1610 1616
rect 1557 1548 1565 1582
rect 1599 1548 1610 1582
rect 1557 1514 1610 1548
rect 1557 1480 1565 1514
rect 1599 1480 1610 1514
rect 1557 1446 1610 1480
rect 1557 1412 1565 1446
rect 1599 1412 1610 1446
rect 1557 1378 1610 1412
rect 1557 1344 1565 1378
rect 1599 1344 1610 1378
rect 1557 1332 1610 1344
rect 1710 1854 1766 1932
rect 1710 1820 1721 1854
rect 1755 1820 1766 1854
rect 1710 1786 1766 1820
rect 1710 1752 1721 1786
rect 1755 1752 1766 1786
rect 1710 1718 1766 1752
rect 1710 1684 1721 1718
rect 1755 1684 1766 1718
rect 1710 1650 1766 1684
rect 1710 1616 1721 1650
rect 1755 1616 1766 1650
rect 1710 1582 1766 1616
rect 1710 1548 1721 1582
rect 1755 1548 1766 1582
rect 1710 1514 1766 1548
rect 1710 1480 1721 1514
rect 1755 1480 1766 1514
rect 1710 1446 1766 1480
rect 1710 1412 1721 1446
rect 1755 1412 1766 1446
rect 1710 1378 1766 1412
rect 1710 1344 1721 1378
rect 1755 1344 1766 1378
rect 1710 1332 1766 1344
rect 1866 1854 1919 1932
rect 1866 1820 1877 1854
rect 1911 1820 1919 1854
rect 1866 1786 1919 1820
rect 1866 1752 1877 1786
rect 1911 1752 1919 1786
rect 1866 1718 1919 1752
rect 1866 1684 1877 1718
rect 1911 1684 1919 1718
rect 1866 1650 1919 1684
rect 1866 1616 1877 1650
rect 1911 1616 1919 1650
rect 1866 1582 1919 1616
rect 1866 1548 1877 1582
rect 1911 1548 1919 1582
rect 1866 1514 1919 1548
rect 1866 1480 1877 1514
rect 1911 1480 1919 1514
rect 1866 1446 1919 1480
rect 1866 1412 1877 1446
rect 1911 1412 1919 1446
rect 1866 1378 1919 1412
rect 1866 1344 1877 1378
rect 1911 1344 1919 1378
rect 1866 1332 1919 1344
<< mvpdiff >>
rect 1257 3003 1310 3081
rect 1257 2969 1265 3003
rect 1299 2969 1310 3003
rect 1257 2935 1310 2969
rect 1257 2901 1265 2935
rect 1299 2901 1310 2935
rect 1257 2867 1310 2901
rect 1257 2833 1265 2867
rect 1299 2833 1310 2867
rect 1257 2799 1310 2833
rect 1257 2765 1265 2799
rect 1299 2765 1310 2799
rect 1257 2731 1310 2765
rect 1257 2697 1265 2731
rect 1299 2697 1310 2731
rect 1257 2663 1310 2697
rect 1257 2629 1265 2663
rect 1299 2629 1310 2663
rect 1257 2595 1310 2629
rect 1257 2561 1265 2595
rect 1299 2561 1310 2595
rect 1257 2527 1310 2561
rect 1257 2493 1265 2527
rect 1299 2493 1310 2527
rect 1257 2481 1310 2493
rect 1410 3003 1466 3081
rect 1410 2969 1421 3003
rect 1455 2969 1466 3003
rect 1410 2935 1466 2969
rect 1410 2901 1421 2935
rect 1455 2901 1466 2935
rect 1410 2867 1466 2901
rect 1410 2833 1421 2867
rect 1455 2833 1466 2867
rect 1410 2799 1466 2833
rect 1410 2765 1421 2799
rect 1455 2765 1466 2799
rect 1410 2731 1466 2765
rect 1410 2697 1421 2731
rect 1455 2697 1466 2731
rect 1410 2663 1466 2697
rect 1410 2629 1421 2663
rect 1455 2629 1466 2663
rect 1410 2595 1466 2629
rect 1410 2561 1421 2595
rect 1455 2561 1466 2595
rect 1410 2527 1466 2561
rect 1410 2493 1421 2527
rect 1455 2493 1466 2527
rect 1410 2481 1466 2493
rect 1566 3003 1619 3081
rect 1566 2969 1577 3003
rect 1611 2969 1619 3003
rect 1566 2935 1619 2969
rect 1566 2901 1577 2935
rect 1611 2901 1619 2935
rect 1566 2867 1619 2901
rect 1566 2833 1577 2867
rect 1611 2833 1619 2867
rect 1566 2799 1619 2833
rect 1566 2765 1577 2799
rect 1611 2765 1619 2799
rect 1566 2731 1619 2765
rect 1566 2697 1577 2731
rect 1611 2697 1619 2731
rect 1566 2663 1619 2697
rect 1566 2629 1577 2663
rect 1611 2629 1619 2663
rect 1566 2595 1619 2629
rect 1566 2561 1577 2595
rect 1611 2561 1619 2595
rect 1566 2527 1619 2561
rect 1566 2493 1577 2527
rect 1611 2493 1619 2527
rect 1566 2481 1619 2493
<< mvndiffc >>
rect 1565 1820 1599 1854
rect 1565 1752 1599 1786
rect 1565 1684 1599 1718
rect 1565 1616 1599 1650
rect 1565 1548 1599 1582
rect 1565 1480 1599 1514
rect 1565 1412 1599 1446
rect 1565 1344 1599 1378
rect 1721 1820 1755 1854
rect 1721 1752 1755 1786
rect 1721 1684 1755 1718
rect 1721 1616 1755 1650
rect 1721 1548 1755 1582
rect 1721 1480 1755 1514
rect 1721 1412 1755 1446
rect 1721 1344 1755 1378
rect 1877 1820 1911 1854
rect 1877 1752 1911 1786
rect 1877 1684 1911 1718
rect 1877 1616 1911 1650
rect 1877 1548 1911 1582
rect 1877 1480 1911 1514
rect 1877 1412 1911 1446
rect 1877 1344 1911 1378
<< mvpdiffc >>
rect 1265 2969 1299 3003
rect 1265 2901 1299 2935
rect 1265 2833 1299 2867
rect 1265 2765 1299 2799
rect 1265 2697 1299 2731
rect 1265 2629 1299 2663
rect 1265 2561 1299 2595
rect 1265 2493 1299 2527
rect 1421 2969 1455 3003
rect 1421 2901 1455 2935
rect 1421 2833 1455 2867
rect 1421 2765 1455 2799
rect 1421 2697 1455 2731
rect 1421 2629 1455 2663
rect 1421 2561 1455 2595
rect 1421 2493 1455 2527
rect 1577 2969 1611 3003
rect 1577 2901 1611 2935
rect 1577 2833 1611 2867
rect 1577 2765 1611 2799
rect 1577 2697 1611 2731
rect 1577 2629 1611 2663
rect 1577 2561 1611 2595
rect 1577 2493 1611 2527
<< psubdiff >>
rect 1266 1918 1482 1942
rect 1266 1884 1267 1918
rect 1301 1884 1357 1918
rect 1391 1884 1447 1918
rect 1481 1884 1482 1918
rect 1266 1806 1482 1884
rect 1266 1772 1267 1806
rect 1301 1772 1357 1806
rect 1391 1772 1447 1806
rect 1481 1772 1482 1806
rect 1266 1694 1482 1772
rect 1266 1660 1267 1694
rect 1301 1660 1357 1694
rect 1391 1660 1447 1694
rect 1481 1660 1482 1694
rect 1266 1582 1482 1660
rect 1266 1548 1267 1582
rect 1301 1548 1357 1582
rect 1391 1548 1447 1582
rect 1481 1548 1482 1582
rect 1266 1469 1482 1548
rect 1266 1435 1267 1469
rect 1301 1435 1357 1469
rect 1391 1435 1447 1469
rect 1481 1435 1482 1469
rect 1266 1356 1482 1435
rect 1266 1322 1267 1356
rect 1301 1322 1357 1356
rect 1391 1322 1447 1356
rect 1481 1322 1482 1356
rect 1266 1243 1482 1322
rect 1266 1209 1267 1243
rect 1301 1209 1357 1243
rect 1391 1209 1447 1243
rect 1481 1209 1482 1243
rect 1266 1185 1482 1209
<< psubdiffcont >>
rect 1267 1884 1301 1918
rect 1357 1884 1391 1918
rect 1447 1884 1481 1918
rect 1267 1772 1301 1806
rect 1357 1772 1391 1806
rect 1447 1772 1481 1806
rect 1267 1660 1301 1694
rect 1357 1660 1391 1694
rect 1447 1660 1481 1694
rect 1267 1548 1301 1582
rect 1357 1548 1391 1582
rect 1447 1548 1481 1582
rect 1267 1435 1301 1469
rect 1357 1435 1391 1469
rect 1447 1435 1481 1469
rect 1267 1322 1301 1356
rect 1357 1322 1391 1356
rect 1447 1322 1481 1356
rect 1267 1209 1301 1243
rect 1357 1209 1391 1243
rect 1447 1209 1481 1243
<< poly >>
rect 1310 3081 1410 3113
rect 1466 3081 1566 3113
rect 1310 2449 1410 2481
rect 1276 2433 1410 2449
rect 1276 2399 1292 2433
rect 1326 2399 1360 2433
rect 1394 2399 1410 2433
rect 1276 2383 1410 2399
rect 1466 2449 1566 2481
rect 1466 2433 1600 2449
rect 1466 2399 1482 2433
rect 1516 2399 1550 2433
rect 1584 2399 1600 2433
rect 1466 2383 1600 2399
rect 1576 2014 1710 2030
rect 1576 1980 1592 2014
rect 1626 1980 1660 2014
rect 1694 1980 1710 2014
rect 1576 1964 1710 1980
rect 1610 1932 1710 1964
rect 1766 2014 1900 2030
rect 1766 1980 1782 2014
rect 1816 1980 1850 2014
rect 1884 1980 1900 2014
rect 1766 1964 1900 1980
rect 1766 1932 1866 1964
rect 1610 1300 1710 1332
rect 1766 1300 1866 1332
<< polycont >>
rect 1292 2399 1326 2433
rect 1360 2399 1394 2433
rect 1482 2399 1516 2433
rect 1550 2399 1584 2433
rect 1592 1980 1626 2014
rect 1660 1980 1694 2014
rect 1782 1980 1816 2014
rect 1850 1980 1884 2014
<< locali >>
rect 1265 3003 1299 3019
rect 1265 2935 1299 2969
rect 1265 2867 1299 2901
rect 1265 2799 1299 2833
rect 1265 2731 1299 2765
rect 1265 2685 1299 2697
rect 1265 2604 1299 2629
rect 1265 2527 1299 2561
rect 1421 3003 1455 3019
rect 1421 2935 1455 2969
rect 1421 2867 1455 2901
rect 1421 2799 1455 2833
rect 1421 2731 1455 2765
rect 1421 2663 1455 2697
rect 1421 2626 1455 2629
rect 1421 2554 1455 2561
rect 1265 2477 1299 2489
rect 1577 3003 1611 3019
rect 1577 2935 1611 2969
rect 1577 2867 1611 2901
rect 1577 2799 1611 2833
rect 1577 2731 1611 2765
rect 1577 2663 1611 2697
rect 1577 2604 1611 2629
rect 1577 2532 1611 2561
rect 1421 2477 1455 2493
rect 1343 2438 1377 2476
rect 1577 2477 1611 2493
rect 1502 2438 1536 2476
rect 1276 2399 1292 2433
rect 1326 2404 1343 2433
rect 1326 2399 1360 2404
rect 1394 2399 1410 2433
rect 1466 2399 1482 2433
rect 1536 2404 1550 2433
rect 1516 2399 1550 2404
rect 1584 2399 1600 2433
rect 1588 2014 1622 2052
rect 1803 2014 1837 2021
rect 1576 1980 1588 2014
rect 1626 1980 1660 2014
rect 1694 1980 1710 2014
rect 1766 1980 1782 2014
rect 1816 1983 1850 2014
rect 1837 1980 1850 1983
rect 1884 1980 1900 2014
rect 1266 1918 1482 1942
rect 1266 1884 1267 1918
rect 1301 1884 1357 1918
rect 1391 1884 1447 1918
rect 1481 1884 1482 1918
rect 1266 1806 1482 1884
rect 1266 1772 1267 1806
rect 1301 1772 1357 1806
rect 1391 1772 1447 1806
rect 1481 1772 1482 1806
rect 1266 1694 1482 1772
rect 1266 1660 1267 1694
rect 1301 1660 1357 1694
rect 1391 1660 1447 1694
rect 1481 1660 1482 1694
rect 1266 1651 1482 1660
rect 1266 1617 1275 1651
rect 1309 1617 1393 1651
rect 1427 1617 1482 1651
rect 1266 1582 1482 1617
rect 1266 1548 1267 1582
rect 1301 1567 1357 1582
rect 1309 1548 1357 1567
rect 1391 1567 1447 1582
rect 1391 1548 1393 1567
rect 1266 1533 1275 1548
rect 1309 1533 1393 1548
rect 1427 1548 1447 1567
rect 1481 1548 1482 1582
rect 1427 1533 1482 1548
rect 1266 1483 1482 1533
rect 1266 1469 1275 1483
rect 1309 1469 1393 1483
rect 1266 1435 1267 1469
rect 1309 1449 1357 1469
rect 1301 1435 1357 1449
rect 1391 1449 1393 1469
rect 1427 1469 1482 1483
rect 1427 1449 1447 1469
rect 1391 1435 1447 1449
rect 1481 1435 1482 1469
rect 1266 1398 1482 1435
rect 1266 1364 1275 1398
rect 1309 1364 1393 1398
rect 1427 1364 1482 1398
rect 1266 1356 1482 1364
rect 1266 1322 1267 1356
rect 1301 1322 1357 1356
rect 1391 1322 1447 1356
rect 1481 1322 1482 1356
rect 1565 1854 1577 1880
rect 1599 1820 1611 1846
rect 1565 1808 1611 1820
rect 1565 1786 1577 1808
rect 1721 1854 1755 1868
rect 1721 1786 1755 1796
rect 1565 1718 1599 1752
rect 1565 1650 1599 1684
rect 1565 1582 1599 1616
rect 1565 1514 1599 1548
rect 1565 1446 1599 1480
rect 1565 1378 1599 1412
rect 1565 1328 1599 1344
rect 1721 1718 1755 1752
rect 1721 1650 1755 1684
rect 1721 1582 1755 1616
rect 1721 1514 1755 1548
rect 1721 1446 1755 1480
rect 1721 1378 1755 1412
rect 1721 1328 1755 1344
rect 1877 1854 1911 1860
rect 1877 1786 1911 1788
rect 1877 1718 1911 1752
rect 1877 1650 1911 1684
rect 1877 1582 1911 1616
rect 1877 1514 1911 1548
rect 1877 1446 1911 1480
rect 1877 1378 1911 1412
rect 1877 1328 1911 1344
rect 1266 1313 1482 1322
rect 1266 1279 1275 1313
rect 1309 1279 1393 1313
rect 1427 1279 1482 1313
rect 1266 1243 1482 1279
rect 1266 1209 1267 1243
rect 1301 1228 1357 1243
rect 1309 1209 1357 1228
rect 1391 1228 1447 1243
rect 1391 1209 1393 1228
rect 1266 1194 1275 1209
rect 1309 1194 1393 1209
rect 1427 1209 1447 1228
rect 1481 1209 1482 1243
rect 1427 1194 1482 1209
rect 1266 1185 1482 1194
<< viali >>
rect 1265 2663 1299 2685
rect 1265 2651 1299 2663
rect 1265 2595 1299 2604
rect 1265 2570 1299 2595
rect 1265 2493 1299 2523
rect 1421 2595 1455 2626
rect 1421 2592 1455 2595
rect 1421 2527 1455 2554
rect 1421 2520 1455 2527
rect 1265 2489 1299 2493
rect 1343 2476 1377 2510
rect 1577 2595 1611 2604
rect 1577 2570 1611 2595
rect 1577 2527 1611 2532
rect 1343 2433 1377 2438
rect 1502 2476 1536 2510
rect 1577 2498 1611 2527
rect 1502 2433 1536 2438
rect 1343 2404 1360 2433
rect 1360 2404 1377 2433
rect 1502 2404 1516 2433
rect 1516 2404 1536 2433
rect 1588 2052 1622 2086
rect 1803 2021 1837 2055
rect 1588 1980 1592 2014
rect 1592 1980 1622 2014
rect 1803 1980 1816 1983
rect 1816 1980 1837 1983
rect 1803 1949 1837 1980
rect 1275 1617 1309 1651
rect 1393 1617 1427 1651
rect 1275 1548 1301 1567
rect 1301 1548 1309 1567
rect 1275 1533 1309 1548
rect 1393 1533 1427 1567
rect 1275 1469 1309 1483
rect 1275 1449 1301 1469
rect 1301 1449 1309 1469
rect 1393 1449 1427 1483
rect 1275 1364 1309 1398
rect 1393 1364 1427 1398
rect 1577 1854 1611 1880
rect 1577 1846 1599 1854
rect 1599 1846 1611 1854
rect 1577 1786 1611 1808
rect 1577 1774 1599 1786
rect 1599 1774 1611 1786
rect 1721 1868 1755 1902
rect 1721 1820 1755 1830
rect 1721 1796 1755 1820
rect 1877 1860 1911 1894
rect 1877 1820 1911 1822
rect 1877 1788 1911 1820
rect 1275 1279 1309 1313
rect 1393 1279 1427 1313
rect 1275 1209 1301 1228
rect 1301 1209 1309 1228
rect 1275 1194 1309 1209
rect 1393 1194 1427 1228
<< metal1 >>
rect 1259 2685 1305 2697
rect 1259 2651 1265 2685
rect 1299 2651 1305 2685
rect 1259 2604 1305 2651
rect 1259 2570 1265 2604
rect 1299 2570 1305 2604
rect 1259 2523 1305 2570
rect 1259 2489 1265 2523
rect 1299 2489 1305 2523
rect 1415 2626 1461 2638
rect 1415 2592 1421 2626
rect 1455 2592 1461 2626
rect 1415 2554 1461 2592
rect 1259 2111 1305 2489
rect 1337 2510 1383 2522
rect 1337 2476 1343 2510
rect 1377 2476 1383 2510
rect 1337 2438 1383 2476
rect 1337 2404 1343 2438
rect 1377 2404 1383 2438
rect 1337 2218 1383 2404
rect 1415 2520 1421 2554
rect 1455 2520 1461 2554
rect 1571 2604 1623 2616
rect 1571 2570 1577 2604
rect 1611 2570 1623 2604
rect 1571 2532 1623 2570
rect 1415 2246 1461 2520
rect 1496 2510 1542 2522
rect 1496 2476 1502 2510
rect 1536 2476 1542 2510
rect 1496 2438 1542 2476
rect 1496 2404 1502 2438
rect 1536 2404 1542 2438
rect 1496 2281 1542 2404
rect 1571 2498 1577 2532
rect 1611 2498 1623 2532
rect 1571 2441 1623 2498
rect 1571 2377 1623 2389
rect 1571 2319 1623 2325
tri 1542 2281 1557 2296 sw
rect 1496 2268 1557 2281
tri 1557 2268 1570 2281 sw
tri 1496 2263 1501 2268 ne
rect 1501 2263 1570 2268
tri 1415 2242 1419 2246 ne
rect 1419 2242 1461 2246
tri 1461 2242 1482 2263 sw
tri 1501 2242 1522 2263 ne
rect 1522 2253 1570 2263
tri 1570 2253 1585 2268 sw
rect 1522 2242 1761 2253
tri 1419 2237 1424 2242 ne
rect 1424 2237 1482 2242
tri 1383 2218 1402 2237 sw
tri 1424 2218 1443 2237 ne
rect 1443 2228 1482 2237
tri 1482 2228 1496 2242 sw
tri 1522 2228 1536 2242 ne
rect 1536 2228 1761 2242
rect 1443 2218 1496 2228
rect 1337 2217 1402 2218
tri 1337 2177 1377 2217 ne
rect 1377 2200 1402 2217
tri 1402 2200 1420 2218 sw
tri 1443 2200 1461 2218 ne
rect 1461 2207 1496 2218
tri 1496 2207 1517 2228 sw
tri 1536 2207 1557 2228 ne
rect 1557 2217 1761 2228
tri 1761 2217 1797 2253 sw
rect 1557 2207 1797 2217
tri 1797 2207 1807 2217 sw
rect 1461 2200 1517 2207
rect 1377 2179 1420 2200
tri 1420 2179 1441 2200 sw
tri 1461 2179 1482 2200 ne
rect 1482 2179 1517 2200
tri 1517 2179 1545 2207 sw
tri 1741 2179 1769 2207 ne
rect 1769 2179 1807 2207
rect 1377 2178 1441 2179
tri 1441 2178 1442 2179 sw
tri 1482 2178 1483 2179 ne
rect 1483 2178 1694 2179
tri 1694 2178 1695 2179 sw
tri 1769 2178 1770 2179 ne
rect 1770 2178 1807 2179
rect 1377 2177 1442 2178
tri 1442 2177 1443 2178 sw
tri 1483 2177 1484 2178 ne
rect 1484 2177 1695 2178
tri 1377 2171 1383 2177 ne
rect 1383 2171 1443 2177
tri 1383 2112 1442 2171 ne
rect 1442 2152 1443 2171
tri 1443 2152 1468 2177 sw
tri 1484 2152 1509 2177 ne
rect 1509 2152 1695 2177
rect 1442 2139 1468 2152
tri 1468 2139 1481 2152 sw
tri 1509 2139 1522 2152 ne
rect 1522 2151 1695 2152
tri 1695 2151 1722 2178 sw
tri 1770 2151 1797 2178 ne
rect 1797 2171 1807 2178
tri 1807 2171 1843 2207 sw
rect 1522 2139 1722 2151
rect 1442 2112 1481 2139
tri 1481 2112 1508 2139 sw
tri 1668 2112 1695 2139 ne
rect 1695 2112 1722 2139
tri 1722 2112 1761 2151 sw
tri 1305 2111 1306 2112 sw
tri 1442 2111 1443 2112 ne
rect 1443 2111 1508 2112
tri 1508 2111 1509 2112 sw
tri 1695 2111 1696 2112 ne
rect 1696 2111 1761 2112
rect 1259 2097 1306 2111
tri 1306 2097 1320 2111 sw
tri 1443 2097 1457 2111 ne
rect 1457 2098 1575 2111
tri 1575 2098 1588 2111 sw
tri 1696 2098 1709 2111 ne
rect 1709 2098 1761 2111
rect 1457 2097 1628 2098
rect 1259 2092 1320 2097
tri 1259 2086 1265 2092 ne
rect 1265 2086 1320 2092
tri 1320 2086 1331 2097 sw
tri 1457 2086 1468 2097 ne
rect 1468 2086 1628 2097
tri 1709 2092 1715 2098 ne
tri 1265 2052 1299 2086 ne
rect 1299 2065 1331 2086
tri 1331 2065 1352 2086 sw
tri 1468 2065 1489 2086 ne
rect 1489 2065 1588 2086
rect 1299 2058 1352 2065
tri 1352 2058 1359 2065 sw
tri 1555 2058 1562 2065 ne
rect 1562 2058 1588 2065
rect 1299 2052 1359 2058
tri 1359 2052 1365 2058 sw
tri 1562 2052 1568 2058 ne
rect 1568 2052 1588 2058
rect 1622 2052 1628 2086
tri 1299 2031 1320 2052 ne
rect 1320 2045 1365 2052
tri 1365 2045 1372 2052 sw
tri 1568 2045 1575 2052 ne
rect 1575 2045 1628 2052
rect 1320 2038 1372 2045
tri 1372 2038 1379 2045 sw
tri 1575 2038 1582 2045 ne
rect 1320 2031 1379 2038
tri 1379 2031 1386 2038 sw
tri 1320 2021 1330 2031 ne
rect 1330 2021 1386 2031
tri 1386 2021 1396 2031 sw
tri 1330 2014 1337 2021 ne
rect 1337 2014 1396 2021
tri 1396 2014 1403 2021 sw
rect 1582 2014 1628 2045
tri 1337 1980 1371 2014 ne
rect 1371 1980 1403 2014
tri 1403 1980 1437 2014 sw
rect 1582 1980 1588 2014
rect 1622 1980 1628 2014
tri 1371 1965 1386 1980 ne
rect 1386 1968 1437 1980
tri 1437 1968 1449 1980 sw
rect 1582 1968 1628 1980
rect 1386 1965 1449 1968
tri 1449 1965 1452 1968 sw
tri 1386 1949 1402 1965 ne
rect 1402 1949 1452 1965
tri 1452 1949 1468 1965 sw
tri 1402 1902 1449 1949 ne
rect 1449 1902 1468 1949
tri 1468 1902 1515 1949 sw
rect 1715 1902 1761 2098
rect 1797 2055 1843 2171
rect 1797 2021 1803 2055
rect 1837 2021 1843 2055
rect 1797 1983 1843 2021
rect 1797 1949 1803 1983
rect 1837 1949 1843 1983
rect 1797 1937 1843 1949
tri 1449 1899 1452 1902 ne
rect 1452 1899 1515 1902
tri 1515 1899 1518 1902 sw
tri 1452 1885 1466 1899 ne
rect 1466 1774 1518 1899
rect 1571 1886 1623 1892
rect 1571 1820 1623 1834
tri 1518 1774 1519 1775 sw
rect 1715 1868 1721 1902
rect 1755 1868 1761 1902
rect 1715 1830 1761 1868
rect 1715 1796 1721 1830
rect 1755 1796 1761 1830
rect 1715 1784 1761 1796
rect 1871 1894 1917 1906
rect 1871 1860 1877 1894
rect 1911 1860 1917 1894
rect 1871 1822 1917 1860
tri 1865 1788 1871 1794 se
rect 1871 1788 1877 1822
rect 1911 1788 1917 1822
tri 1861 1784 1865 1788 se
rect 1865 1784 1917 1788
rect 1466 1768 1519 1774
tri 1466 1730 1504 1768 ne
rect 1504 1730 1519 1768
tri 1519 1730 1563 1774 sw
rect 1571 1762 1623 1768
tri 1839 1762 1861 1784 se
rect 1861 1774 1917 1784
rect 1861 1762 1873 1774
tri 1807 1730 1839 1762 se
rect 1839 1730 1873 1762
tri 1873 1730 1917 1774 nw
tri 1504 1716 1518 1730 ne
rect 1518 1716 1859 1730
tri 1859 1716 1873 1730 nw
tri 1518 1684 1550 1716 ne
rect 1550 1684 1827 1716
tri 1827 1684 1859 1716 nw
rect 1267 1655 1433 1663
tri 1433 1655 1441 1663 sw
rect 1267 1651 1441 1655
rect 1267 1617 1275 1651
rect 1309 1617 1393 1651
rect 1427 1617 1441 1651
rect 1267 1567 1441 1617
rect 1267 1533 1275 1567
rect 1309 1533 1393 1567
rect 1427 1533 1441 1567
rect 1267 1483 1441 1533
rect 1267 1449 1275 1483
rect 1309 1449 1393 1483
rect 1427 1449 1441 1483
rect 1267 1398 1441 1449
rect 1267 1364 1275 1398
rect 1309 1364 1393 1398
rect 1427 1364 1441 1398
rect 1267 1313 1441 1364
rect 1267 1279 1275 1313
rect 1309 1279 1393 1313
rect 1427 1279 1441 1313
rect 1267 1242 1441 1279
tri 1441 1242 1612 1413 sw
rect 1267 1228 1627 1242
rect 1267 1194 1275 1228
rect 1309 1194 1393 1228
rect 1427 1194 1627 1228
rect 1267 1040 1627 1194
<< via1 >>
rect 1571 2389 1623 2441
rect 1571 2325 1623 2377
rect 1571 1880 1623 1886
rect 1571 1846 1577 1880
rect 1577 1846 1611 1880
rect 1611 1846 1623 1880
rect 1571 1834 1623 1846
rect 1571 1808 1623 1820
rect 1571 1774 1577 1808
rect 1577 1774 1611 1808
rect 1611 1774 1623 1808
rect 1571 1768 1623 1774
<< metal2 >>
rect 1571 2441 1623 2447
rect 1571 2377 1623 2389
rect 1571 1886 1623 2325
rect 1571 1820 1623 1834
rect 1571 1762 1623 1768
use sky130_fd_pr__nfet_01v8__example_5595914180888  sky130_fd_pr__nfet_01v8__example_5595914180888_0
timestamp 1624884095
transform 1 0 1766 0 1 1332
box -28 0 128 267
use sky130_fd_pr__nfet_01v8__example_5595914180888  sky130_fd_pr__nfet_01v8__example_5595914180888_1
timestamp 1624884095
transform -1 0 1710 0 1 1332
box -28 0 128 267
use sky130_fd_pr__pfet_01v8__example_55959141808628  sky130_fd_pr__pfet_01v8__example_55959141808628_0
timestamp 1624884095
transform -1 0 1566 0 1 2481
box -28 0 128 267
use sky130_fd_pr__pfet_01v8__example_55959141808628  sky130_fd_pr__pfet_01v8__example_55959141808628_1
timestamp 1624884095
transform 1 0 1310 0 1 2481
box -28 0 128 267
<< labels >>
flabel metal1 s 1806 1938 1826 1958 3 FreeSans 200 0 0 0 SEL_H_N
port 1 nsew
flabel metal1 s 1575 1798 1595 1818 3 FreeSans 200 0 0 0 A_H
port 2 nsew
flabel metal1 s 1731 1831 1751 1851 3 FreeSans 200 0 0 0 Y_H
port 3 nsew
flabel metal1 s 1269 2500 1289 2520 3 FreeSans 200 0 0 0 B_H
port 4 nsew
flabel metal1 s 1346 2321 1372 2354 3 FreeSans 520 0 0 0 SEL_H
port 5 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 12181438
string GDS_START 12172596
<< end >>
