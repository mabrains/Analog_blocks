magic
tech sky130A
magscale 1 2
timestamp 1624884095
<< checkpaint >>
rect -1987 -891 4137 3170
<< nwell >>
rect -439 1874 2086 1910
rect -439 1847 2606 1874
rect 2611 1847 2827 1867
rect -439 1112 2827 1847
rect 434 1052 1568 1112
rect 2606 829 2827 1112
<< pwell >>
rect -727 986 363 1052
rect -727 400 471 986
rect -727 370 -641 400
rect 385 369 471 400
<< mvnmos >>
rect -540 426 -420 1026
rect -364 426 -244 1026
rect -188 426 -68 1026
rect -12 426 108 1026
rect 164 426 284 1026
<< mvpmos >>
rect -189 1208 -89 1808
rect -33 1208 67 1808
rect 123 1208 223 1808
rect 279 1208 379 1808
rect 653 1608 753 1808
rect 809 1608 1009 1808
rect 1065 1608 1265 1808
rect 1687 1608 2487 1808
rect 653 1118 753 1318
rect 809 1118 1009 1318
rect 1065 1118 1265 1318
rect 1687 1314 2487 1514
rect 2677 948 2761 1748
<< mvndiff >>
rect -593 948 -540 1026
rect -593 914 -585 948
rect -551 914 -540 948
rect -593 880 -540 914
rect -593 846 -585 880
rect -551 846 -540 880
rect -593 812 -540 846
rect -593 778 -585 812
rect -551 778 -540 812
rect -593 744 -540 778
rect -593 710 -585 744
rect -551 710 -540 744
rect -593 676 -540 710
rect -593 642 -585 676
rect -551 642 -540 676
rect -593 608 -540 642
rect -593 574 -585 608
rect -551 574 -540 608
rect -593 540 -540 574
rect -593 506 -585 540
rect -551 506 -540 540
rect -593 472 -540 506
rect -593 438 -585 472
rect -551 438 -540 472
rect -593 426 -540 438
rect -420 948 -364 1026
rect -420 914 -409 948
rect -375 914 -364 948
rect -420 880 -364 914
rect -420 846 -409 880
rect -375 846 -364 880
rect -420 812 -364 846
rect -420 778 -409 812
rect -375 778 -364 812
rect -420 744 -364 778
rect -420 710 -409 744
rect -375 710 -364 744
rect -420 676 -364 710
rect -420 642 -409 676
rect -375 642 -364 676
rect -420 608 -364 642
rect -420 574 -409 608
rect -375 574 -364 608
rect -420 540 -364 574
rect -420 506 -409 540
rect -375 506 -364 540
rect -420 472 -364 506
rect -420 438 -409 472
rect -375 438 -364 472
rect -420 426 -364 438
rect -244 948 -188 1026
rect -244 914 -233 948
rect -199 914 -188 948
rect -244 880 -188 914
rect -244 846 -233 880
rect -199 846 -188 880
rect -244 812 -188 846
rect -244 778 -233 812
rect -199 778 -188 812
rect -244 744 -188 778
rect -244 710 -233 744
rect -199 710 -188 744
rect -244 676 -188 710
rect -244 642 -233 676
rect -199 642 -188 676
rect -244 608 -188 642
rect -244 574 -233 608
rect -199 574 -188 608
rect -244 540 -188 574
rect -244 506 -233 540
rect -199 506 -188 540
rect -244 472 -188 506
rect -244 438 -233 472
rect -199 438 -188 472
rect -244 426 -188 438
rect -68 948 -12 1026
rect -68 914 -57 948
rect -23 914 -12 948
rect -68 880 -12 914
rect -68 846 -57 880
rect -23 846 -12 880
rect -68 812 -12 846
rect -68 778 -57 812
rect -23 778 -12 812
rect -68 744 -12 778
rect -68 710 -57 744
rect -23 710 -12 744
rect -68 676 -12 710
rect -68 642 -57 676
rect -23 642 -12 676
rect -68 608 -12 642
rect -68 574 -57 608
rect -23 574 -12 608
rect -68 540 -12 574
rect -68 506 -57 540
rect -23 506 -12 540
rect -68 472 -12 506
rect -68 438 -57 472
rect -23 438 -12 472
rect -68 426 -12 438
rect 108 948 164 1026
rect 108 914 119 948
rect 153 914 164 948
rect 108 880 164 914
rect 108 846 119 880
rect 153 846 164 880
rect 108 812 164 846
rect 108 778 119 812
rect 153 778 164 812
rect 108 744 164 778
rect 108 710 119 744
rect 153 710 164 744
rect 108 676 164 710
rect 108 642 119 676
rect 153 642 164 676
rect 108 608 164 642
rect 108 574 119 608
rect 153 574 164 608
rect 108 540 164 574
rect 108 506 119 540
rect 153 506 164 540
rect 108 472 164 506
rect 108 438 119 472
rect 153 438 164 472
rect 108 426 164 438
rect 284 948 337 1026
rect 284 914 295 948
rect 329 914 337 948
rect 284 880 337 914
rect 284 846 295 880
rect 329 846 337 880
rect 284 812 337 846
rect 284 778 295 812
rect 329 778 337 812
rect 284 744 337 778
rect 284 710 295 744
rect 329 710 337 744
rect 284 676 337 710
rect 284 642 295 676
rect 329 642 337 676
rect 284 608 337 642
rect 284 574 295 608
rect 329 574 337 608
rect 284 540 337 574
rect 284 506 295 540
rect 329 506 337 540
rect 284 472 337 506
rect 284 438 295 472
rect 329 438 337 472
rect 284 426 337 438
<< mvpdiff >>
rect -242 1730 -189 1808
rect -242 1696 -234 1730
rect -200 1696 -189 1730
rect -242 1662 -189 1696
rect -242 1628 -234 1662
rect -200 1628 -189 1662
rect -242 1594 -189 1628
rect -242 1560 -234 1594
rect -200 1560 -189 1594
rect -242 1526 -189 1560
rect -242 1492 -234 1526
rect -200 1492 -189 1526
rect -242 1458 -189 1492
rect -242 1424 -234 1458
rect -200 1424 -189 1458
rect -242 1390 -189 1424
rect -242 1356 -234 1390
rect -200 1356 -189 1390
rect -242 1322 -189 1356
rect -242 1288 -234 1322
rect -200 1288 -189 1322
rect -242 1254 -189 1288
rect -242 1220 -234 1254
rect -200 1220 -189 1254
rect -242 1208 -189 1220
rect -89 1730 -33 1808
rect -89 1696 -78 1730
rect -44 1696 -33 1730
rect -89 1662 -33 1696
rect -89 1628 -78 1662
rect -44 1628 -33 1662
rect -89 1594 -33 1628
rect -89 1560 -78 1594
rect -44 1560 -33 1594
rect -89 1526 -33 1560
rect -89 1492 -78 1526
rect -44 1492 -33 1526
rect -89 1458 -33 1492
rect -89 1424 -78 1458
rect -44 1424 -33 1458
rect -89 1390 -33 1424
rect -89 1356 -78 1390
rect -44 1356 -33 1390
rect -89 1322 -33 1356
rect -89 1288 -78 1322
rect -44 1288 -33 1322
rect -89 1254 -33 1288
rect -89 1220 -78 1254
rect -44 1220 -33 1254
rect -89 1208 -33 1220
rect 67 1730 123 1808
rect 67 1696 78 1730
rect 112 1696 123 1730
rect 67 1662 123 1696
rect 67 1628 78 1662
rect 112 1628 123 1662
rect 67 1594 123 1628
rect 67 1560 78 1594
rect 112 1560 123 1594
rect 67 1526 123 1560
rect 67 1492 78 1526
rect 112 1492 123 1526
rect 67 1458 123 1492
rect 67 1424 78 1458
rect 112 1424 123 1458
rect 67 1390 123 1424
rect 67 1356 78 1390
rect 112 1356 123 1390
rect 67 1322 123 1356
rect 67 1288 78 1322
rect 112 1288 123 1322
rect 67 1254 123 1288
rect 67 1220 78 1254
rect 112 1220 123 1254
rect 67 1208 123 1220
rect 223 1730 279 1808
rect 223 1696 234 1730
rect 268 1696 279 1730
rect 223 1662 279 1696
rect 223 1628 234 1662
rect 268 1628 279 1662
rect 223 1594 279 1628
rect 223 1560 234 1594
rect 268 1560 279 1594
rect 223 1526 279 1560
rect 223 1492 234 1526
rect 268 1492 279 1526
rect 223 1458 279 1492
rect 223 1424 234 1458
rect 268 1424 279 1458
rect 223 1390 279 1424
rect 223 1356 234 1390
rect 268 1356 279 1390
rect 223 1322 279 1356
rect 223 1288 234 1322
rect 268 1288 279 1322
rect 223 1254 279 1288
rect 223 1220 234 1254
rect 268 1220 279 1254
rect 223 1208 279 1220
rect 379 1730 432 1808
rect 379 1696 390 1730
rect 424 1696 432 1730
rect 379 1662 432 1696
rect 379 1628 390 1662
rect 424 1628 432 1662
rect 379 1594 432 1628
rect 600 1796 653 1808
rect 600 1762 608 1796
rect 642 1762 653 1796
rect 600 1728 653 1762
rect 600 1694 608 1728
rect 642 1694 653 1728
rect 600 1660 653 1694
rect 600 1626 608 1660
rect 642 1626 653 1660
rect 600 1608 653 1626
rect 753 1796 809 1808
rect 753 1762 764 1796
rect 798 1762 809 1796
rect 753 1728 809 1762
rect 753 1694 764 1728
rect 798 1694 809 1728
rect 753 1660 809 1694
rect 753 1626 764 1660
rect 798 1626 809 1660
rect 753 1608 809 1626
rect 1009 1796 1065 1808
rect 1009 1762 1020 1796
rect 1054 1762 1065 1796
rect 1009 1728 1065 1762
rect 1009 1694 1020 1728
rect 1054 1694 1065 1728
rect 1009 1660 1065 1694
rect 1009 1626 1020 1660
rect 1054 1626 1065 1660
rect 1009 1608 1065 1626
rect 1265 1796 1318 1808
rect 1265 1762 1276 1796
rect 1310 1762 1318 1796
rect 1265 1728 1318 1762
rect 1265 1694 1276 1728
rect 1310 1694 1318 1728
rect 1265 1660 1318 1694
rect 1265 1626 1276 1660
rect 1310 1626 1318 1660
rect 1265 1608 1318 1626
rect 1634 1796 1687 1808
rect 1634 1762 1642 1796
rect 1676 1762 1687 1796
rect 1634 1728 1687 1762
rect 1634 1694 1642 1728
rect 1676 1694 1687 1728
rect 1634 1660 1687 1694
rect 1634 1626 1642 1660
rect 1676 1626 1687 1660
rect 1634 1608 1687 1626
rect 2487 1796 2540 1808
rect 2487 1762 2498 1796
rect 2532 1762 2540 1796
rect 2487 1728 2540 1762
rect 2677 1793 2761 1801
rect 2677 1759 2715 1793
rect 2749 1759 2761 1793
rect 2677 1748 2761 1759
rect 2487 1694 2498 1728
rect 2532 1694 2540 1728
rect 2487 1660 2540 1694
rect 2487 1626 2498 1660
rect 2532 1626 2540 1660
rect 2487 1608 2540 1626
rect 379 1560 390 1594
rect 424 1560 432 1594
rect 379 1526 432 1560
rect 379 1492 390 1526
rect 424 1492 432 1526
rect 379 1458 432 1492
rect 379 1424 390 1458
rect 424 1424 432 1458
rect 379 1390 432 1424
rect 379 1356 390 1390
rect 424 1356 432 1390
rect 379 1322 432 1356
rect 1634 1496 1687 1514
rect 1634 1462 1642 1496
rect 1676 1462 1687 1496
rect 1634 1428 1687 1462
rect 1634 1394 1642 1428
rect 1676 1394 1687 1428
rect 1634 1360 1687 1394
rect 379 1288 390 1322
rect 424 1288 432 1322
rect 1634 1326 1642 1360
rect 1676 1326 1687 1360
rect 379 1254 432 1288
rect 379 1220 390 1254
rect 424 1220 432 1254
rect 379 1208 432 1220
rect 600 1300 653 1318
rect 600 1266 608 1300
rect 642 1266 653 1300
rect 600 1232 653 1266
rect 600 1198 608 1232
rect 642 1198 653 1232
rect 600 1164 653 1198
rect 600 1130 608 1164
rect 642 1130 653 1164
rect 600 1118 653 1130
rect 753 1300 809 1318
rect 753 1266 764 1300
rect 798 1266 809 1300
rect 753 1232 809 1266
rect 753 1198 764 1232
rect 798 1198 809 1232
rect 753 1164 809 1198
rect 753 1130 764 1164
rect 798 1130 809 1164
rect 753 1118 809 1130
rect 1009 1300 1065 1318
rect 1009 1266 1020 1300
rect 1054 1266 1065 1300
rect 1009 1232 1065 1266
rect 1009 1198 1020 1232
rect 1054 1198 1065 1232
rect 1009 1164 1065 1198
rect 1009 1130 1020 1164
rect 1054 1130 1065 1164
rect 1009 1118 1065 1130
rect 1265 1300 1318 1318
rect 1634 1314 1687 1326
rect 2487 1496 2540 1514
rect 2487 1462 2498 1496
rect 2532 1462 2540 1496
rect 2487 1428 2540 1462
rect 2487 1394 2498 1428
rect 2532 1394 2540 1428
rect 2487 1360 2540 1394
rect 2487 1326 2498 1360
rect 2532 1326 2540 1360
rect 2487 1314 2540 1326
rect 1265 1266 1276 1300
rect 1310 1266 1318 1300
rect 1265 1232 1318 1266
rect 1265 1198 1276 1232
rect 1310 1198 1318 1232
rect 1265 1164 1318 1198
rect 1265 1130 1276 1164
rect 1310 1130 1318 1164
rect 1265 1118 1318 1130
rect 2677 937 2761 948
rect 2677 903 2715 937
rect 2749 903 2761 937
rect 2677 895 2761 903
<< mvndiffc >>
rect -585 914 -551 948
rect -585 846 -551 880
rect -585 778 -551 812
rect -585 710 -551 744
rect -585 642 -551 676
rect -585 574 -551 608
rect -585 506 -551 540
rect -585 438 -551 472
rect -409 914 -375 948
rect -409 846 -375 880
rect -409 778 -375 812
rect -409 710 -375 744
rect -409 642 -375 676
rect -409 574 -375 608
rect -409 506 -375 540
rect -409 438 -375 472
rect -233 914 -199 948
rect -233 846 -199 880
rect -233 778 -199 812
rect -233 710 -199 744
rect -233 642 -199 676
rect -233 574 -199 608
rect -233 506 -199 540
rect -233 438 -199 472
rect -57 914 -23 948
rect -57 846 -23 880
rect -57 778 -23 812
rect -57 710 -23 744
rect -57 642 -23 676
rect -57 574 -23 608
rect -57 506 -23 540
rect -57 438 -23 472
rect 119 914 153 948
rect 119 846 153 880
rect 119 778 153 812
rect 119 710 153 744
rect 119 642 153 676
rect 119 574 153 608
rect 119 506 153 540
rect 119 438 153 472
rect 295 914 329 948
rect 295 846 329 880
rect 295 778 329 812
rect 295 710 329 744
rect 295 642 329 676
rect 295 574 329 608
rect 295 506 329 540
rect 295 438 329 472
<< mvpdiffc >>
rect -234 1696 -200 1730
rect -234 1628 -200 1662
rect -234 1560 -200 1594
rect -234 1492 -200 1526
rect -234 1424 -200 1458
rect -234 1356 -200 1390
rect -234 1288 -200 1322
rect -234 1220 -200 1254
rect -78 1696 -44 1730
rect -78 1628 -44 1662
rect -78 1560 -44 1594
rect -78 1492 -44 1526
rect -78 1424 -44 1458
rect -78 1356 -44 1390
rect -78 1288 -44 1322
rect -78 1220 -44 1254
rect 78 1696 112 1730
rect 78 1628 112 1662
rect 78 1560 112 1594
rect 78 1492 112 1526
rect 78 1424 112 1458
rect 78 1356 112 1390
rect 78 1288 112 1322
rect 78 1220 112 1254
rect 234 1696 268 1730
rect 234 1628 268 1662
rect 234 1560 268 1594
rect 234 1492 268 1526
rect 234 1424 268 1458
rect 234 1356 268 1390
rect 234 1288 268 1322
rect 234 1220 268 1254
rect 390 1696 424 1730
rect 390 1628 424 1662
rect 608 1762 642 1796
rect 608 1694 642 1728
rect 608 1626 642 1660
rect 764 1762 798 1796
rect 764 1694 798 1728
rect 764 1626 798 1660
rect 1020 1762 1054 1796
rect 1020 1694 1054 1728
rect 1020 1626 1054 1660
rect 1276 1762 1310 1796
rect 1276 1694 1310 1728
rect 1276 1626 1310 1660
rect 1642 1762 1676 1796
rect 1642 1694 1676 1728
rect 1642 1626 1676 1660
rect 2498 1762 2532 1796
rect 2715 1759 2749 1793
rect 2498 1694 2532 1728
rect 2498 1626 2532 1660
rect 390 1560 424 1594
rect 390 1492 424 1526
rect 390 1424 424 1458
rect 390 1356 424 1390
rect 1642 1462 1676 1496
rect 1642 1394 1676 1428
rect 390 1288 424 1322
rect 1642 1326 1676 1360
rect 390 1220 424 1254
rect 608 1266 642 1300
rect 608 1198 642 1232
rect 608 1130 642 1164
rect 764 1266 798 1300
rect 764 1198 798 1232
rect 764 1130 798 1164
rect 1020 1266 1054 1300
rect 1020 1198 1054 1232
rect 1020 1130 1054 1164
rect 2498 1462 2532 1496
rect 2498 1394 2532 1428
rect 2498 1326 2532 1360
rect 1276 1266 1310 1300
rect 1276 1198 1310 1232
rect 1276 1130 1310 1164
rect 2715 903 2749 937
<< mvpsubdiff >>
rect -701 992 -667 1026
rect -701 924 -667 958
rect -701 856 -667 890
rect -701 788 -667 822
rect -701 720 -667 754
rect -701 652 -667 686
rect -701 584 -667 618
rect -701 516 -667 550
rect -701 396 -667 482
rect 411 936 445 960
rect 411 867 445 902
rect 411 798 445 833
rect 411 729 445 764
rect 411 660 445 695
rect 411 591 445 626
rect 411 522 445 557
rect 411 453 445 488
rect 411 395 445 419
<< mvnsubdiff >>
rect -350 1814 -316 1838
rect -350 1745 -316 1780
rect -350 1676 -316 1711
rect -350 1607 -316 1642
rect -350 1538 -316 1573
rect -350 1470 -316 1504
rect -350 1402 -316 1436
rect -350 1334 -316 1368
rect -350 1266 -316 1300
rect -350 1208 -316 1232
<< mvpsubdiffcont >>
rect -701 958 -667 992
rect -701 890 -667 924
rect -701 822 -667 856
rect -701 754 -667 788
rect -701 686 -667 720
rect -701 618 -667 652
rect -701 550 -667 584
rect -701 482 -667 516
rect 411 902 445 936
rect 411 833 445 867
rect 411 764 445 798
rect 411 695 445 729
rect 411 626 445 660
rect 411 557 445 591
rect 411 488 445 522
rect 411 419 445 453
<< mvnsubdiffcont >>
rect -350 1780 -316 1814
rect -350 1711 -316 1745
rect -350 1642 -316 1676
rect -350 1573 -316 1607
rect -350 1504 -316 1538
rect -350 1436 -316 1470
rect -350 1368 -316 1402
rect -350 1300 -316 1334
rect -350 1232 -316 1266
<< poly >>
rect -189 1890 379 1906
rect -189 1856 -158 1890
rect -124 1856 -90 1890
rect -56 1856 -22 1890
rect 12 1856 46 1890
rect 80 1856 114 1890
rect 148 1856 182 1890
rect 216 1856 250 1890
rect 284 1856 318 1890
rect 352 1856 379 1890
rect -189 1834 379 1856
rect -189 1808 -89 1834
rect -33 1808 67 1834
rect 123 1808 223 1834
rect 279 1808 379 1834
rect 653 1890 1265 1906
rect 653 1856 675 1890
rect 709 1856 753 1890
rect 787 1856 830 1890
rect 864 1856 907 1890
rect 941 1856 984 1890
rect 1018 1856 1061 1890
rect 1095 1856 1138 1890
rect 1172 1856 1215 1890
rect 1249 1856 1265 1890
rect 653 1840 1265 1856
rect 653 1834 1009 1840
rect 653 1808 753 1834
rect 809 1808 1009 1834
rect 1065 1808 1265 1840
rect 1687 1890 2487 1906
rect 1687 1856 1718 1890
rect 1752 1856 1786 1890
rect 1820 1856 1854 1890
rect 1888 1856 1922 1890
rect 1956 1856 1990 1890
rect 2024 1856 2058 1890
rect 2092 1856 2126 1890
rect 2160 1856 2194 1890
rect 2228 1856 2262 1890
rect 2296 1856 2330 1890
rect 2364 1856 2398 1890
rect 2432 1856 2487 1890
rect 1687 1808 2487 1856
rect 2579 1707 2677 1748
rect 2579 1673 2595 1707
rect 2629 1673 2677 1707
rect 2579 1637 2677 1673
rect 653 1582 753 1608
rect 809 1582 1009 1608
rect 1065 1582 1265 1608
rect 1687 1582 2487 1608
rect 2579 1603 2595 1637
rect 2629 1603 2677 1637
rect 2579 1566 2677 1603
rect 1687 1514 2487 1540
rect 2579 1532 2595 1566
rect 2629 1532 2677 1566
rect 653 1318 753 1344
rect 809 1318 1009 1344
rect 1065 1318 1265 1344
rect -189 1182 -89 1208
rect -33 1182 67 1208
rect 123 1182 223 1208
rect 279 1182 379 1208
rect -540 1108 284 1124
rect 2579 1495 2677 1532
rect 2579 1461 2595 1495
rect 2629 1461 2677 1495
rect 2579 1424 2677 1461
rect 2579 1390 2595 1424
rect 2629 1390 2677 1424
rect 2579 1353 2677 1390
rect 2579 1319 2595 1353
rect 2629 1319 2677 1353
rect 1687 1266 2487 1314
rect 1687 1232 1735 1266
rect 1769 1232 1803 1266
rect 1837 1232 1871 1266
rect 1905 1232 1939 1266
rect 1973 1232 2007 1266
rect 2041 1232 2075 1266
rect 2109 1232 2143 1266
rect 2177 1232 2211 1266
rect 2245 1232 2279 1266
rect 2313 1232 2347 1266
rect 2381 1232 2415 1266
rect 2449 1232 2487 1266
rect 1687 1216 2487 1232
rect 2579 1282 2677 1319
rect 2579 1248 2595 1282
rect 2629 1248 2677 1282
rect 2579 1211 2677 1248
rect 2579 1177 2595 1211
rect 2629 1177 2677 1211
rect 2579 1140 2677 1177
rect -540 1074 -524 1108
rect -490 1074 -455 1108
rect -421 1074 -386 1108
rect -352 1074 -317 1108
rect -283 1074 -248 1108
rect -214 1074 -179 1108
rect -145 1074 -110 1108
rect -76 1074 -41 1108
rect -7 1074 28 1108
rect 62 1074 97 1108
rect 131 1074 166 1108
rect 200 1074 234 1108
rect 268 1074 284 1108
rect -540 1052 284 1074
rect -540 1026 -420 1052
rect -364 1026 -244 1052
rect -188 1026 -68 1052
rect -12 1026 108 1052
rect 164 1026 284 1052
rect 653 1092 753 1118
rect 809 1092 1009 1118
rect 1065 1092 1265 1118
rect 653 1013 1265 1092
rect 653 979 669 1013
rect 703 979 738 1013
rect 772 979 807 1013
rect 841 979 875 1013
rect 909 979 943 1013
rect 977 979 1011 1013
rect 1045 979 1079 1013
rect 1113 979 1147 1013
rect 1181 979 1215 1013
rect 1249 979 1265 1013
rect 653 963 1265 979
rect 2579 1106 2595 1140
rect 2629 1106 2677 1140
rect 2579 1069 2677 1106
rect 2579 1035 2595 1069
rect 2629 1035 2677 1069
rect 2579 998 2677 1035
rect 2579 964 2595 998
rect 2629 964 2677 998
rect 2579 948 2677 964
rect 2761 948 2793 1748
rect -540 400 -420 426
rect -364 400 -244 426
rect -188 400 -68 426
rect -12 400 108 426
rect 164 400 284 426
<< polycont >>
rect -158 1856 -124 1890
rect -90 1856 -56 1890
rect -22 1856 12 1890
rect 46 1856 80 1890
rect 114 1856 148 1890
rect 182 1856 216 1890
rect 250 1856 284 1890
rect 318 1856 352 1890
rect 675 1856 709 1890
rect 753 1856 787 1890
rect 830 1856 864 1890
rect 907 1856 941 1890
rect 984 1856 1018 1890
rect 1061 1856 1095 1890
rect 1138 1856 1172 1890
rect 1215 1856 1249 1890
rect 1718 1856 1752 1890
rect 1786 1856 1820 1890
rect 1854 1856 1888 1890
rect 1922 1856 1956 1890
rect 1990 1856 2024 1890
rect 2058 1856 2092 1890
rect 2126 1856 2160 1890
rect 2194 1856 2228 1890
rect 2262 1856 2296 1890
rect 2330 1856 2364 1890
rect 2398 1856 2432 1890
rect 2595 1673 2629 1707
rect 2595 1603 2629 1637
rect 2595 1532 2629 1566
rect 2595 1461 2629 1495
rect 2595 1390 2629 1424
rect 2595 1319 2629 1353
rect 1735 1232 1769 1266
rect 1803 1232 1837 1266
rect 1871 1232 1905 1266
rect 1939 1232 1973 1266
rect 2007 1232 2041 1266
rect 2075 1232 2109 1266
rect 2143 1232 2177 1266
rect 2211 1232 2245 1266
rect 2279 1232 2313 1266
rect 2347 1232 2381 1266
rect 2415 1232 2449 1266
rect 2595 1248 2629 1282
rect 2595 1177 2629 1211
rect -524 1074 -490 1108
rect -455 1074 -421 1108
rect -386 1074 -352 1108
rect -317 1074 -283 1108
rect -248 1074 -214 1108
rect -179 1074 -145 1108
rect -110 1074 -76 1108
rect -41 1074 -7 1108
rect 28 1074 62 1108
rect 97 1074 131 1108
rect 166 1074 200 1108
rect 234 1074 268 1108
rect 669 979 703 1013
rect 738 979 772 1013
rect 807 979 841 1013
rect 875 979 909 1013
rect 943 979 977 1013
rect 1011 979 1045 1013
rect 1079 979 1113 1013
rect 1147 979 1181 1013
rect 1215 979 1249 1013
rect 2595 1106 2629 1140
rect 2595 1035 2629 1069
rect 2595 964 2629 998
<< locali >>
rect -175 1859 -158 1890
rect -124 1859 -90 1890
rect -56 1859 -22 1890
rect 12 1859 46 1890
rect -350 1814 -316 1838
rect -175 1825 -174 1859
rect -124 1856 -102 1859
rect -56 1856 -30 1859
rect 12 1856 42 1859
rect 80 1856 114 1890
rect 148 1856 182 1890
rect 216 1859 250 1890
rect 284 1859 318 1890
rect 352 1859 368 1890
rect 220 1856 250 1859
rect 292 1856 318 1859
rect -140 1825 -102 1856
rect -68 1825 -30 1856
rect 4 1825 42 1856
rect 76 1825 114 1856
rect 148 1825 186 1856
rect 220 1825 258 1856
rect 292 1825 330 1856
rect 364 1825 368 1859
rect 659 1856 675 1890
rect 709 1856 753 1890
rect 787 1856 830 1890
rect 864 1856 907 1890
rect 941 1856 984 1890
rect 1018 1856 1061 1890
rect 1095 1856 1138 1890
rect 1172 1856 1215 1890
rect 1249 1856 1265 1890
rect 1702 1859 1718 1890
rect 1752 1859 1786 1890
rect 1702 1856 1710 1859
rect 1752 1856 1782 1859
rect 1820 1856 1854 1890
rect 1888 1856 1922 1890
rect 1956 1859 1990 1890
rect 2024 1859 2058 1890
rect 2092 1859 2126 1890
rect 2160 1859 2194 1890
rect 2228 1859 2262 1890
rect 2296 1859 2330 1890
rect 2364 1859 2398 1890
rect 2432 1859 2456 1890
rect 1960 1856 1990 1859
rect 2032 1856 2058 1859
rect 2104 1856 2126 1859
rect 2176 1856 2194 1859
rect 2248 1856 2262 1859
rect 2320 1856 2330 1859
rect 2392 1856 2398 1859
rect 1744 1825 1782 1856
rect 1816 1825 1854 1856
rect 1888 1825 1926 1856
rect 1960 1825 1998 1856
rect 2032 1825 2070 1856
rect 2104 1825 2142 1856
rect 2176 1825 2214 1856
rect 2248 1825 2286 1856
rect 2320 1825 2358 1856
rect 2392 1825 2430 1856
rect -350 1745 -316 1780
rect 547 1796 653 1812
rect 547 1762 608 1796
rect 642 1762 653 1796
rect -350 1676 -316 1711
rect -350 1607 -316 1642
rect -350 1538 -316 1573
rect -350 1470 -316 1504
rect -350 1402 -316 1436
rect -350 1334 -316 1368
rect -350 1266 -316 1300
rect -350 1181 -316 1219
rect -234 1730 -200 1746
rect -234 1662 -200 1696
rect -234 1594 -200 1628
rect -234 1555 -200 1560
rect -78 1730 -44 1746
rect -78 1662 -44 1696
rect -78 1594 -44 1628
rect -200 1521 -162 1555
rect -78 1526 -44 1560
rect 78 1730 112 1746
rect 78 1662 112 1696
rect 78 1594 112 1628
rect 78 1555 112 1560
rect 234 1730 268 1746
rect 234 1662 268 1696
rect 234 1594 268 1628
rect -234 1458 -200 1492
rect -234 1390 -200 1424
rect 77 1526 115 1555
rect 77 1521 78 1526
rect -78 1458 -44 1492
rect -78 1401 -44 1424
rect 112 1521 115 1526
rect 234 1526 268 1560
rect 390 1730 424 1746
rect 390 1662 424 1696
rect 390 1594 424 1628
rect 390 1555 424 1560
rect 547 1728 653 1762
rect 547 1694 608 1728
rect 642 1694 653 1728
rect 547 1660 653 1694
rect 547 1626 608 1660
rect 642 1626 653 1660
rect 78 1458 112 1492
rect 354 1526 392 1555
rect 354 1521 390 1526
rect 234 1475 268 1492
rect 234 1458 272 1475
rect -62 1390 -24 1401
rect -44 1367 -24 1390
rect 78 1390 112 1424
rect -234 1322 -200 1356
rect -234 1254 -200 1288
rect -234 1204 -200 1220
rect -78 1322 -44 1356
rect -78 1254 -44 1288
rect -78 1204 -44 1220
rect 78 1322 112 1356
rect 78 1254 112 1288
rect 78 1204 112 1220
rect 268 1441 272 1458
rect 390 1458 424 1492
rect 234 1390 268 1424
rect 234 1322 268 1356
rect 234 1254 268 1288
rect 234 1204 268 1220
rect 390 1390 424 1424
rect 390 1322 424 1356
rect 390 1254 424 1288
rect 390 1204 424 1220
rect 547 1475 653 1626
rect 581 1441 619 1475
rect 547 1300 653 1441
rect 547 1266 608 1300
rect 642 1266 653 1300
rect 547 1232 653 1266
rect 547 1198 608 1232
rect 642 1198 653 1232
rect 547 1164 653 1198
rect 547 1130 608 1164
rect 642 1130 653 1164
rect 547 1114 653 1130
rect 700 1796 830 1812
rect 700 1762 764 1796
rect 798 1762 830 1796
rect 700 1728 830 1762
rect 700 1694 764 1728
rect 798 1694 830 1728
rect 700 1660 830 1694
rect 700 1626 764 1660
rect 798 1626 830 1660
rect 700 1300 830 1626
rect 700 1266 764 1300
rect 798 1266 830 1300
rect 700 1259 830 1266
rect 700 1225 712 1259
rect 746 1232 784 1259
rect 746 1225 764 1232
rect 818 1225 830 1259
rect 700 1198 764 1225
rect 798 1198 830 1225
rect 700 1181 830 1198
rect 700 1147 712 1181
rect 746 1164 784 1181
rect 746 1147 764 1164
rect 818 1147 830 1181
rect 700 1130 764 1147
rect 798 1130 830 1147
rect -540 1074 -524 1108
rect -490 1074 -455 1108
rect -421 1074 -386 1108
rect -352 1074 -317 1108
rect -283 1074 -248 1108
rect -214 1074 -179 1108
rect -145 1074 -110 1108
rect -76 1074 -41 1108
rect -7 1074 28 1108
rect 62 1074 97 1108
rect 131 1074 166 1108
rect 200 1074 234 1108
rect 268 1074 284 1108
rect 700 1103 830 1130
rect 999 1796 1105 1812
rect 999 1762 1020 1796
rect 1054 1762 1105 1796
rect 999 1728 1105 1762
rect 999 1694 1020 1728
rect 1054 1694 1105 1728
rect 999 1660 1105 1694
rect 999 1626 1020 1660
rect 1054 1626 1105 1660
rect 999 1401 1105 1626
rect 1033 1367 1071 1401
rect 999 1300 1105 1367
rect 999 1266 1020 1300
rect 1054 1266 1105 1300
rect 999 1232 1105 1266
rect 999 1198 1020 1232
rect 1054 1198 1105 1232
rect 999 1164 1105 1198
rect 999 1130 1020 1164
rect 1054 1130 1105 1164
rect 999 1114 1105 1130
rect 1152 1796 1347 1812
rect 1152 1762 1276 1796
rect 1310 1762 1347 1796
rect 1152 1728 1347 1762
rect 1152 1694 1276 1728
rect 1310 1694 1347 1728
rect 1152 1660 1347 1694
rect 1152 1626 1276 1660
rect 1310 1626 1347 1660
rect 1152 1300 1347 1626
rect 1152 1266 1276 1300
rect 1310 1266 1347 1300
rect 1152 1259 1347 1266
rect 1152 1225 1164 1259
rect 1198 1232 1301 1259
rect 1198 1225 1276 1232
rect 1335 1225 1347 1259
rect 1152 1198 1276 1225
rect 1310 1198 1347 1225
rect 1152 1181 1347 1198
rect 1152 1147 1164 1181
rect 1198 1164 1301 1181
rect 1198 1147 1276 1164
rect 1335 1147 1347 1181
rect 1152 1130 1276 1147
rect 1310 1130 1347 1147
rect -701 992 -667 1026
rect -321 1023 -268 1074
rect -321 989 -311 1023
rect -277 989 -268 1023
rect -701 924 -667 958
rect -701 856 -667 890
rect -701 788 -667 822
rect -701 720 -667 754
rect -701 656 -667 686
rect -671 652 -667 656
rect -705 618 -701 622
rect -705 584 -667 618
rect -701 516 -667 550
rect -701 396 -667 482
rect -585 948 -479 964
rect -551 914 -479 948
rect -585 880 -479 914
rect -551 871 -479 880
rect -551 837 -513 871
rect -585 812 -479 837
rect -551 778 -479 812
rect -585 744 -479 778
rect -551 710 -479 744
rect -585 676 -479 710
rect -551 642 -479 676
rect -585 608 -479 642
rect -551 574 -479 608
rect -585 540 -479 574
rect -551 506 -479 540
rect -585 472 -479 506
rect -551 438 -479 472
rect -585 422 -479 438
rect -429 948 -355 964
rect -429 914 -409 948
rect -375 914 -355 948
rect -429 880 -355 914
rect -321 951 -268 989
rect -162 1023 -91 1074
rect -162 989 -143 1023
rect -109 989 -91 1023
rect -321 917 -311 951
rect -277 917 -268 951
rect -321 905 -268 917
rect -233 948 -199 964
rect -429 846 -409 880
rect -375 846 -355 880
rect -233 880 -199 914
rect -162 951 -91 989
rect 11 1023 85 1074
rect 11 989 33 1023
rect 67 989 85 1023
rect -162 917 -143 951
rect -109 917 -91 951
rect -162 905 -91 917
rect -57 948 -23 964
rect -57 880 -23 914
rect 11 951 85 989
rect 187 1023 240 1074
rect 700 1069 712 1103
rect 746 1069 784 1103
rect 818 1069 830 1103
rect 700 1063 830 1069
rect 1152 1103 1347 1130
rect 1152 1069 1164 1103
rect 1198 1069 1301 1103
rect 1335 1069 1347 1103
rect 1152 1063 1347 1069
rect 1410 1259 1586 1812
rect 1642 1796 1676 1812
rect 2498 1796 2765 1874
rect 1676 1762 1828 1791
rect 1642 1728 1828 1762
rect 1676 1694 1828 1728
rect 1642 1660 1828 1694
rect 1676 1626 1828 1660
rect 1642 1555 1828 1626
rect 1756 1521 1794 1555
rect 2532 1793 2765 1796
rect 2532 1762 2715 1793
rect 2498 1759 2715 1762
rect 2749 1759 2765 1793
rect 2498 1728 2532 1759
rect 2498 1660 2532 1694
rect 1410 1225 1422 1259
rect 1456 1225 1540 1259
rect 1574 1225 1586 1259
rect 1410 1181 1586 1225
rect 1410 1147 1422 1181
rect 1456 1147 1540 1181
rect 1574 1147 1586 1181
rect 1642 1496 1676 1512
rect 1642 1428 1676 1462
rect 1642 1360 1676 1394
rect 2498 1496 2532 1626
rect 2498 1428 2532 1462
rect 2498 1360 2532 1394
rect 1642 1253 1676 1326
rect 1642 1181 1676 1219
rect 1719 1333 2464 1339
rect 1719 1299 1743 1333
rect 1777 1299 1815 1333
rect 1849 1299 1887 1333
rect 1921 1299 1959 1333
rect 1993 1299 2031 1333
rect 2065 1299 2103 1333
rect 2137 1299 2175 1333
rect 2209 1299 2247 1333
rect 2281 1299 2319 1333
rect 2353 1299 2391 1333
rect 2425 1299 2464 1333
rect 2498 1310 2532 1326
rect 2595 1707 2629 1723
rect 2595 1637 2629 1673
rect 2595 1566 2629 1603
rect 2595 1495 2629 1532
rect 2595 1424 2629 1461
rect 2595 1353 2629 1390
rect 1719 1275 2464 1299
rect 2595 1282 2629 1319
rect 1719 1266 2595 1275
rect 1719 1232 1735 1266
rect 1769 1232 1803 1266
rect 1837 1232 1871 1266
rect 1905 1232 1939 1266
rect 1973 1232 2007 1266
rect 2041 1232 2075 1266
rect 2109 1232 2143 1266
rect 2177 1232 2211 1266
rect 2245 1232 2279 1266
rect 2313 1232 2347 1266
rect 2381 1232 2415 1266
rect 2449 1248 2595 1266
rect 2449 1232 2629 1248
rect 1719 1211 2629 1232
rect 1719 1187 2595 1211
rect 1410 1103 1586 1147
rect 1410 1069 1422 1103
rect 1456 1069 1540 1103
rect 1574 1069 1586 1103
rect 187 989 201 1023
rect 235 989 240 1023
rect 11 917 33 951
rect 67 917 85 951
rect 11 905 85 917
rect 119 948 153 964
rect -429 812 -355 846
rect -199 846 -191 871
rect -229 837 -191 846
rect -77 846 -57 871
rect 119 880 153 914
rect 187 951 240 989
rect 187 917 201 951
rect 235 917 240 951
rect 187 905 240 917
rect 275 948 450 1035
rect 653 979 669 1013
rect 703 979 738 1013
rect 772 979 807 1013
rect 841 979 875 1013
rect 909 979 943 1013
rect 977 979 1011 1013
rect 1045 979 1079 1013
rect 1113 979 1147 1013
rect 1181 979 1215 1013
rect 1249 979 1265 1013
rect 275 914 295 948
rect 329 936 450 948
rect 329 914 411 936
rect 275 902 411 914
rect 445 902 450 936
rect 275 880 450 902
rect -23 846 -3 871
rect -429 778 -409 812
rect -375 778 -355 812
rect -429 744 -355 778
rect -429 710 -409 744
rect -375 710 -355 744
rect -429 676 -355 710
rect -429 622 -409 676
rect -375 622 -355 676
rect -429 608 -355 622
rect -429 550 -409 608
rect -375 550 -355 608
rect -429 540 -355 550
rect -429 506 -409 540
rect -375 506 -355 540
rect -429 472 -355 506
rect -429 438 -409 472
rect -375 438 -355 472
rect -429 422 -355 438
rect -233 812 -199 837
rect -233 744 -199 778
rect -233 676 -199 710
rect -233 608 -199 642
rect -233 540 -199 574
rect -233 472 -199 506
rect -233 422 -199 438
rect -77 812 -3 846
rect -77 778 -57 812
rect -23 778 -3 812
rect -77 744 -3 778
rect -77 710 -57 744
rect -23 710 -3 744
rect -77 676 -3 710
rect -77 622 -57 676
rect -23 622 -3 676
rect -77 608 -3 622
rect -77 550 -57 608
rect -23 550 -3 608
rect -77 540 -3 550
rect -77 506 -57 540
rect -23 506 -3 540
rect -77 472 -3 506
rect -77 438 -57 472
rect -23 438 -3 472
rect -77 422 -3 438
rect 81 837 119 871
rect 153 837 173 871
rect 47 812 173 837
rect 47 778 119 812
rect 153 778 173 812
rect 47 744 173 778
rect 47 710 119 744
rect 153 710 173 744
rect 47 676 173 710
rect 47 642 119 676
rect 153 642 173 676
rect 47 608 173 642
rect 47 574 119 608
rect 153 574 173 608
rect 47 540 173 574
rect 47 506 119 540
rect 153 506 173 540
rect 47 472 173 506
rect 47 438 119 472
rect 153 438 173 472
rect 47 422 173 438
rect 275 846 295 880
rect 329 867 450 880
rect 329 846 411 867
rect 275 833 411 846
rect 445 833 450 867
rect 275 812 450 833
rect 275 778 295 812
rect 329 798 450 812
rect 329 778 411 798
rect 275 764 411 778
rect 445 764 450 798
rect 275 744 450 764
rect 275 710 295 744
rect 329 729 450 744
rect 329 710 411 729
rect 275 695 411 710
rect 445 695 450 729
rect 275 676 450 695
rect 275 656 295 676
rect 329 660 450 676
rect 275 622 294 656
rect 329 642 411 660
rect 328 622 411 642
rect 445 622 450 660
rect 275 608 450 622
rect 275 584 295 608
rect 329 591 450 608
rect 275 550 294 584
rect 329 574 411 591
rect 328 550 411 574
rect 445 550 450 591
rect 275 540 450 550
rect 1410 542 1586 1069
rect 2595 1140 2629 1177
rect 2595 1069 2629 1106
rect 2595 998 2629 1035
rect 2595 948 2629 964
rect 2663 1251 2827 1265
rect 2663 1217 2667 1251
rect 2701 1217 2793 1251
rect 2663 1110 2827 1217
rect 2663 1076 2667 1110
rect 2701 1076 2793 1110
rect 2663 937 2827 1076
rect 2663 903 2715 937
rect 2749 903 2827 937
rect 2663 898 2827 903
rect 275 506 295 540
rect 329 522 450 540
rect 329 506 411 522
rect 275 488 411 506
rect 445 488 450 522
rect 275 472 450 488
rect 275 438 295 472
rect 329 453 450 472
rect 329 438 411 453
rect 275 419 411 438
rect 445 419 450 453
rect 275 396 450 419
rect 411 395 445 396
<< viali >>
rect -174 1856 -158 1859
rect -158 1856 -140 1859
rect -102 1856 -90 1859
rect -90 1856 -68 1859
rect -30 1856 -22 1859
rect -22 1856 4 1859
rect 42 1856 46 1859
rect 46 1856 76 1859
rect 114 1856 148 1859
rect 186 1856 216 1859
rect 216 1856 220 1859
rect 258 1856 284 1859
rect 284 1856 292 1859
rect 330 1856 352 1859
rect 352 1856 364 1859
rect -174 1825 -140 1856
rect -102 1825 -68 1856
rect -30 1825 4 1856
rect 42 1825 76 1856
rect 114 1825 148 1856
rect 186 1825 220 1856
rect 258 1825 292 1856
rect 330 1825 364 1856
rect 1710 1856 1718 1859
rect 1718 1856 1744 1859
rect 1782 1856 1786 1859
rect 1786 1856 1816 1859
rect 1854 1856 1888 1859
rect 1926 1856 1956 1859
rect 1956 1856 1960 1859
rect 1998 1856 2024 1859
rect 2024 1856 2032 1859
rect 2070 1856 2092 1859
rect 2092 1856 2104 1859
rect 2142 1856 2160 1859
rect 2160 1856 2176 1859
rect 2214 1856 2228 1859
rect 2228 1856 2248 1859
rect 2286 1856 2296 1859
rect 2296 1856 2320 1859
rect 2358 1856 2364 1859
rect 2364 1856 2392 1859
rect 2430 1856 2432 1859
rect 2432 1856 2464 1859
rect 1710 1825 1744 1856
rect 1782 1825 1816 1856
rect 1854 1825 1888 1856
rect 1926 1825 1960 1856
rect 1998 1825 2032 1856
rect 2070 1825 2104 1856
rect 2142 1825 2176 1856
rect 2214 1825 2248 1856
rect 2286 1825 2320 1856
rect 2358 1825 2392 1856
rect 2430 1825 2464 1856
rect -350 1232 -316 1253
rect -350 1219 -316 1232
rect -234 1526 -200 1555
rect -234 1521 -200 1526
rect -162 1521 -128 1555
rect 43 1521 77 1555
rect 115 1521 149 1555
rect 320 1521 354 1555
rect 392 1526 426 1555
rect 392 1521 424 1526
rect 424 1521 426 1526
rect 200 1441 234 1475
rect -96 1390 -62 1401
rect -96 1367 -78 1390
rect -78 1367 -62 1390
rect -24 1367 10 1401
rect 272 1441 306 1475
rect 547 1441 581 1475
rect 619 1441 653 1475
rect -350 1147 -316 1181
rect 712 1225 746 1259
rect 784 1232 818 1259
rect 784 1225 798 1232
rect 798 1225 818 1232
rect 712 1147 746 1181
rect 784 1164 818 1181
rect 784 1147 798 1164
rect 798 1147 818 1164
rect 999 1367 1033 1401
rect 1071 1367 1105 1401
rect 1164 1225 1198 1259
rect 1301 1232 1335 1259
rect 1301 1225 1310 1232
rect 1310 1225 1335 1232
rect 1164 1147 1198 1181
rect 1301 1164 1335 1181
rect 1301 1147 1310 1164
rect 1310 1147 1335 1164
rect -311 989 -277 1023
rect -705 652 -671 656
rect -705 622 -701 652
rect -701 622 -671 652
rect -705 550 -701 584
rect -701 550 -671 584
rect -585 846 -551 871
rect -585 837 -551 846
rect -513 837 -479 871
rect -143 989 -109 1023
rect -311 917 -277 951
rect 33 989 67 1023
rect -143 917 -109 951
rect 712 1069 746 1103
rect 784 1069 818 1103
rect 1164 1069 1198 1103
rect 1301 1069 1335 1103
rect 1722 1521 1756 1555
rect 1794 1521 1828 1555
rect 1422 1225 1456 1259
rect 1540 1225 1574 1259
rect 1422 1147 1456 1181
rect 1540 1147 1574 1181
rect 1642 1219 1676 1253
rect 1743 1299 1777 1333
rect 1815 1299 1849 1333
rect 1887 1299 1921 1333
rect 1959 1299 1993 1333
rect 2031 1299 2065 1333
rect 2103 1299 2137 1333
rect 2175 1299 2209 1333
rect 2247 1299 2281 1333
rect 2319 1299 2353 1333
rect 2391 1299 2425 1333
rect 1642 1147 1676 1181
rect 1422 1069 1456 1103
rect 1540 1069 1574 1103
rect 201 989 235 1023
rect 33 917 67 951
rect -263 846 -233 871
rect -233 846 -229 871
rect -263 837 -229 846
rect -191 837 -157 871
rect 201 917 235 951
rect -409 642 -375 656
rect -409 622 -375 642
rect -409 574 -375 584
rect -409 550 -375 574
rect -57 642 -23 656
rect -57 622 -23 642
rect -57 574 -23 584
rect -57 550 -23 574
rect 47 837 81 871
rect 119 846 153 871
rect 119 837 153 846
rect 294 642 295 656
rect 295 642 328 656
rect 294 622 328 642
rect 411 626 445 656
rect 411 622 445 626
rect 294 574 295 584
rect 295 574 328 584
rect 294 550 328 574
rect 411 557 445 584
rect 411 550 445 557
rect 2667 1217 2701 1251
rect 2793 1217 2827 1251
rect 2667 1076 2701 1110
rect 2793 1076 2827 1110
<< metal1 >>
rect -528 1819 -522 1871
rect -470 1819 -458 1871
rect -406 1859 2476 1871
rect -406 1825 -174 1859
rect -140 1825 -102 1859
rect -68 1825 -30 1859
rect 4 1825 42 1859
rect 76 1825 114 1859
rect 148 1825 186 1859
rect 220 1825 258 1859
rect 292 1825 330 1859
rect 364 1825 1710 1859
rect 1744 1825 1782 1859
rect 1816 1825 1854 1859
rect 1888 1825 1926 1859
rect 1960 1825 1998 1859
rect 2032 1825 2070 1859
rect 2104 1825 2142 1859
rect 2176 1825 2214 1859
rect 2248 1825 2286 1859
rect 2320 1825 2358 1859
rect 2392 1825 2430 1859
rect 2464 1825 2476 1859
rect -406 1819 2476 1825
rect -520 1589 2606 1791
rect -246 1555 1718 1561
rect -246 1521 -234 1555
rect -200 1521 -162 1555
rect -128 1521 43 1555
rect 77 1521 115 1555
rect 149 1521 320 1555
rect 354 1521 392 1555
rect 426 1521 1718 1555
rect -246 1509 1718 1521
rect 1770 1509 1782 1561
rect 1834 1509 1840 1561
rect -124 1475 1359 1481
rect -124 1441 200 1475
rect 234 1441 272 1475
rect 306 1441 547 1475
rect 581 1441 619 1475
rect 653 1441 1359 1475
rect -124 1435 1359 1441
rect 2187 1415 2239 1421
rect -108 1401 1359 1407
rect -108 1367 -96 1401
rect -62 1367 -24 1401
rect 10 1367 999 1401
rect 1033 1367 1071 1401
rect 1105 1367 1359 1401
rect -108 1361 1359 1367
tri 2184 1361 2187 1364 se
rect 2187 1361 2239 1363
tri 2239 1361 2242 1364 sw
tri 2162 1339 2184 1361 se
rect 2184 1351 2242 1361
rect 2184 1339 2187 1351
rect 1731 1333 2187 1339
rect 2239 1339 2242 1351
tri 2242 1339 2264 1361 sw
rect 2239 1333 2437 1339
rect 1731 1299 1743 1333
rect 1777 1299 1815 1333
rect 1849 1299 1887 1333
rect 1921 1299 1959 1333
rect 1993 1299 2031 1333
rect 2065 1299 2103 1333
rect 2137 1299 2175 1333
rect 2239 1299 2247 1333
rect 2281 1299 2319 1333
rect 2353 1299 2391 1333
rect 2425 1299 2437 1333
rect 1731 1293 2437 1299
rect -520 1259 2877 1265
rect -520 1253 712 1259
rect -520 1219 -350 1253
rect -316 1225 712 1253
rect 746 1225 784 1259
rect 818 1225 1164 1259
rect 1198 1225 1301 1259
rect 1335 1225 1422 1259
rect 1456 1225 1540 1259
rect 1574 1253 2877 1259
rect 1574 1225 1642 1253
rect -316 1219 1642 1225
rect 1676 1251 2877 1253
rect 1676 1219 2667 1251
rect -520 1217 2667 1219
rect 2701 1217 2793 1251
rect 2827 1217 2877 1251
rect -520 1181 2877 1217
rect -520 1147 -350 1181
rect -316 1147 712 1181
rect 746 1147 784 1181
rect 818 1147 1164 1181
rect 1198 1147 1301 1181
rect 1335 1147 1422 1181
rect 1456 1147 1540 1181
rect 1574 1147 1642 1181
rect 1676 1147 2877 1181
rect -520 1110 2877 1147
rect -520 1103 2667 1110
rect -520 1069 712 1103
rect 746 1069 784 1103
rect 818 1069 1164 1103
rect 1198 1069 1301 1103
rect 1335 1069 1422 1103
rect 1456 1069 1540 1103
rect 1574 1076 2667 1103
rect 2701 1076 2793 1110
rect 2827 1076 2877 1110
rect 1574 1069 2877 1076
rect -520 1063 2877 1069
rect -528 919 -522 1035
rect -406 1023 241 1035
rect -406 989 -311 1023
rect -277 989 -143 1023
rect -109 989 33 1023
rect 67 989 201 1023
rect 235 989 241 1023
rect -406 951 241 989
rect -406 919 -311 951
rect -528 917 -311 919
rect -277 917 -143 951
rect -109 917 33 951
rect 67 917 201 951
rect 235 917 241 951
rect -528 905 241 917
rect 2187 1027 2239 1035
rect 2187 963 2239 975
rect 2187 905 2239 911
rect -597 871 1718 877
rect -597 837 -585 871
rect -551 837 -513 871
rect -479 837 -263 871
rect -229 837 -191 871
rect -157 837 47 871
rect 81 837 119 871
rect 153 837 1718 871
rect -597 825 1718 837
rect 1770 825 1782 877
rect 1834 825 1840 877
rect -711 656 2606 668
rect -711 622 -705 656
rect -671 622 -409 656
rect -375 622 -57 656
rect -23 622 294 656
rect 328 622 411 656
rect 445 622 2606 656
rect -711 584 2606 622
rect -711 550 -705 584
rect -671 550 -409 584
rect -375 550 -57 584
rect -23 550 294 584
rect 328 550 411 584
rect 445 550 2606 584
rect -711 538 2606 550
<< via1 >>
rect -522 1819 -470 1871
rect -458 1819 -406 1871
rect 1718 1555 1770 1561
rect 1718 1521 1722 1555
rect 1722 1521 1756 1555
rect 1756 1521 1770 1555
rect 1718 1509 1770 1521
rect 1782 1555 1834 1561
rect 1782 1521 1794 1555
rect 1794 1521 1828 1555
rect 1828 1521 1834 1555
rect 1782 1509 1834 1521
rect 2187 1363 2239 1415
rect 2187 1333 2239 1351
rect 2187 1299 2209 1333
rect 2209 1299 2239 1333
rect -522 919 -406 1035
rect 2187 975 2239 1027
rect 2187 911 2239 963
rect 1718 825 1770 877
rect 1782 825 1834 877
<< metal2 >>
rect -528 1819 -522 1871
rect -470 1819 -458 1871
rect -406 1819 -400 1871
rect -528 1035 -400 1819
rect -528 919 -522 1035
rect -406 919 -400 1035
rect 1712 1509 1718 1561
rect 1770 1509 1782 1561
rect 1834 1509 1840 1561
rect 1712 877 1840 1509
rect 2187 1415 2239 1421
rect 2187 1351 2239 1363
rect 2187 1027 2239 1299
rect 2187 963 2239 975
rect 2187 905 2239 911
rect 1712 825 1718 877
rect 1770 825 1782 877
rect 1834 825 1840 877
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_0
timestamp 1624884095
transform 1 0 -528 0 -1 1035
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_0
timestamp 1624884095
transform 0 -1 2239 1 0 1293
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_1
timestamp 1624884095
transform 0 -1 2239 1 0 905
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_2
timestamp 1624884095
transform 1 0 -528 0 1 1819
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_3
timestamp 1624884095
transform -1 0 1840 0 -1 1561
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_4
timestamp 1624884095
transform 1 0 1712 0 1 825
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808294  sky130_fd_pr__via_pol1__example_55959141808294_0
timestamp 1624884095
transform 0 -1 368 -1 0 1906
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_0
timestamp 1624884095
transform 0 -1 2465 -1 0 1282
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_1
timestamp 1624884095
transform 0 -1 2448 1 0 1840
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808349  sky130_fd_pr__via_l1m1__example_55959141808349_0
timestamp 1624884095
transform 1 0 1743 0 1 1299
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808290  sky130_fd_pr__via_l1m1__example_55959141808290_0
timestamp 1624884095
transform 1 0 -174 0 1 1825
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808326  sky130_fd_pr__via_l1m1__example_55959141808326_0
timestamp 1624884095
transform -1 0 2464 0 1 1825
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1624884095
transform 0 -1 -277 1 0 917
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1624884095
transform 0 1 294 -1 0 656
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1624884095
transform 0 -1 -109 1 0 917
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1624884095
transform 0 1 411 -1 0 656
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_4
timestamp 1624884095
transform 1 0 320 0 1 1521
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_5
timestamp 1624884095
transform 0 -1 67 1 0 917
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_6
timestamp 1624884095
transform 0 -1 235 1 0 917
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_7
timestamp 1624884095
transform 0 -1 1676 1 0 1147
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_8
timestamp 1624884095
transform 1 0 1722 0 1 1521
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_9
timestamp 1624884095
transform 1 0 43 0 1 1521
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_10
timestamp 1624884095
transform -1 0 10 0 1 1367
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_11
timestamp 1624884095
transform -1 0 1105 0 1 1367
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_12
timestamp 1624884095
transform -1 0 306 0 1 1441
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_13
timestamp 1624884095
transform 1 0 -234 0 1 1521
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_14
timestamp 1624884095
transform -1 0 653 0 1 1441
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_15
timestamp 1624884095
transform -1 0 153 0 1 837
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_16
timestamp 1624884095
transform -1 0 -157 0 1 837
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_17
timestamp 1624884095
transform -1 0 -479 0 1 837
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_18
timestamp 1624884095
transform 0 1 -705 -1 0 656
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_19
timestamp 1624884095
transform 0 1 -409 -1 0 656
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_20
timestamp 1624884095
transform 0 1 -57 -1 0 656
box 0 0 1 1
use sky130_fd_pr__pfet_01v8__example_55959141808356  sky130_fd_pr__pfet_01v8__example_55959141808356_0
timestamp 1624884095
transform 1 0 1687 0 1 1314
box -28 0 828 97
use sky130_fd_pr__pfet_01v8__example_55959141808356  sky130_fd_pr__pfet_01v8__example_55959141808356_1
timestamp 1624884095
transform -1 0 2487 0 -1 1808
box -28 0 828 97
use sky130_fd_pr__pfet_01v8__example_55959141808355  sky130_fd_pr__pfet_01v8__example_55959141808355_0
timestamp 1624884095
transform 1 0 123 0 1 1208
box -28 0 284 267
use sky130_fd_pr__pfet_01v8__example_55959141808355  sky130_fd_pr__pfet_01v8__example_55959141808355_1
timestamp 1624884095
transform -1 0 67 0 1 1208
box -28 0 284 267
use sky130_fd_pr__pfet_01v8__example_55959141808354  sky130_fd_pr__pfet_01v8__example_55959141808354_0
timestamp 1624884095
transform 0 -1 2761 -1 0 1748
box -28 0 828 29
use sky130_fd_pr__pfet_01v8__example_55959141808353  sky130_fd_pr__pfet_01v8__example_55959141808353_0
timestamp 1624884095
transform 1 0 809 0 1 1118
box -28 0 228 97
use sky130_fd_pr__pfet_01v8__example_55959141808353  sky130_fd_pr__pfet_01v8__example_55959141808353_1
timestamp 1624884095
transform -1 0 1265 0 1 1118
box -28 0 228 97
use sky130_fd_pr__pfet_01v8__example_55959141808353  sky130_fd_pr__pfet_01v8__example_55959141808353_2
timestamp 1624884095
transform 1 0 809 0 -1 1808
box -28 0 228 97
use sky130_fd_pr__pfet_01v8__example_55959141808353  sky130_fd_pr__pfet_01v8__example_55959141808353_3
timestamp 1624884095
transform -1 0 1265 0 -1 1808
box -28 0 228 97
use sky130_fd_pr__pfet_01v8__example_55959141808352  sky130_fd_pr__pfet_01v8__example_55959141808352_0
timestamp 1624884095
transform -1 0 753 0 1 1118
box -28 0 128 97
use sky130_fd_pr__pfet_01v8__example_55959141808352  sky130_fd_pr__pfet_01v8__example_55959141808352_1
timestamp 1624884095
transform -1 0 753 0 -1 1808
box -28 0 128 97
use sky130_fd_pr__nfet_01v8__example_55959141808351  sky130_fd_pr__nfet_01v8__example_55959141808351_0
timestamp 1624884095
transform -1 0 284 0 1 426
box -28 0 852 267
<< labels >>
flabel locali s 1190 979 1236 1013 0 FreeSans 300 180 0 0 EN_FAST_N[1]
port 1 nsew
flabel metal1 s 2564 1589 2606 1791 7 FreeSans 300 180 0 0 VGND_IO
port 2 nsew
flabel metal1 s -520 1589 -478 1791 3 FreeSans 300 180 0 0 VGND_IO
port 2 nsew
flabel metal1 s 2187 905 2239 954 7 FreeSans 300 180 0 0 PDEN_H_N
port 3 nsew
flabel metal1 s 1793 825 1840 877 7 FreeSans 300 180 0 0 PD_H
port 4 nsew
flabel metal1 s -528 1819 -481 1871 3 FreeSans 300 180 0 0 DRVLO_H_N
port 5 nsew
flabel metal1 s 2564 538 2606 668 7 FreeSans 300 180 0 0 VGND_IO
port 2 nsew
flabel metal1 s -516 538 -474 668 3 FreeSans 300 180 0 0 VGND_IO
port 2 nsew
flabel metal1 s -520 1063 -480 1265 3 FreeSans 300 180 0 0 VCC_IO
port 6 nsew
flabel metal1 s 2837 1063 2877 1265 7 FreeSans 300 180 0 0 VCC_IO
port 6 nsew
flabel comment s 2114 1228 2114 1228 0 FreeSans 300 0 0 0 PDEN_H_N
flabel comment s 20 1142 20 1142 0 FreeSans 300 0 0 0 DRVLO_H_N
flabel comment s 42 1547 42 1547 0 FreeSans 300 0 0 0 PD_H
flabel comment s -201 861 -201 861 0 FreeSans 300 0 0 0 PD_H
flabel comment s 2071 1905 2071 1905 0 FreeSans 300 0 0 0 DRVLO_H_N
flabel comment s 1236 1009 1236 1009 0 FreeSans 300 0 0 0 EN_FAST_N[1]
flabel comment s 761 1890 761 1890 0 FreeSans 300 0 0 0 EN_FAST_N<0>
flabel comment s 2512 1553 2512 1553 0 FreeSans 300 90 0 0 INT_SLOW
flabel comment s 366 1122 366 1122 0 FreeSans 300 0 0 0 PDEN_H_N
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 36974220
string GDS_START 36956782
<< end >>
