magic
tech sky130A
magscale 1 2
timestamp 1624884095
<< checkpaint >>
rect -1245 -1247 1545 1274
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_0
timestamp 1624884095
transform -1 0 16 0 1 13
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_1
timestamp 1624884095
transform 1 0 284 0 1 13
box 0 0 1 1
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 39006
string GDS_START 38524
<< end >>
