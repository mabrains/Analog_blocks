magic
tech sky130A
magscale 1 2
timestamp 1624884095
<< checkpaint >>
rect -1288 -1260 1544 1391
use sky130_fd_pr__dfl1sd__example_55959141808504  sky130_fd_pr__dfl1sd__example_55959141808504_0
timestamp 1624884095
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808462  sky130_fd_pr__hvdfl1sd2__example_55959141808462_0
timestamp 1624884095
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808278  sky130_fd_pr__hvdfl1sd__example_55959141808278_0
timestamp 1624884095
transform -1 0 0 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 284 131 284 131 0 FreeSans 300 0 0 0 S
flabel comment s 128 131 128 131 0 FreeSans 300 0 0 0 D
flabel comment s -28 131 -28 131 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 48364024
string GDS_START 48362582
<< end >>
