magic
tech sky130A
magscale 1 2
timestamp 1624884114
<< metal3 >>
rect 11966 18347 14932 18592
rect 11788 18333 11966 18347
rect 11982 18333 14932 18347
rect 11788 18169 14932 18333
rect 11530 18153 11788 18169
rect 11802 18153 14932 18169
rect 11530 17911 14932 18153
rect 11283 17883 11530 17911
rect 11532 17883 14932 17911
rect 11283 17664 14932 17883
rect 11027 17643 11283 17664
rect 11292 17643 14932 17664
rect 11027 17408 14932 17643
rect 10742 17403 11027 17408
rect 11052 17403 14932 17408
rect 10742 17123 14932 17403
rect 10481 17103 10742 17123
rect 10752 17103 14932 17123
rect 10481 16862 14932 17103
rect 10152 16833 10481 16862
rect 10482 16833 14932 16862
rect 10152 13607 14932 16833
rect 10151 12418 14931 13306
rect 120 3558 4900 4486
rect 10151 3558 14931 4486
<< obsm3 >>
rect 119 18427 11886 18591
rect 119 18249 11708 18427
rect 119 17991 11450 18249
rect 119 17744 11203 17991
rect 119 17488 10947 17744
rect 119 17203 10662 17488
rect 119 16942 10401 17203
rect 119 13527 10072 16942
rect 119 13386 11982 13527
rect 119 12418 10071 13386
<< metal4 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 0 18592 254 18600
rect 0 16558 2821 18592
rect 14746 18593 15000 18600
rect 2851 18190 3073 18342
rect 2854 17669 3250 18164
rect 11978 18190 12200 18342
rect 3283 17673 3505 17906
rect 2875 16598 3771 17628
rect 11546 17673 11768 17906
rect 11801 17669 12197 18164
rect 3799 17162 4013 17403
rect 3834 16589 4290 17118
rect 11038 17162 11252 17403
rect 4330 16571 4554 16857
rect 0 16525 254 16558
rect 0 13612 4900 16525
rect 0 13607 254 13612
rect 10497 16571 10721 16857
rect 10761 16589 11217 17118
rect 11280 16598 12176 17628
rect 12230 16557 15000 18593
rect 14746 16525 15000 16557
rect 10151 13612 15000 16525
rect 14746 13607 15000 13612
rect 0 12417 4895 13307
rect 10156 12417 15000 13307
rect 0 11247 254 12137
rect 14746 11247 15000 12137
rect 0 10881 15000 10947
rect 0 10225 15000 10821
rect 0 9929 254 10165
rect 14746 9929 15000 10165
rect 0 9273 15000 9869
rect 0 9147 15000 9213
rect 0 7917 254 8847
rect 14746 7917 15000 8847
rect 0 6947 254 7637
rect 14746 6947 15000 7637
rect 0 5977 254 6667
rect 14746 5977 15000 6667
rect 0 4767 254 5697
rect 14746 4767 15000 5697
rect 0 3557 4895 4487
rect 10156 3557 15000 4487
rect 0 2587 193 3277
rect 14807 2587 15000 3277
rect 0 1377 254 2307
rect 14746 1377 15000 2307
rect 0 7 254 1097
rect 14746 7 15000 1097
<< obsm4 >>
rect 334 34677 14666 39600
rect 193 18680 14807 34677
rect 334 18673 14666 18680
rect 334 18672 12150 18673
rect 2901 18422 12150 18672
rect 3153 18244 11898 18422
rect 3330 17986 11721 18244
rect 3585 17708 11466 17986
rect 3851 17483 11200 17708
rect 4093 17198 10958 17483
rect 4370 16937 10681 17198
rect 4634 16605 10417 16937
rect 4980 13532 10071 16605
rect 334 13527 14666 13532
rect 193 13387 14807 13527
rect 4975 12337 10076 13387
rect 193 12217 14807 12337
rect 334 11167 14666 12217
rect 193 11027 14807 11167
rect 334 9949 14666 10145
rect 193 8927 14807 9067
rect 334 7837 14666 8927
rect 193 7717 14807 7837
rect 334 6867 14666 7717
rect 193 6747 14807 6867
rect 334 5897 14666 6747
rect 193 5777 14807 5897
rect 334 4687 14666 5777
rect 193 4567 14807 4687
rect 4975 3477 10076 4567
rect 193 3357 14807 3477
rect 273 2507 14727 3357
rect 193 2387 14807 2507
rect 334 1297 14666 2387
rect 193 1177 14807 1297
rect 334 7 14666 1177
<< metal5 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 0 13607 254 18597
rect 0 12437 254 13287
rect 0 11267 254 12117
rect 0 9147 254 10947
rect 0 7937 254 8827
rect 0 6968 254 7617
rect 14746 13607 15000 18597
rect 14746 12437 15000 13287
rect 14746 11267 15000 12117
rect 14746 9147 15000 10947
rect 14746 7937 15000 8827
rect 14746 6968 15000 7617
rect 0 5997 254 6647
rect 0 4787 254 5677
rect 0 3577 254 4467
rect 14746 5997 15000 6647
rect 14746 4787 15000 5677
rect 14746 3577 15000 4467
rect 0 2607 193 3257
rect 14807 2607 15000 3257
rect 0 1397 254 2287
rect 0 27 254 1077
rect 14746 1397 15000 2287
rect 14746 27 15000 1077
<< obsm5 >>
rect 574 34437 14426 39600
rect 0 18917 15000 34437
rect 574 6968 14426 18917
rect 0 6967 15000 6968
rect 574 3257 14426 6967
rect 513 2607 14487 3257
rect 574 27 14426 2607
<< labels >>
rlabel metal5 s 14746 12437 15000 13287 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal5 s 0 12437 254 13287 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 0 12417 254 13307 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 14746 12417 15000 13307 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10151 12418 14931 13306 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 0 12417 4895 13307 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10156 12417 15000 13307 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal5 s 0 12437 254 13287 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal5 s 14746 12437 15000 13287 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 13252 14913 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 13170 14913 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 13088 14913 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 13006 14913 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 12924 14913 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 12842 14913 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 12760 14913 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 12678 14913 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 12596 14913 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 12514 14913 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 12432 14913 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 13252 14831 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 13170 14831 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 13088 14831 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 13006 14831 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 12924 14831 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 12842 14831 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 12760 14831 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 12678 14831 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 12596 14831 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 12514 14831 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 12432 14831 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 13252 14749 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 13170 14749 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 13088 14749 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 13006 14749 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 12924 14749 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 12842 14749 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 12760 14749 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 12678 14749 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 12596 14749 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 12514 14749 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 12432 14749 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 13252 14667 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 13170 14667 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 13088 14667 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 13006 14667 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 12924 14667 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 12842 14667 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 12760 14667 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 12678 14667 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 12596 14667 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 12514 14667 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 12432 14667 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 13252 14585 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 13170 14585 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 13088 14585 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 13006 14585 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 12924 14585 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 12842 14585 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 12760 14585 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 12678 14585 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 12596 14585 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 12514 14585 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 12432 14585 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 13252 14503 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 13170 14503 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 13088 14503 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 13006 14503 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 12924 14503 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 12842 14503 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 12760 14503 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 12678 14503 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 12596 14503 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 12514 14503 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 12432 14503 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 13252 14421 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 13170 14421 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 13088 14421 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 13006 14421 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 12924 14421 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 12842 14421 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 12760 14421 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 12678 14421 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 12596 14421 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 12514 14421 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 12432 14421 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 13252 14340 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 13170 14340 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 13088 14340 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 13006 14340 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 12924 14340 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 12842 14340 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 12760 14340 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 12678 14340 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 12596 14340 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 12514 14340 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 12432 14340 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 13252 14259 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 13170 14259 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 13088 14259 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 13006 14259 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 12924 14259 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 12842 14259 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 12760 14259 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 12678 14259 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 12596 14259 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 12514 14259 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 12432 14259 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 13252 14178 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 13170 14178 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 13088 14178 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 13006 14178 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 12924 14178 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 12842 14178 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 12760 14178 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 12678 14178 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 12596 14178 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 12514 14178 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 12432 14178 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 13252 14097 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 13170 14097 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 13088 14097 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 13006 14097 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 12924 14097 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 12842 14097 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 12760 14097 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 12678 14097 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 12596 14097 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 12514 14097 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 12432 14097 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 13252 14016 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 13170 14016 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 13088 14016 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 13006 14016 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 12924 14016 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 12842 14016 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 12760 14016 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 12678 14016 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 12596 14016 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 12514 14016 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 12432 14016 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 13252 13935 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 13170 13935 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 13088 13935 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 13006 13935 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 12924 13935 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 12842 13935 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 12760 13935 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 12678 13935 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 12596 13935 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 12514 13935 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 12432 13935 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 13252 13854 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 13170 13854 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 13088 13854 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 13006 13854 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 12924 13854 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 12842 13854 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 12760 13854 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 12678 13854 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 12596 13854 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 12514 13854 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 12432 13854 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 13252 13773 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 13170 13773 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 13088 13773 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 13006 13773 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 12924 13773 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 12842 13773 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 12760 13773 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 12678 13773 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 12596 13773 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 12514 13773 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 12432 13773 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 13252 13692 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 13170 13692 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 13088 13692 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 13006 13692 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 12924 13692 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 12842 13692 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 12760 13692 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 12678 13692 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 12596 13692 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 12514 13692 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 12432 13692 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 13252 13611 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 13170 13611 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 13088 13611 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 13006 13611 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 12924 13611 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 12842 13611 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 12760 13611 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 12678 13611 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 12596 13611 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 12514 13611 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 12432 13611 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 13252 13530 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 13170 13530 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 13088 13530 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 13006 13530 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 12924 13530 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 12842 13530 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 12760 13530 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 12678 13530 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 12596 13530 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 12514 13530 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 12432 13530 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 13252 13449 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 13170 13449 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 13088 13449 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 13006 13449 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 12924 13449 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 12842 13449 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 12760 13449 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 12678 13449 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 12596 13449 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 12514 13449 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 12432 13449 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 13252 13368 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 13170 13368 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 13088 13368 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 13006 13368 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 12924 13368 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 12842 13368 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 12760 13368 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 12678 13368 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 12596 13368 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 12514 13368 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 12432 13368 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 13252 13287 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 13170 13287 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 13088 13287 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 13006 13287 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 12924 13287 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 12842 13287 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 12760 13287 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 12678 13287 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 12596 13287 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 12514 13287 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 12432 13287 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 13252 13206 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 13170 13206 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 13088 13206 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 13006 13206 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 12924 13206 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 12842 13206 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 12760 13206 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 12678 13206 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 12596 13206 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 12514 13206 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 12432 13206 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 13252 13125 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 13170 13125 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 13088 13125 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 13006 13125 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 12924 13125 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 12842 13125 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 12760 13125 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 12678 13125 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 12596 13125 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 12514 13125 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 12432 13125 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 13252 13044 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 13170 13044 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 13088 13044 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 13006 13044 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 12924 13044 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 12842 13044 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 12760 13044 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 12678 13044 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 12596 13044 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 12514 13044 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 12432 13044 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 13252 12963 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 13170 12963 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 13088 12963 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 13006 12963 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 12924 12963 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 12842 12963 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 12760 12963 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 12678 12963 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 12596 12963 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 12514 12963 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 12432 12963 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 13252 12882 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 13170 12882 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 13088 12882 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 13006 12882 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 12924 12882 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 12842 12882 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 12760 12882 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 12678 12882 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 12596 12882 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 12514 12882 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 12432 12882 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 13252 12801 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 13170 12801 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 13088 12801 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 13006 12801 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 12924 12801 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 12842 12801 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 12760 12801 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 12678 12801 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 12596 12801 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 12514 12801 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 12432 12801 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 13252 12720 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 13170 12720 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 13088 12720 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 13006 12720 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 12924 12720 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 12842 12720 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 12760 12720 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 12678 12720 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 12596 12720 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 12514 12720 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 12432 12720 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 13252 12639 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 13170 12639 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 13088 12639 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 13006 12639 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 12924 12639 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 12842 12639 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 12760 12639 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 12678 12639 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 12596 12639 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 12514 12639 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 12432 12639 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 13252 12558 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 13170 12558 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 13088 12558 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 13006 12558 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 12924 12558 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 12842 12558 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 12760 12558 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 12678 12558 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 12596 12558 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 12514 12558 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 12432 12558 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 13252 12477 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 13170 12477 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 13088 12477 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 13006 12477 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 12924 12477 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 12842 12477 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 12760 12477 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 12678 12477 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 12596 12477 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 12514 12477 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 12432 12477 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 13252 12396 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 13170 12396 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 13088 12396 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 13006 12396 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 12924 12396 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 12842 12396 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 12760 12396 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 12678 12396 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 12596 12396 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 12514 12396 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 12432 12396 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 13252 12315 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 13170 12315 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 13088 12315 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 13006 12315 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 12924 12315 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 12842 12315 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 12760 12315 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 12678 12315 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 12596 12315 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 12514 12315 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 12432 12315 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 13252 12234 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 13170 12234 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 13088 12234 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 13006 12234 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 12924 12234 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 12842 12234 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 12760 12234 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 12678 12234 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 12596 12234 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 12514 12234 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 12432 12234 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 13252 12153 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 13170 12153 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 13088 12153 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 13006 12153 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 12924 12153 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 12842 12153 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 12760 12153 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 12678 12153 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 12596 12153 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 12514 12153 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 12432 12153 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 13252 12072 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 13170 12072 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 13088 12072 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 13006 12072 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 12924 12072 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 12842 12072 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 12760 12072 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 12678 12072 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 12596 12072 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 12514 12072 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 12432 12072 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 13252 11991 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 13170 11991 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 13088 11991 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 13006 11991 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 12924 11991 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 12842 11991 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 12760 11991 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 12678 11991 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 12596 11991 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 12514 11991 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 12432 11991 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 13252 11910 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 13170 11910 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 13088 11910 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 13006 11910 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 12924 11910 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 12842 11910 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 12760 11910 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 12678 11910 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 12596 11910 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 12514 11910 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 12432 11910 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 13252 11829 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 13170 11829 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 13088 11829 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 13006 11829 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 12924 11829 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 12842 11829 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 12760 11829 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 12678 11829 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 12596 11829 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 12514 11829 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 12432 11829 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 13252 11748 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 13170 11748 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 13088 11748 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 13006 11748 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 12924 11748 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 12842 11748 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 12760 11748 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 12678 11748 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 12596 11748 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 12514 11748 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 12432 11748 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 13252 11667 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 13170 11667 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 13088 11667 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 13006 11667 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 12924 11667 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 12842 11667 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 12760 11667 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 12678 11667 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 12596 11667 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 12514 11667 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 12432 11667 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 13252 11586 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 13170 11586 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 13088 11586 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 13006 11586 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 12924 11586 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 12842 11586 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 12760 11586 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 12678 11586 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 12596 11586 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 12514 11586 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 12432 11586 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 13252 11505 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 13170 11505 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 13088 11505 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 13006 11505 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 12924 11505 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 12842 11505 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 12760 11505 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 12678 11505 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 12596 11505 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 12514 11505 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 12432 11505 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 13252 11424 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 13170 11424 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 13088 11424 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 13006 11424 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 12924 11424 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 12842 11424 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 12760 11424 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 12678 11424 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 12596 11424 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 12514 11424 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 12432 11424 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 13252 11343 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 13170 11343 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 13088 11343 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 13006 11343 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 12924 11343 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 12842 11343 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 12760 11343 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 12678 11343 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 12596 11343 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 12514 11343 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 12432 11343 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 13252 11262 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 13170 11262 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 13088 11262 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 13006 11262 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 12924 11262 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 12842 11262 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 12760 11262 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 12678 11262 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 12596 11262 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 12514 11262 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 12432 11262 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 13252 11181 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 13170 11181 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 13088 11181 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 13006 11181 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 12924 11181 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 12842 11181 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 12760 11181 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 12678 11181 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 12596 11181 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 12514 11181 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 12432 11181 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 13252 11100 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 13170 11100 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 13088 11100 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 13006 11100 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 12924 11100 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 12842 11100 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 12760 11100 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 12678 11100 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 12596 11100 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 12514 11100 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 12432 11100 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 13252 11019 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 13170 11019 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 13088 11019 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 13006 11019 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 12924 11019 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 12842 11019 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 12760 11019 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 12678 11019 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 12596 11019 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 12514 11019 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 12432 11019 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 13252 10938 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 13170 10938 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 13088 10938 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 13006 10938 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 12924 10938 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 12842 10938 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 12760 10938 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 12678 10938 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 12596 10938 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 12514 10938 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 12432 10938 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 13252 10857 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 13170 10857 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 13088 10857 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 13006 10857 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 12924 10857 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 12842 10857 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 12760 10857 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 12678 10857 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 12596 10857 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 12514 10857 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 12432 10857 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 13252 10776 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 13170 10776 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 13088 10776 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 13006 10776 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 12924 10776 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 12842 10776 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 12760 10776 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 12678 10776 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 12596 10776 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 12514 10776 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 12432 10776 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 13252 10695 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 13170 10695 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 13088 10695 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 13006 10695 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 12924 10695 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 12842 10695 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 12760 10695 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 12678 10695 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 12596 10695 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 12514 10695 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 12432 10695 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 13252 10614 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 13170 10614 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 13088 10614 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 13006 10614 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 12924 10614 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 12842 10614 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 12760 10614 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 12678 10614 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 12596 10614 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 12514 10614 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 12432 10614 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 13252 10533 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 13170 10533 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 13088 10533 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 13006 10533 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 12924 10533 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 12842 10533 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 12760 10533 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 12678 10533 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 12596 10533 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 12514 10533 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 12432 10533 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 13252 10452 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 13170 10452 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 13088 10452 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 13006 10452 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 12924 10452 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 12842 10452 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 12760 10452 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 12678 10452 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 12596 10452 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 12514 10452 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 12432 10452 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 13252 10371 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 13170 10371 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 13088 10371 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 13006 10371 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 12924 10371 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 12842 10371 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 12760 10371 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 12678 10371 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 12596 10371 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 12514 10371 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 12432 10371 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 13252 10290 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 13170 10290 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 13088 10290 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 13006 10290 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 12924 10290 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 12842 10290 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 12760 10290 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 12678 10290 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 12596 10290 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 12514 10290 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 12432 10290 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 13252 10209 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 13170 10209 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 13088 10209 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 13006 10209 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 12924 10209 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 12842 10209 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 12760 10209 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 12678 10209 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 12596 10209 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 12514 10209 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 12432 10209 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 13240 4894 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 13158 4894 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 13076 4894 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 12994 4894 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 12912 4894 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 12830 4894 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 12748 4894 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 12666 4894 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 12584 4894 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 12502 4894 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4830 12420 4894 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 13240 4812 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 13158 4812 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 13076 4812 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 12994 4812 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 12912 4812 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 12830 4812 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 12748 4812 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 12666 4812 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 12584 4812 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 12502 4812 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4748 12420 4812 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 13240 4730 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 13158 4730 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 13076 4730 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 12994 4730 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 12912 4730 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 12830 4730 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 12748 4730 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 12666 4730 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 12584 4730 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 12502 4730 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4666 12420 4730 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 13240 4648 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 13158 4648 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 13076 4648 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 12994 4648 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 12912 4648 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 12830 4648 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 12748 4648 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 12666 4648 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 12584 4648 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 12502 4648 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4584 12420 4648 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 13240 4566 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 13158 4566 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 13076 4566 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 12994 4566 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 12912 4566 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 12830 4566 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 12748 4566 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 12666 4566 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 12584 4566 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 12502 4566 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4502 12420 4566 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 13240 4484 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 13158 4484 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 13076 4484 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 12994 4484 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 12912 4484 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 12830 4484 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 12748 4484 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 12666 4484 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 12584 4484 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 12502 4484 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4420 12420 4484 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 13240 4402 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 13158 4402 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 13076 4402 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 12994 4402 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 12912 4402 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 12830 4402 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 12748 4402 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 12666 4402 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 12584 4402 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 12502 4402 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4338 12420 4402 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 13240 4321 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 13158 4321 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 13076 4321 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 12994 4321 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 12912 4321 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 12830 4321 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 12748 4321 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 12666 4321 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 12584 4321 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 12502 4321 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4257 12420 4321 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 13240 4240 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 13158 4240 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 13076 4240 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 12994 4240 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 12912 4240 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 12830 4240 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 12748 4240 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 12666 4240 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 12584 4240 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 12502 4240 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4176 12420 4240 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 13240 4159 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 13158 4159 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 13076 4159 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 12994 4159 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 12912 4159 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 12830 4159 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 12748 4159 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 12666 4159 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 12584 4159 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 12502 4159 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4095 12420 4159 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 13240 4078 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 13158 4078 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 13076 4078 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 12994 4078 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 12912 4078 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 12830 4078 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 12748 4078 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 12666 4078 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 12584 4078 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 12502 4078 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4014 12420 4078 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 13240 3997 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 13158 3997 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 13076 3997 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 12994 3997 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 12912 3997 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 12830 3997 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 12748 3997 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 12666 3997 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 12584 3997 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 12502 3997 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3933 12420 3997 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 13240 3916 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 13158 3916 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 13076 3916 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 12994 3916 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 12912 3916 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 12830 3916 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 12748 3916 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 12666 3916 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 12584 3916 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 12502 3916 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3852 12420 3916 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 13240 3835 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 13158 3835 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 13076 3835 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 12994 3835 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 12912 3835 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 12830 3835 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 12748 3835 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 12666 3835 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 12584 3835 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 12502 3835 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3771 12420 3835 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 13240 3754 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 13158 3754 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 13076 3754 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 12994 3754 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 12912 3754 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 12830 3754 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 12748 3754 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 12666 3754 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 12584 3754 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 12502 3754 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3690 12420 3754 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 13240 3673 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 13158 3673 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 13076 3673 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 12994 3673 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 12912 3673 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 12830 3673 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 12748 3673 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 12666 3673 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 12584 3673 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 12502 3673 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3609 12420 3673 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 13240 3592 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 13158 3592 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 13076 3592 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 12994 3592 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 12912 3592 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 12830 3592 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 12748 3592 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 12666 3592 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 12584 3592 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 12502 3592 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3528 12420 3592 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 13240 3511 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 13158 3511 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 13076 3511 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 12994 3511 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 12912 3511 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 12830 3511 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 12748 3511 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 12666 3511 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 12584 3511 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 12502 3511 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3447 12420 3511 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 13240 3430 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 13158 3430 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 13076 3430 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 12994 3430 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 12912 3430 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 12830 3430 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 12748 3430 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 12666 3430 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 12584 3430 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 12502 3430 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3366 12420 3430 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 13240 3349 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 13158 3349 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 13076 3349 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 12994 3349 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 12912 3349 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 12830 3349 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 12748 3349 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 12666 3349 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 12584 3349 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 12502 3349 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3285 12420 3349 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 13240 3268 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 13158 3268 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 13076 3268 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 12994 3268 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 12912 3268 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 12830 3268 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 12748 3268 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 12666 3268 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 12584 3268 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 12502 3268 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3204 12420 3268 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 13240 3187 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 13158 3187 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 13076 3187 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 12994 3187 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 12912 3187 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 12830 3187 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 12748 3187 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 12666 3187 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 12584 3187 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 12502 3187 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3123 12420 3187 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 13240 3106 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 13158 3106 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 13076 3106 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 12994 3106 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 12912 3106 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 12830 3106 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 12748 3106 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 12666 3106 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 12584 3106 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 12502 3106 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3042 12420 3106 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 13240 3025 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 13158 3025 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 13076 3025 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 12994 3025 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 12912 3025 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 12830 3025 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 12748 3025 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 12666 3025 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 12584 3025 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 12502 3025 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2961 12420 3025 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 13240 2944 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 13158 2944 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 13076 2944 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 12994 2944 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 12912 2944 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 12830 2944 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 12748 2944 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 12666 2944 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 12584 2944 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 12502 2944 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2880 12420 2944 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 13240 2863 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 13158 2863 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 13076 2863 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 12994 2863 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 12912 2863 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 12830 2863 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 12748 2863 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 12666 2863 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 12584 2863 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 12502 2863 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2799 12420 2863 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 13240 2782 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 13158 2782 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 13076 2782 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 12994 2782 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 12912 2782 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 12830 2782 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 12748 2782 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 12666 2782 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 12584 2782 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 12502 2782 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2718 12420 2782 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 13240 2701 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 13158 2701 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 13076 2701 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 12994 2701 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 12912 2701 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 12830 2701 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 12748 2701 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 12666 2701 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 12584 2701 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 12502 2701 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2637 12420 2701 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 13240 2620 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 13158 2620 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 13076 2620 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 12994 2620 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 12912 2620 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 12830 2620 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 12748 2620 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 12666 2620 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 12584 2620 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 12502 2620 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2556 12420 2620 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 13240 2539 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 13158 2539 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 13076 2539 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 12994 2539 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 12912 2539 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 12830 2539 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 12748 2539 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 12666 2539 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 12584 2539 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 12502 2539 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2475 12420 2539 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 13240 2458 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 13158 2458 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 13076 2458 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 12994 2458 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 12912 2458 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 12830 2458 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 12748 2458 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 12666 2458 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 12584 2458 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 12502 2458 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2394 12420 2458 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 13240 2377 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 13158 2377 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 13076 2377 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 12994 2377 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 12912 2377 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 12830 2377 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 12748 2377 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 12666 2377 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 12584 2377 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 12502 2377 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2313 12420 2377 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 13240 2296 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 13158 2296 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 13076 2296 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 12994 2296 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 12912 2296 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 12830 2296 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 12748 2296 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 12666 2296 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 12584 2296 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 12502 2296 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2232 12420 2296 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 13240 2215 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 13158 2215 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 13076 2215 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 12994 2215 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 12912 2215 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 12830 2215 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 12748 2215 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 12666 2215 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 12584 2215 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 12502 2215 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2151 12420 2215 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 13240 2134 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 13158 2134 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 13076 2134 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 12994 2134 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 12912 2134 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 12830 2134 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 12748 2134 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 12666 2134 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 12584 2134 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 12502 2134 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2070 12420 2134 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 13240 2053 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 13158 2053 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 13076 2053 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 12994 2053 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 12912 2053 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 12830 2053 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 12748 2053 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 12666 2053 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 12584 2053 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 12502 2053 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1989 12420 2053 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 13240 1972 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 13158 1972 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 13076 1972 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 12994 1972 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 12912 1972 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 12830 1972 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 12748 1972 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 12666 1972 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 12584 1972 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 12502 1972 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1908 12420 1972 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 13240 1891 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 13158 1891 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 13076 1891 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 12994 1891 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 12912 1891 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 12830 1891 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 12748 1891 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 12666 1891 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 12584 1891 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 12502 1891 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1827 12420 1891 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 13240 1810 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 13158 1810 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 13076 1810 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 12994 1810 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 12912 1810 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 12830 1810 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 12748 1810 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 12666 1810 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 12584 1810 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 12502 1810 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1746 12420 1810 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 13240 1729 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 13158 1729 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 13076 1729 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 12994 1729 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 12912 1729 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 12830 1729 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 12748 1729 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 12666 1729 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 12584 1729 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 12502 1729 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1665 12420 1729 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 13240 1648 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 13158 1648 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 13076 1648 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 12994 1648 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 12912 1648 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 12830 1648 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 12748 1648 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 12666 1648 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 12584 1648 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 12502 1648 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1584 12420 1648 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 13240 1567 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 13158 1567 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 13076 1567 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 12994 1567 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 12912 1567 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 12830 1567 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 12748 1567 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 12666 1567 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 12584 1567 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 12502 1567 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1503 12420 1567 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 13240 1486 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 13158 1486 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 13076 1486 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 12994 1486 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 12912 1486 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 12830 1486 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 12748 1486 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 12666 1486 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 12584 1486 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 12502 1486 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1422 12420 1486 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 13240 1405 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 13158 1405 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 13076 1405 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 12994 1405 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 12912 1405 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 12830 1405 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 12748 1405 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 12666 1405 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 12584 1405 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 12502 1405 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1341 12420 1405 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 13240 1324 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 13158 1324 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 13076 1324 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 12994 1324 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 12912 1324 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 12830 1324 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 12748 1324 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 12666 1324 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 12584 1324 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 12502 1324 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1260 12420 1324 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 13240 1243 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 13158 1243 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 13076 1243 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 12994 1243 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 12912 1243 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 12830 1243 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 12748 1243 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 12666 1243 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 12584 1243 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 12502 1243 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1179 12420 1243 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 13240 1162 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 13158 1162 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 13076 1162 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 12994 1162 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 12912 1162 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 12830 1162 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 12748 1162 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 12666 1162 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 12584 1162 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 12502 1162 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1098 12420 1162 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 13240 1081 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 13158 1081 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 13076 1081 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 12994 1081 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 12912 1081 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 12830 1081 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 12748 1081 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 12666 1081 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 12584 1081 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 12502 1081 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1017 12420 1081 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 13240 1000 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 13158 1000 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 13076 1000 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 12994 1000 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 12912 1000 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 12830 1000 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 12748 1000 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 12666 1000 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 12584 1000 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 12502 1000 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 936 12420 1000 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 13240 919 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 13158 919 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 13076 919 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 12994 919 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 12912 919 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 12830 919 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 12748 919 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 12666 919 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 12584 919 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 12502 919 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 855 12420 919 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 13240 838 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 13158 838 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 13076 838 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 12994 838 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 12912 838 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 12830 838 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 12748 838 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 12666 838 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 12584 838 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 12502 838 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 774 12420 838 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 13240 757 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 13158 757 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 13076 757 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 12994 757 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 12912 757 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 12830 757 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 12748 757 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 12666 757 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 12584 757 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 12502 757 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 693 12420 757 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 13240 676 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 13158 676 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 13076 676 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 12994 676 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 12912 676 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 12830 676 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 12748 676 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 12666 676 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 12584 676 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 12502 676 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 612 12420 676 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 13240 595 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 13158 595 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 13076 595 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 12994 595 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 12912 595 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 12830 595 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 12748 595 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 12666 595 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 12584 595 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 12502 595 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 531 12420 595 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 13240 514 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 13158 514 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 13076 514 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 12994 514 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 12912 514 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 12830 514 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 12748 514 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 12666 514 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 12584 514 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 12502 514 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 450 12420 514 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 13240 433 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 13158 433 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 13076 433 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 12994 433 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 12912 433 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 12830 433 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 12748 433 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 12666 433 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 12584 433 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 12502 433 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 369 12420 433 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 13240 352 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 13158 352 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 13076 352 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 12994 352 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 12912 352 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 12830 352 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 12748 352 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 12666 352 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 12584 352 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 12502 352 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 288 12420 352 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 13240 271 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 13158 271 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 13076 271 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 12994 271 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 12912 271 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 12830 271 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 12748 271 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 12666 271 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 12584 271 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 12502 271 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 207 12420 271 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 13240 190 13304 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 13158 190 13222 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 13076 190 13140 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 12994 190 13058 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 12912 190 12976 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 12830 190 12894 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 12748 190 12812 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 12666 190 12730 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 12584 190 12648 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 12502 190 12566 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 126 12420 190 12484 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10151 12418 14931 13306 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 0 12417 4895 13307 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal4 s 10156 12417 15000 13307 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal5 s 0 12437 254 13287 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal5 s 14746 12437 15000 13287 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 13252 14913 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 13170 14913 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 13088 14913 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 13006 14913 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 12924 14913 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 12842 14913 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 12760 14913 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 12678 14913 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 12596 14913 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 12514 14913 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14873 12432 14913 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 13252 14831 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 13170 14831 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 13088 14831 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 13006 14831 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 12924 14831 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 12842 14831 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 12760 14831 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 12678 14831 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 12596 14831 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 12514 14831 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14791 12432 14831 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 13252 14749 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 13170 14749 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 13088 14749 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 13006 14749 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 12924 14749 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 12842 14749 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 12760 14749 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 12678 14749 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 12596 14749 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 12514 14749 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14709 12432 14749 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 13252 14667 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 13170 14667 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 13088 14667 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 13006 14667 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 12924 14667 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 12842 14667 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 12760 14667 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 12678 14667 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 12596 14667 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 12514 14667 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14627 12432 14667 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 13252 14585 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 13170 14585 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 13088 14585 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 13006 14585 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 12924 14585 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 12842 14585 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 12760 14585 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 12678 14585 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 12596 14585 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 12514 14585 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14545 12432 14585 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 13252 14503 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 13170 14503 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 13088 14503 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 13006 14503 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 12924 14503 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 12842 14503 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 12760 14503 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 12678 14503 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 12596 14503 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 12514 14503 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14463 12432 14503 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 13252 14421 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 13170 14421 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 13088 14421 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 13006 14421 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 12924 14421 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 12842 14421 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 12760 14421 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 12678 14421 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 12596 14421 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 12514 14421 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14381 12432 14421 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 13252 14340 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 13170 14340 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 13088 14340 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 13006 14340 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 12924 14340 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 12842 14340 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 12760 14340 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 12678 14340 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 12596 14340 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 12514 14340 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14300 12432 14340 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 13252 14259 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 13170 14259 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 13088 14259 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 13006 14259 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 12924 14259 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 12842 14259 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 12760 14259 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 12678 14259 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 12596 14259 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 12514 14259 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14219 12432 14259 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 13252 14178 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 13170 14178 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 13088 14178 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 13006 14178 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 12924 14178 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 12842 14178 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 12760 14178 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 12678 14178 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 12596 14178 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 12514 14178 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14138 12432 14178 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 13252 14097 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 13170 14097 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 13088 14097 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 13006 14097 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 12924 14097 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 12842 14097 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 12760 14097 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 12678 14097 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 12596 14097 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 12514 14097 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 14057 12432 14097 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 13252 14016 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 13170 14016 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 13088 14016 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 13006 14016 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 12924 14016 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 12842 14016 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 12760 14016 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 12678 14016 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 12596 14016 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 12514 14016 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13976 12432 14016 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 13252 13935 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 13170 13935 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 13088 13935 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 13006 13935 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 12924 13935 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 12842 13935 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 12760 13935 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 12678 13935 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 12596 13935 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 12514 13935 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13895 12432 13935 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 13252 13854 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 13170 13854 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 13088 13854 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 13006 13854 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 12924 13854 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 12842 13854 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 12760 13854 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 12678 13854 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 12596 13854 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 12514 13854 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13814 12432 13854 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 13252 13773 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 13170 13773 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 13088 13773 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 13006 13773 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 12924 13773 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 12842 13773 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 12760 13773 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 12678 13773 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 12596 13773 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 12514 13773 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13733 12432 13773 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 13252 13692 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 13170 13692 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 13088 13692 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 13006 13692 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 12924 13692 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 12842 13692 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 12760 13692 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 12678 13692 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 12596 13692 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 12514 13692 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13652 12432 13692 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 13252 13611 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 13170 13611 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 13088 13611 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 13006 13611 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 12924 13611 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 12842 13611 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 12760 13611 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 12678 13611 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 12596 13611 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 12514 13611 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13571 12432 13611 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 13252 13530 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 13170 13530 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 13088 13530 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 13006 13530 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 12924 13530 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 12842 13530 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 12760 13530 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 12678 13530 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 12596 13530 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 12514 13530 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13490 12432 13530 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 13252 13449 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 13170 13449 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 13088 13449 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 13006 13449 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 12924 13449 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 12842 13449 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 12760 13449 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 12678 13449 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 12596 13449 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 12514 13449 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13409 12432 13449 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 13252 13368 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 13170 13368 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 13088 13368 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 13006 13368 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 12924 13368 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 12842 13368 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 12760 13368 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 12678 13368 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 12596 13368 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 12514 13368 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13328 12432 13368 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 13252 13287 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 13170 13287 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 13088 13287 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 13006 13287 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 12924 13287 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 12842 13287 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 12760 13287 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 12678 13287 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 12596 13287 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 12514 13287 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13247 12432 13287 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 13252 13206 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 13170 13206 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 13088 13206 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 13006 13206 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 12924 13206 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 12842 13206 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 12760 13206 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 12678 13206 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 12596 13206 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 12514 13206 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13166 12432 13206 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 13252 13125 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 13170 13125 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 13088 13125 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 13006 13125 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 12924 13125 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 12842 13125 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 12760 13125 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 12678 13125 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 12596 13125 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 12514 13125 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13085 12432 13125 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 13252 13044 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 13170 13044 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 13088 13044 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 13006 13044 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 12924 13044 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 12842 13044 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 12760 13044 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 12678 13044 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 12596 13044 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 12514 13044 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 13004 12432 13044 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 13252 12963 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 13170 12963 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 13088 12963 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 13006 12963 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 12924 12963 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 12842 12963 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 12760 12963 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 12678 12963 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 12596 12963 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 12514 12963 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12923 12432 12963 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 13252 12882 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 13170 12882 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 13088 12882 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 13006 12882 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 12924 12882 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 12842 12882 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 12760 12882 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 12678 12882 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 12596 12882 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 12514 12882 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12842 12432 12882 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 13252 12801 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 13170 12801 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 13088 12801 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 13006 12801 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 12924 12801 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 12842 12801 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 12760 12801 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 12678 12801 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 12596 12801 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 12514 12801 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12761 12432 12801 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 13252 12720 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 13170 12720 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 13088 12720 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 13006 12720 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 12924 12720 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 12842 12720 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 12760 12720 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 12678 12720 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 12596 12720 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 12514 12720 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12680 12432 12720 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 13252 12639 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 13170 12639 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 13088 12639 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 13006 12639 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 12924 12639 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 12842 12639 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 12760 12639 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 12678 12639 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 12596 12639 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 12514 12639 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12599 12432 12639 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 13252 12558 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 13170 12558 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 13088 12558 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 13006 12558 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 12924 12558 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 12842 12558 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 12760 12558 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 12678 12558 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 12596 12558 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 12514 12558 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12518 12432 12558 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 13252 12477 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 13170 12477 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 13088 12477 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 13006 12477 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 12924 12477 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 12842 12477 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 12760 12477 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 12678 12477 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 12596 12477 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 12514 12477 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12437 12432 12477 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 13252 12396 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 13170 12396 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 13088 12396 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 13006 12396 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 12924 12396 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 12842 12396 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 12760 12396 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 12678 12396 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 12596 12396 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 12514 12396 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12356 12432 12396 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 13252 12315 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 13170 12315 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 13088 12315 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 13006 12315 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 12924 12315 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 12842 12315 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 12760 12315 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 12678 12315 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 12596 12315 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 12514 12315 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12275 12432 12315 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 13252 12234 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 13170 12234 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 13088 12234 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 13006 12234 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 12924 12234 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 12842 12234 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 12760 12234 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 12678 12234 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 12596 12234 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 12514 12234 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12194 12432 12234 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 13252 12153 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 13170 12153 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 13088 12153 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 13006 12153 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 12924 12153 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 12842 12153 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 12760 12153 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 12678 12153 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 12596 12153 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 12514 12153 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12113 12432 12153 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 13252 12072 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 13170 12072 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 13088 12072 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 13006 12072 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 12924 12072 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 12842 12072 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 12760 12072 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 12678 12072 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 12596 12072 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 12514 12072 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 12032 12432 12072 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 13252 11991 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 13170 11991 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 13088 11991 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 13006 11991 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 12924 11991 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 12842 11991 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 12760 11991 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 12678 11991 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 12596 11991 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 12514 11991 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11951 12432 11991 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 13252 11910 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 13170 11910 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 13088 11910 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 13006 11910 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 12924 11910 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 12842 11910 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 12760 11910 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 12678 11910 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 12596 11910 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 12514 11910 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11870 12432 11910 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 13252 11829 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 13170 11829 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 13088 11829 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 13006 11829 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 12924 11829 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 12842 11829 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 12760 11829 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 12678 11829 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 12596 11829 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 12514 11829 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11789 12432 11829 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 13252 11748 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 13170 11748 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 13088 11748 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 13006 11748 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 12924 11748 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 12842 11748 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 12760 11748 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 12678 11748 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 12596 11748 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 12514 11748 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11708 12432 11748 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 13252 11667 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 13170 11667 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 13088 11667 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 13006 11667 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 12924 11667 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 12842 11667 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 12760 11667 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 12678 11667 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 12596 11667 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 12514 11667 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11627 12432 11667 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 13252 11586 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 13170 11586 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 13088 11586 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 13006 11586 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 12924 11586 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 12842 11586 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 12760 11586 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 12678 11586 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 12596 11586 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 12514 11586 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11546 12432 11586 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 13252 11505 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 13170 11505 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 13088 11505 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 13006 11505 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 12924 11505 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 12842 11505 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 12760 11505 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 12678 11505 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 12596 11505 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 12514 11505 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11465 12432 11505 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 13252 11424 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 13170 11424 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 13088 11424 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 13006 11424 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 12924 11424 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 12842 11424 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 12760 11424 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 12678 11424 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 12596 11424 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 12514 11424 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11384 12432 11424 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 13252 11343 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 13170 11343 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 13088 11343 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 13006 11343 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 12924 11343 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 12842 11343 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 12760 11343 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 12678 11343 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 12596 11343 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 12514 11343 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11303 12432 11343 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 13252 11262 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 13170 11262 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 13088 11262 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 13006 11262 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 12924 11262 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 12842 11262 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 12760 11262 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 12678 11262 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 12596 11262 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 12514 11262 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11222 12432 11262 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 13252 11181 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 13170 11181 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 13088 11181 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 13006 11181 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 12924 11181 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 12842 11181 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 12760 11181 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 12678 11181 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 12596 11181 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 12514 11181 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11141 12432 11181 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 13252 11100 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 13170 11100 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 13088 11100 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 13006 11100 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 12924 11100 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 12842 11100 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 12760 11100 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 12678 11100 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 12596 11100 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 12514 11100 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 11060 12432 11100 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 13252 11019 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 13170 11019 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 13088 11019 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 13006 11019 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 12924 11019 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 12842 11019 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 12760 11019 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 12678 11019 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 12596 11019 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 12514 11019 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10979 12432 11019 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 13252 10938 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 13170 10938 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 13088 10938 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 13006 10938 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 12924 10938 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 12842 10938 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 12760 10938 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 12678 10938 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 12596 10938 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 12514 10938 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10898 12432 10938 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 13252 10857 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 13170 10857 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 13088 10857 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 13006 10857 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 12924 10857 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 12842 10857 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 12760 10857 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 12678 10857 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 12596 10857 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 12514 10857 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10817 12432 10857 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 13252 10776 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 13170 10776 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 13088 10776 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 13006 10776 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 12924 10776 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 12842 10776 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 12760 10776 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 12678 10776 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 12596 10776 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 12514 10776 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10736 12432 10776 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 13252 10695 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 13170 10695 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 13088 10695 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 13006 10695 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 12924 10695 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 12842 10695 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 12760 10695 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 12678 10695 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 12596 10695 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 12514 10695 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10655 12432 10695 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 13252 10614 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 13170 10614 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 13088 10614 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 13006 10614 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 12924 10614 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 12842 10614 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 12760 10614 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 12678 10614 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 12596 10614 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 12514 10614 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10574 12432 10614 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 13252 10533 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 13170 10533 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 13088 10533 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 13006 10533 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 12924 10533 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 12842 10533 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 12760 10533 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 12678 10533 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 12596 10533 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 12514 10533 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10493 12432 10533 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 13252 10452 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 13170 10452 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 13088 10452 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 13006 10452 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 12924 10452 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 12842 10452 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 12760 10452 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 12678 10452 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 12596 10452 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 12514 10452 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10412 12432 10452 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 13252 10371 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 13170 10371 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 13088 10371 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 13006 10371 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 12924 10371 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 12842 10371 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 12760 10371 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 12678 10371 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 12596 10371 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 12514 10371 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10331 12432 10371 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 13252 10290 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 13170 10290 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 13088 10290 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 13006 10290 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 12924 10290 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 12842 10290 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 12760 10290 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 12678 10290 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 12596 10290 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 12514 10290 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10250 12432 10290 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 13252 10209 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 13170 10209 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 13088 10209 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 13006 10209 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 12924 10209 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 12842 10209 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 12760 10209 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 12678 10209 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 12596 10209 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 12514 10209 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 10169 12432 10209 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4842 13252 4882 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4842 13170 4882 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4842 13088 4882 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4842 13006 4882 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4842 12924 4882 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4842 12842 4882 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4842 12760 4882 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4842 12678 4882 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4842 12596 4882 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4842 12514 4882 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4842 12432 4882 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4760 13252 4800 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4760 13170 4800 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4760 13088 4800 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4760 13006 4800 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4760 12924 4800 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4760 12842 4800 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4760 12760 4800 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4760 12678 4800 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4760 12596 4800 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4760 12514 4800 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4760 12432 4800 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4678 13252 4718 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4678 13170 4718 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4678 13088 4718 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4678 13006 4718 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4678 12924 4718 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4678 12842 4718 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4678 12760 4718 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4678 12678 4718 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4678 12596 4718 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4678 12514 4718 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4678 12432 4718 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4596 13252 4636 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4596 13170 4636 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4596 13088 4636 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4596 13006 4636 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4596 12924 4636 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4596 12842 4636 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4596 12760 4636 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4596 12678 4636 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4596 12596 4636 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4596 12514 4636 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4596 12432 4636 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4514 13252 4554 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4514 13170 4554 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4514 13088 4554 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4514 13006 4554 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4514 12924 4554 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4514 12842 4554 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4514 12760 4554 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4514 12678 4554 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4514 12596 4554 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4514 12514 4554 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4514 12432 4554 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4432 13252 4472 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4432 13170 4472 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4432 13088 4472 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4432 13006 4472 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4432 12924 4472 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4432 12842 4472 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4432 12760 4472 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4432 12678 4472 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4432 12596 4472 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4432 12514 4472 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4432 12432 4472 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4350 13252 4390 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4350 13170 4390 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4350 13088 4390 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4350 13006 4390 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4350 12924 4390 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4350 12842 4390 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4350 12760 4390 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4350 12678 4390 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4350 12596 4390 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4350 12514 4390 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4350 12432 4390 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4269 13252 4309 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4269 13170 4309 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4269 13088 4309 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4269 13006 4309 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4269 12924 4309 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4269 12842 4309 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4269 12760 4309 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4269 12678 4309 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4269 12596 4309 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4269 12514 4309 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4269 12432 4309 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4188 13252 4228 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4188 13170 4228 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4188 13088 4228 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4188 13006 4228 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4188 12924 4228 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4188 12842 4228 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4188 12760 4228 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4188 12678 4228 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4188 12596 4228 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4188 12514 4228 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4188 12432 4228 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4107 13252 4147 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4107 13170 4147 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4107 13088 4147 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4107 13006 4147 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4107 12924 4147 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4107 12842 4147 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4107 12760 4147 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4107 12678 4147 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4107 12596 4147 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4107 12514 4147 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4107 12432 4147 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4026 13252 4066 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4026 13170 4066 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4026 13088 4066 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4026 13006 4066 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4026 12924 4066 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4026 12842 4066 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4026 12760 4066 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4026 12678 4066 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4026 12596 4066 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4026 12514 4066 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 4026 12432 4066 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3945 13252 3985 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3945 13170 3985 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3945 13088 3985 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3945 13006 3985 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3945 12924 3985 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3945 12842 3985 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3945 12760 3985 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3945 12678 3985 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3945 12596 3985 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3945 12514 3985 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3945 12432 3985 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3864 13252 3904 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3864 13170 3904 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3864 13088 3904 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3864 13006 3904 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3864 12924 3904 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3864 12842 3904 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3864 12760 3904 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3864 12678 3904 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3864 12596 3904 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3864 12514 3904 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3864 12432 3904 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3783 13252 3823 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3783 13170 3823 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3783 13088 3823 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3783 13006 3823 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3783 12924 3823 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3783 12842 3823 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3783 12760 3823 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3783 12678 3823 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3783 12596 3823 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3783 12514 3823 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3783 12432 3823 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3702 13252 3742 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3702 13170 3742 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3702 13088 3742 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3702 13006 3742 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3702 12924 3742 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3702 12842 3742 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3702 12760 3742 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3702 12678 3742 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3702 12596 3742 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3702 12514 3742 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3702 12432 3742 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3621 13252 3661 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3621 13170 3661 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3621 13088 3661 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3621 13006 3661 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3621 12924 3661 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3621 12842 3661 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3621 12760 3661 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3621 12678 3661 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3621 12596 3661 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3621 12514 3661 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3621 12432 3661 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3540 13252 3580 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3540 13170 3580 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3540 13088 3580 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3540 13006 3580 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3540 12924 3580 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3540 12842 3580 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3540 12760 3580 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3540 12678 3580 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3540 12596 3580 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3540 12514 3580 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3540 12432 3580 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3459 13252 3499 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3459 13170 3499 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3459 13088 3499 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3459 13006 3499 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3459 12924 3499 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3459 12842 3499 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3459 12760 3499 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3459 12678 3499 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3459 12596 3499 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3459 12514 3499 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3459 12432 3499 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3378 13252 3418 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3378 13170 3418 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3378 13088 3418 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3378 13006 3418 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3378 12924 3418 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3378 12842 3418 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3378 12760 3418 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3378 12678 3418 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3378 12596 3418 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3378 12514 3418 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3378 12432 3418 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3297 13252 3337 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3297 13170 3337 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3297 13088 3337 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3297 13006 3337 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3297 12924 3337 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3297 12842 3337 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3297 12760 3337 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3297 12678 3337 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3297 12596 3337 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3297 12514 3337 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3297 12432 3337 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3216 13252 3256 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3216 13170 3256 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3216 13088 3256 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3216 13006 3256 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3216 12924 3256 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3216 12842 3256 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3216 12760 3256 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3216 12678 3256 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3216 12596 3256 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3216 12514 3256 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3216 12432 3256 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3135 13252 3175 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3135 13170 3175 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3135 13088 3175 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3135 13006 3175 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3135 12924 3175 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3135 12842 3175 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3135 12760 3175 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3135 12678 3175 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3135 12596 3175 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3135 12514 3175 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3135 12432 3175 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3054 13252 3094 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3054 13170 3094 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3054 13088 3094 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3054 13006 3094 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3054 12924 3094 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3054 12842 3094 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3054 12760 3094 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3054 12678 3094 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3054 12596 3094 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3054 12514 3094 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 3054 12432 3094 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2973 13252 3013 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2973 13170 3013 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2973 13088 3013 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2973 13006 3013 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2973 12924 3013 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2973 12842 3013 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2973 12760 3013 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2973 12678 3013 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2973 12596 3013 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2973 12514 3013 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2973 12432 3013 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2892 13252 2932 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2892 13170 2932 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2892 13088 2932 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2892 13006 2932 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2892 12924 2932 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2892 12842 2932 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2892 12760 2932 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2892 12678 2932 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2892 12596 2932 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2892 12514 2932 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2892 12432 2932 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2811 13252 2851 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2811 13170 2851 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2811 13088 2851 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2811 13006 2851 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2811 12924 2851 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2811 12842 2851 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2811 12760 2851 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2811 12678 2851 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2811 12596 2851 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2811 12514 2851 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2811 12432 2851 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2730 13252 2770 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2730 13170 2770 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2730 13088 2770 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2730 13006 2770 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2730 12924 2770 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2730 12842 2770 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2730 12760 2770 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2730 12678 2770 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2730 12596 2770 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2730 12514 2770 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2730 12432 2770 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2649 13252 2689 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2649 13170 2689 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2649 13088 2689 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2649 13006 2689 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2649 12924 2689 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2649 12842 2689 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2649 12760 2689 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2649 12678 2689 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2649 12596 2689 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2649 12514 2689 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2649 12432 2689 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2568 13252 2608 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2568 13170 2608 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2568 13088 2608 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2568 13006 2608 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2568 12924 2608 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2568 12842 2608 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2568 12760 2608 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2568 12678 2608 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2568 12596 2608 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2568 12514 2608 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2568 12432 2608 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2487 13252 2527 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2487 13170 2527 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2487 13088 2527 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2487 13006 2527 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2487 12924 2527 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2487 12842 2527 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2487 12760 2527 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2487 12678 2527 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2487 12596 2527 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2487 12514 2527 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2487 12432 2527 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2406 13252 2446 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2406 13170 2446 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2406 13088 2446 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2406 13006 2446 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2406 12924 2446 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2406 12842 2446 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2406 12760 2446 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2406 12678 2446 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2406 12596 2446 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2406 12514 2446 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2406 12432 2446 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2325 13252 2365 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2325 13170 2365 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2325 13088 2365 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2325 13006 2365 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2325 12924 2365 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2325 12842 2365 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2325 12760 2365 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2325 12678 2365 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2325 12596 2365 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2325 12514 2365 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2325 12432 2365 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2244 13252 2284 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2244 13170 2284 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2244 13088 2284 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2244 13006 2284 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2244 12924 2284 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2244 12842 2284 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2244 12760 2284 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2244 12678 2284 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2244 12596 2284 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2244 12514 2284 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2244 12432 2284 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2163 13252 2203 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2163 13170 2203 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2163 13088 2203 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2163 13006 2203 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2163 12924 2203 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2163 12842 2203 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2163 12760 2203 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2163 12678 2203 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2163 12596 2203 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2163 12514 2203 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2163 12432 2203 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2082 13252 2122 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2082 13170 2122 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2082 13088 2122 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2082 13006 2122 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2082 12924 2122 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2082 12842 2122 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2082 12760 2122 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2082 12678 2122 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2082 12596 2122 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2082 12514 2122 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2082 12432 2122 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2001 13252 2041 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2001 13170 2041 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2001 13088 2041 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2001 13006 2041 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2001 12924 2041 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2001 12842 2041 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2001 12760 2041 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2001 12678 2041 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2001 12596 2041 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2001 12514 2041 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 2001 12432 2041 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1920 13252 1960 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1920 13170 1960 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1920 13088 1960 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1920 13006 1960 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1920 12924 1960 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1920 12842 1960 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1920 12760 1960 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1920 12678 1960 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1920 12596 1960 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1920 12514 1960 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1920 12432 1960 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1839 13252 1879 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1839 13170 1879 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1839 13088 1879 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1839 13006 1879 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1839 12924 1879 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1839 12842 1879 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1839 12760 1879 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1839 12678 1879 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1839 12596 1879 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1839 12514 1879 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1839 12432 1879 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1758 13252 1798 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1758 13170 1798 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1758 13088 1798 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1758 13006 1798 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1758 12924 1798 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1758 12842 1798 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1758 12760 1798 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1758 12678 1798 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1758 12596 1798 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1758 12514 1798 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1758 12432 1798 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1677 13252 1717 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1677 13170 1717 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1677 13088 1717 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1677 13006 1717 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1677 12924 1717 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1677 12842 1717 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1677 12760 1717 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1677 12678 1717 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1677 12596 1717 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1677 12514 1717 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1677 12432 1717 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1596 13252 1636 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1596 13170 1636 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1596 13088 1636 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1596 13006 1636 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1596 12924 1636 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1596 12842 1636 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1596 12760 1636 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1596 12678 1636 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1596 12596 1636 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1596 12514 1636 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1596 12432 1636 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1515 13252 1555 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1515 13170 1555 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1515 13088 1555 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1515 13006 1555 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1515 12924 1555 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1515 12842 1555 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1515 12760 1555 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1515 12678 1555 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1515 12596 1555 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1515 12514 1555 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1515 12432 1555 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1434 13252 1474 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1434 13170 1474 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1434 13088 1474 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1434 13006 1474 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1434 12924 1474 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1434 12842 1474 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1434 12760 1474 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1434 12678 1474 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1434 12596 1474 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1434 12514 1474 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1434 12432 1474 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1353 13252 1393 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1353 13170 1393 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1353 13088 1393 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1353 13006 1393 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1353 12924 1393 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1353 12842 1393 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1353 12760 1393 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1353 12678 1393 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1353 12596 1393 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1353 12514 1393 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1353 12432 1393 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1272 13252 1312 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1272 13170 1312 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1272 13088 1312 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1272 13006 1312 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1272 12924 1312 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1272 12842 1312 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1272 12760 1312 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1272 12678 1312 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1272 12596 1312 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1272 12514 1312 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1272 12432 1312 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1191 13252 1231 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1191 13170 1231 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1191 13088 1231 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1191 13006 1231 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1191 12924 1231 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1191 12842 1231 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1191 12760 1231 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1191 12678 1231 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1191 12596 1231 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1191 12514 1231 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1191 12432 1231 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1110 13252 1150 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1110 13170 1150 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1110 13088 1150 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1110 13006 1150 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1110 12924 1150 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1110 12842 1150 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1110 12760 1150 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1110 12678 1150 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1110 12596 1150 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1110 12514 1150 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1110 12432 1150 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1029 13252 1069 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1029 13170 1069 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1029 13088 1069 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1029 13006 1069 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1029 12924 1069 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1029 12842 1069 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1029 12760 1069 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1029 12678 1069 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1029 12596 1069 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1029 12514 1069 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 1029 12432 1069 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 948 13252 988 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 948 13170 988 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 948 13088 988 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 948 13006 988 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 948 12924 988 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 948 12842 988 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 948 12760 988 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 948 12678 988 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 948 12596 988 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 948 12514 988 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 948 12432 988 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 867 13252 907 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 867 13170 907 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 867 13088 907 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 867 13006 907 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 867 12924 907 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 867 12842 907 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 867 12760 907 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 867 12678 907 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 867 12596 907 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 867 12514 907 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 867 12432 907 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 786 13252 826 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 786 13170 826 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 786 13088 826 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 786 13006 826 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 786 12924 826 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 786 12842 826 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 786 12760 826 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 786 12678 826 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 786 12596 826 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 786 12514 826 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 786 12432 826 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 705 13252 745 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 705 13170 745 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 705 13088 745 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 705 13006 745 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 705 12924 745 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 705 12842 745 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 705 12760 745 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 705 12678 745 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 705 12596 745 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 705 12514 745 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 705 12432 745 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 624 13252 664 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 624 13170 664 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 624 13088 664 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 624 13006 664 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 624 12924 664 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 624 12842 664 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 624 12760 664 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 624 12678 664 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 624 12596 664 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 624 12514 664 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 624 12432 664 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 543 13252 583 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 543 13170 583 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 543 13088 583 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 543 13006 583 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 543 12924 583 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 543 12842 583 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 543 12760 583 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 543 12678 583 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 543 12596 583 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 543 12514 583 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 543 12432 583 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 462 13252 502 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 462 13170 502 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 462 13088 502 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 462 13006 502 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 462 12924 502 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 462 12842 502 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 462 12760 502 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 462 12678 502 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 462 12596 502 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 462 12514 502 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 462 12432 502 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 381 13252 421 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 381 13170 421 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 381 13088 421 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 381 13006 421 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 381 12924 421 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 381 12842 421 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 381 12760 421 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 381 12678 421 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 381 12596 421 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 381 12514 421 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 381 12432 421 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 300 13252 340 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 300 13170 340 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 300 13088 340 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 300 13006 340 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 300 12924 340 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 300 12842 340 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 300 12760 340 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 300 12678 340 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 300 12596 340 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 300 12514 340 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 300 12432 340 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 219 13252 259 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 219 13170 259 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 219 13088 259 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 219 13006 259 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 219 12924 259 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 219 12842 259 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 219 12760 259 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 219 12678 259 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 219 12596 259 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 219 12514 259 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 219 12432 259 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 138 13252 178 13292 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 138 13170 178 13210 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 138 13088 178 13128 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 138 13006 178 13046 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 138 12924 178 12964 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 138 12842 178 12882 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 138 12760 178 12800 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 138 12678 178 12718 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 138 12596 178 12636 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 138 12514 178 12554 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal3 s 138 12432 178 12472 6 VDDIO_Q
port 1 nsew power bidirectional
rlabel metal5 s 14807 2607 15000 3257 6 VDDA
port 2 nsew power bidirectional
rlabel metal5 s 0 2607 193 3257 6 VDDA
port 2 nsew power bidirectional
rlabel metal4 s 0 2587 193 3277 6 VDDA
port 2 nsew power bidirectional
rlabel metal4 s 14807 2587 15000 3277 6 VDDA
port 2 nsew power bidirectional
rlabel metal4 s 14807 2587 15000 3277 6 VDDA
port 2 nsew power bidirectional
rlabel metal5 s 0 2607 193 3257 6 VDDA
port 2 nsew power bidirectional
rlabel metal5 s 14807 2607 15000 3257 6 VDDA
port 2 nsew power bidirectional
rlabel metal4 s 14807 2587 15000 3277 6 VDDA
port 2 nsew power bidirectional
rlabel metal5 s 0 2607 193 3257 6 VDDA
port 2 nsew power bidirectional
rlabel metal5 s 14807 2607 15000 3257 6 VDDA
port 2 nsew power bidirectional
rlabel metal5 s 14746 9147 15000 10947 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 14746 6968 15000 7617 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 9147 254 10947 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 6968 254 7617 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 6947 15000 7637 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 9147 15000 9213 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 10881 15000 10947 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 9929 15000 10165 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 9147 254 9213 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 9929 254 10165 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 10881 254 10947 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 6947 254 7637 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 9147 254 9213 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 9929 254 10165 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 10881 254 10947 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 6947 15000 7637 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 9147 15000 9213 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 9929 15000 10165 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 10881 15000 10947 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 6968 254 7617 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 9147 254 10947 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 14746 6968 15000 7617 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 14746 9147 15000 10947 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 9147 254 9213 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 9929 254 10165 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 0 10881 254 10947 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 6947 15000 7637 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 9147 15000 9213 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 9929 15000 10165 6 VSSA
port 3 nsew ground bidirectional
rlabel metal4 s 14746 10881 15000 10947 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 6968 254 7617 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 9147 254 10947 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 14746 6968 15000 7617 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 14746 9147 15000 10947 6 VSSA
port 3 nsew ground bidirectional
rlabel metal5 s 0 1397 254 2287 6 VCCD
port 4 nsew power bidirectional
rlabel metal5 s 14746 1397 15000 2287 6 VCCD
port 4 nsew power bidirectional
rlabel metal4 s 14746 1377 15000 2307 6 VCCD
port 4 nsew power bidirectional
rlabel metal4 s 0 1377 254 2307 6 VCCD
port 4 nsew power bidirectional
rlabel metal4 s 14746 1377 15000 2307 6 VCCD
port 4 nsew power bidirectional
rlabel metal5 s 0 1397 254 2287 6 VCCD
port 4 nsew power bidirectional
rlabel metal5 s 14746 1397 15000 2287 6 VCCD
port 4 nsew power bidirectional
rlabel metal4 s 14746 1377 15000 2307 6 VCCD
port 4 nsew power bidirectional
rlabel metal5 s 0 1397 254 2287 6 VCCD
port 4 nsew power bidirectional
rlabel metal5 s 14746 1397 15000 2287 6 VCCD
port 4 nsew power bidirectional
rlabel metal5 s 0 27 254 1077 6 VCCHIB
port 5 nsew power bidirectional
rlabel metal5 s 14746 27 15000 1077 6 VCCHIB
port 5 nsew power bidirectional
rlabel metal4 s 14746 7 15000 1097 6 VCCHIB
port 5 nsew power bidirectional
rlabel metal4 s 0 7 254 1097 6 VCCHIB
port 5 nsew power bidirectional
rlabel metal4 s 14746 7 15000 1097 6 VCCHIB
port 5 nsew power bidirectional
rlabel metal5 s 0 27 254 1077 6 VCCHIB
port 5 nsew power bidirectional
rlabel metal5 s 14746 27 15000 1077 6 VCCHIB
port 5 nsew power bidirectional
rlabel metal4 s 14746 7 15000 1097 6 VCCHIB
port 5 nsew power bidirectional
rlabel metal5 s 0 27 254 1077 6 VCCHIB
port 5 nsew power bidirectional
rlabel metal5 s 14746 27 15000 1077 6 VCCHIB
port 5 nsew power bidirectional
rlabel metal5 s 14746 7937 15000 8827 6 VSSD
port 6 nsew ground bidirectional
rlabel metal5 s 0 7937 254 8827 6 VSSD
port 6 nsew ground bidirectional
rlabel metal4 s 14746 7917 15000 8847 6 VSSD
port 6 nsew ground bidirectional
rlabel metal4 s 0 7917 254 8847 6 VSSD
port 6 nsew ground bidirectional
rlabel metal4 s 14746 7917 15000 8847 6 VSSD
port 6 nsew ground bidirectional
rlabel metal5 s 0 7937 254 8827 6 VSSD
port 6 nsew ground bidirectional
rlabel metal5 s 14746 7937 15000 8827 6 VSSD
port 6 nsew ground bidirectional
rlabel metal4 s 14746 7917 15000 8847 6 VSSD
port 6 nsew ground bidirectional
rlabel metal5 s 0 7937 254 8827 6 VSSD
port 6 nsew ground bidirectional
rlabel metal5 s 14746 7937 15000 8827 6 VSSD
port 6 nsew ground bidirectional
rlabel metal5 s 14746 13607 15000 18597 6 VDDIO
port 7 nsew power bidirectional
rlabel metal5 s 14746 3577 15000 4467 6 VDDIO
port 7 nsew power bidirectional
rlabel metal5 s 0 13607 254 18597 6 VDDIO
port 7 nsew power bidirectional
rlabel metal5 s 0 3577 254 4467 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14746 3557 15000 4487 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14746 13607 15000 18600 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 0 3557 254 4487 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 0 13607 254 18600 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 120 3558 4900 4486 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10151 3558 14931 4486 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12211 18573 14932 18592 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11966 18347 12211 18592 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12162 18513 14932 18543 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12132 18483 14932 18513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12102 18453 14932 18483 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12072 18423 14932 18453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 18393 14932 18423 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12012 18363 14932 18393 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11982 18333 14932 18363 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11788 18169 11966 18347 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11922 18273 14932 18303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11892 18243 14932 18273 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11862 18213 14932 18243 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11832 18183 14932 18213 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 18153 14932 18183 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11530 17911 11788 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11742 18093 14932 18123 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11712 18063 14932 18093 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11682 18033 14932 18063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11652 18003 14932 18033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11622 17973 14932 18003 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11592 17943 14932 17973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 17913 14932 17943 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11532 17883 14932 17913 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11283 17664 11530 17911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11472 17823 14932 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11442 17793 14932 17823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11412 17763 14932 17793 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11382 17733 14932 17763 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11352 17703 14932 17733 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 17673 14932 17703 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11292 17643 14932 17673 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11027 17408 11283 17664 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11232 17583 14932 17613 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11202 17553 14932 17583 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11172 17523 14932 17553 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11142 17493 14932 17523 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11112 17463 14932 17493 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 17433 14932 17463 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11052 17403 14932 17433 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10742 17123 11027 17408 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10992 17343 14932 17373 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10962 17313 14932 17343 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10932 17283 14932 17313 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10902 17253 14932 17283 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10872 17223 14932 17253 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 17193 14932 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10812 17163 14932 17193 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10782 17133 14932 17163 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10752 17103 14932 17133 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10481 16862 10742 17123 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10692 17043 14932 17073 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10662 17013 14932 17043 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10632 16983 14932 17013 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 16953 14932 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10572 16923 14932 16953 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10542 16893 14932 16923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10512 16863 14932 16893 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10482 16833 14932 16863 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10152 16533 10481 16862 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10422 16773 14932 16803 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10392 16743 14932 16773 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 16713 14932 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10332 16683 14932 16713 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10302 16653 14932 16683 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10272 16623 14932 16653 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10242 16593 14932 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10212 16563 14932 16593 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10182 16533 14932 16563 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10152 13607 14932 16533 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 0 3557 4895 4487 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 0 18592 254 18600 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 0 16558 2821 18592 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 0 16525 254 16558 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 0 13612 4900 16525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 0 13607 254 13612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2851 18190 3073 18342 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2854 17669 3250 18164 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2875 16598 3771 17628 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3283 17673 3505 17906 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3799 17162 4013 17403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3834 16589 4290 17118 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4330 16571 4554 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14746 18593 15000 18600 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14746 16525 15000 16557 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14746 13607 15000 13612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12230 16557 15000 18593 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10151 13612 15000 16525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10156 3557 15000 4487 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10497 16571 10721 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10761 16589 11217 17118 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11038 17162 11252 17403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11280 16598 12176 17628 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11546 17673 11768 17906 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11801 17669 12197 18164 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11978 18190 12200 18342 6 VDDIO
port 7 nsew power bidirectional
rlabel metal5 s 0 3577 254 4467 6 VDDIO
port 7 nsew power bidirectional
rlabel metal5 s 0 13607 254 18597 6 VDDIO
port 7 nsew power bidirectional
rlabel metal5 s 14746 3577 15000 4467 6 VDDIO
port 7 nsew power bidirectional
rlabel metal5 s 14746 13607 15000 18597 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 4432 14913 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 4346 14913 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 4260 14913 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 4174 14913 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 4088 14913 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 4002 14913 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 3916 14913 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 3830 14913 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 3744 14913 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 3658 14913 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 3572 14913 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 18539 14904 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 18457 14904 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 18375 14904 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 18293 14904 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 18211 14904 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 18129 14904 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 18047 14904 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 17965 14904 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 17883 14904 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 17801 14904 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 17719 14904 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 17637 14904 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 17555 14904 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 17473 14904 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 17391 14904 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 17309 14904 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 17227 14904 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 17145 14904 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 17063 14904 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 16981 14904 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 16899 14904 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 16817 14904 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 16735 14904 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 16653 14904 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 16571 14904 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 16472 14882 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 16391 14882 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 16310 14882 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 16229 14882 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 16148 14882 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 16067 14882 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15986 14882 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15905 14882 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15824 14882 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15743 14882 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15662 14882 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15581 14882 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15500 14882 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15419 14882 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15338 14882 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15257 14882 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15176 14882 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15095 14882 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15014 14882 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14933 14882 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14852 14882 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14771 14882 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14690 14882 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14609 14882 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14527 14882 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14445 14882 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14363 14882 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14281 14882 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14199 14882 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14117 14882 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14035 14882 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 13953 14882 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 13871 14882 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 13789 14882 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 13707 14882 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 13625 14882 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 4432 14831 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 4346 14831 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 4260 14831 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 4174 14831 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 4088 14831 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 4002 14831 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 3916 14831 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 3830 14831 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 3744 14831 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 3658 14831 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 3572 14831 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 18539 14822 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 18457 14822 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 18375 14822 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 18293 14822 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 18211 14822 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 18129 14822 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 18047 14822 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 17965 14822 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 17883 14822 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 17801 14822 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 17719 14822 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 17637 14822 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 17555 14822 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 17473 14822 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 17391 14822 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 17309 14822 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 17227 14822 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 17145 14822 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 17063 14822 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 16981 14822 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 16899 14822 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 16817 14822 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 16735 14822 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 16653 14822 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 16571 14822 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 16472 14802 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 16391 14802 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 16310 14802 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 16229 14802 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 16148 14802 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 16067 14802 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15986 14802 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15905 14802 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15824 14802 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15743 14802 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15662 14802 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15581 14802 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15500 14802 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15419 14802 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15338 14802 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15257 14802 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15176 14802 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15095 14802 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15014 14802 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14933 14802 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14852 14802 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14771 14802 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14690 14802 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14609 14802 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14527 14802 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14445 14802 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14363 14802 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14281 14802 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14199 14802 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14117 14802 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14035 14802 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 13953 14802 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 13871 14802 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 13789 14802 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 13707 14802 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 13625 14802 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 4432 14749 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 4346 14749 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 4260 14749 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 4174 14749 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 4088 14749 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 4002 14749 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 3916 14749 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 3830 14749 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 3744 14749 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 3658 14749 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 3572 14749 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 18539 14740 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 18457 14740 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 18375 14740 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 18293 14740 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 18211 14740 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 18129 14740 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 18047 14740 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 17965 14740 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 17883 14740 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 17801 14740 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 17719 14740 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 17637 14740 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 17555 14740 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 17473 14740 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 17391 14740 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 17309 14740 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 17227 14740 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 17145 14740 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 17063 14740 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 16981 14740 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 16899 14740 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 16817 14740 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 16735 14740 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 16653 14740 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 16571 14740 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 16472 14722 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 16391 14722 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 16310 14722 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 16229 14722 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 16148 14722 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 16067 14722 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15986 14722 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15905 14722 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15824 14722 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15743 14722 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15662 14722 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15581 14722 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15500 14722 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15419 14722 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15338 14722 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15257 14722 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15176 14722 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15095 14722 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15014 14722 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14933 14722 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14852 14722 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14771 14722 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14690 14722 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14609 14722 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14527 14722 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14445 14722 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14363 14722 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14281 14722 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14199 14722 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14117 14722 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14035 14722 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 13953 14722 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 13871 14722 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 13789 14722 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 13707 14722 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 13625 14722 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 4432 14667 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 4346 14667 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 4260 14667 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 4174 14667 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 4088 14667 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 4002 14667 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 3916 14667 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 3830 14667 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 3744 14667 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 3658 14667 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 3572 14667 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 18539 14658 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 18457 14658 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 18375 14658 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 18293 14658 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 18211 14658 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 18129 14658 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 18047 14658 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 17965 14658 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 17883 14658 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 17801 14658 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 17719 14658 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 17637 14658 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 17555 14658 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 17473 14658 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 17391 14658 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 17309 14658 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 17227 14658 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 17145 14658 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 17063 14658 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 16981 14658 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 16899 14658 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 16817 14658 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 16735 14658 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 16653 14658 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 16571 14658 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 16472 14642 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 16391 14642 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 16310 14642 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 16229 14642 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 16148 14642 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 16067 14642 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15986 14642 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15905 14642 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15824 14642 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15743 14642 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15662 14642 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15581 14642 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15500 14642 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15419 14642 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15338 14642 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15257 14642 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15176 14642 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15095 14642 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15014 14642 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14933 14642 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14852 14642 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14771 14642 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14690 14642 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14609 14642 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14527 14642 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14445 14642 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14363 14642 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14281 14642 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14199 14642 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14117 14642 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14035 14642 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 13953 14642 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 13871 14642 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 13789 14642 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 13707 14642 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 13625 14642 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 4432 14585 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 4346 14585 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 4260 14585 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 4174 14585 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 4088 14585 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 4002 14585 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 3916 14585 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 3830 14585 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 3744 14585 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 3658 14585 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 3572 14585 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 18539 14576 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 18457 14576 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 18375 14576 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 18293 14576 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 18211 14576 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 18129 14576 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 18047 14576 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 17965 14576 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 17883 14576 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 17801 14576 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 17719 14576 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 17637 14576 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 17555 14576 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 17473 14576 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 17391 14576 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 17309 14576 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 17227 14576 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 17145 14576 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 17063 14576 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 16981 14576 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 16899 14576 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 16817 14576 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 16735 14576 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 16653 14576 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 16571 14576 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 16472 14562 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 16391 14562 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 16310 14562 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 16229 14562 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 16148 14562 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 16067 14562 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15986 14562 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15905 14562 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15824 14562 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15743 14562 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15662 14562 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15581 14562 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15500 14562 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15419 14562 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15338 14562 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15257 14562 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15176 14562 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15095 14562 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15014 14562 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14933 14562 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14852 14562 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14771 14562 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14690 14562 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14609 14562 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14527 14562 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14445 14562 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14363 14562 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14281 14562 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14199 14562 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14117 14562 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14035 14562 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 13953 14562 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 13871 14562 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 13789 14562 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 13707 14562 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 13625 14562 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 4432 14503 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 4346 14503 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 4260 14503 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 4174 14503 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 4088 14503 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 4002 14503 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 3916 14503 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 3830 14503 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 3744 14503 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 3658 14503 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 3572 14503 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 18539 14494 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 18457 14494 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 18375 14494 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 18293 14494 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 18211 14494 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 18129 14494 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 18047 14494 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 17965 14494 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 17883 14494 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 17801 14494 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 17719 14494 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 17637 14494 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 17555 14494 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 17473 14494 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 17391 14494 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 17309 14494 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 17227 14494 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 17145 14494 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 17063 14494 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 16981 14494 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 16899 14494 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 16817 14494 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 16735 14494 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 16653 14494 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 16571 14494 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16472 14482 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16391 14482 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16310 14482 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16229 14482 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16148 14482 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16067 14482 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15986 14482 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15905 14482 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15824 14482 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15743 14482 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15662 14482 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15581 14482 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15500 14482 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15419 14482 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15338 14482 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15257 14482 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15176 14482 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15095 14482 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15014 14482 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14933 14482 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14852 14482 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14771 14482 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14690 14482 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14609 14482 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14527 14482 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14445 14482 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14363 14482 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14281 14482 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14199 14482 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14117 14482 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14035 14482 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 13953 14482 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 13871 14482 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 13789 14482 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 13707 14482 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 13625 14482 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 4432 14421 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 4346 14421 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 4260 14421 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 4174 14421 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 4088 14421 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 4002 14421 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 3916 14421 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 3830 14421 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 3744 14421 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 3658 14421 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 3572 14421 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 18539 14412 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 18457 14412 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 18375 14412 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 18293 14412 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 18211 14412 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 18129 14412 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 18047 14412 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 17965 14412 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 17883 14412 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 17801 14412 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 17719 14412 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 17637 14412 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 17555 14412 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 17473 14412 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 17391 14412 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 17309 14412 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 17227 14412 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 17145 14412 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 17063 14412 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 16981 14412 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 16899 14412 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 16817 14412 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 16735 14412 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 16653 14412 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 16571 14412 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 16472 14402 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 16391 14402 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 16310 14402 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 16229 14402 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 16148 14402 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 16067 14402 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15986 14402 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15905 14402 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15824 14402 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15743 14402 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15662 14402 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15581 14402 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15500 14402 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15419 14402 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15338 14402 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15257 14402 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15176 14402 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15095 14402 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15014 14402 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14933 14402 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14852 14402 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14771 14402 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14690 14402 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14609 14402 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14527 14402 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14445 14402 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14363 14402 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14281 14402 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14199 14402 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14117 14402 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14035 14402 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 13953 14402 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 13871 14402 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 13789 14402 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 13707 14402 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 13625 14402 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 4432 14340 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 4346 14340 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 4260 14340 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 4174 14340 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 4088 14340 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 4002 14340 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 3916 14340 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 3830 14340 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 3744 14340 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 3658 14340 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 3572 14340 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 18539 14330 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 18457 14330 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 18375 14330 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 18293 14330 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 18211 14330 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 18129 14330 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 18047 14330 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 17965 14330 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 17883 14330 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 17801 14330 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 17719 14330 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 17637 14330 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 17555 14330 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 17473 14330 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 17391 14330 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 17309 14330 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 17227 14330 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 17145 14330 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 17063 14330 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 16981 14330 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 16899 14330 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 16817 14330 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 16735 14330 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 16653 14330 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 16571 14330 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 16472 14322 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 16391 14322 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 16310 14322 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 16229 14322 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 16148 14322 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 16067 14322 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15986 14322 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15905 14322 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15824 14322 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15743 14322 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15662 14322 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15581 14322 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15500 14322 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15419 14322 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15338 14322 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15257 14322 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15176 14322 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15095 14322 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15014 14322 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14933 14322 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14852 14322 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14771 14322 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14690 14322 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14609 14322 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14527 14322 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14445 14322 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14363 14322 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14281 14322 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14199 14322 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14117 14322 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14035 14322 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 13953 14322 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 13871 14322 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 13789 14322 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 13707 14322 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 13625 14322 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 4432 14259 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 4346 14259 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 4260 14259 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 4174 14259 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 4088 14259 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 4002 14259 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 3916 14259 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 3830 14259 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 3744 14259 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 3658 14259 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 3572 14259 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 18539 14248 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 18457 14248 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 18375 14248 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 18293 14248 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 18211 14248 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 18129 14248 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 18047 14248 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 17965 14248 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 17883 14248 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 17801 14248 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 17719 14248 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 17637 14248 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 17555 14248 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 17473 14248 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 17391 14248 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 17309 14248 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 17227 14248 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 17145 14248 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 17063 14248 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 16981 14248 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 16899 14248 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 16817 14248 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 16735 14248 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 16653 14248 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 16571 14248 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 16472 14242 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 16391 14242 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 16310 14242 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 16229 14242 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 16148 14242 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 16067 14242 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15986 14242 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15905 14242 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15824 14242 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15743 14242 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15662 14242 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15581 14242 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15500 14242 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15419 14242 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15338 14242 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15257 14242 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15176 14242 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15095 14242 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15014 14242 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14933 14242 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14852 14242 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14771 14242 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14690 14242 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14609 14242 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14527 14242 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14445 14242 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14363 14242 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14281 14242 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14199 14242 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14117 14242 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14035 14242 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 13953 14242 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 13871 14242 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 13789 14242 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 13707 14242 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 13625 14242 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 4432 14178 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 4346 14178 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 4260 14178 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 4174 14178 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 4088 14178 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 4002 14178 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 3916 14178 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 3830 14178 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 3744 14178 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 3658 14178 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 3572 14178 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 18539 14166 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 18457 14166 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 18375 14166 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 18293 14166 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 18211 14166 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 18129 14166 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 18047 14166 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 17965 14166 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 17883 14166 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 17801 14166 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 17719 14166 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 17637 14166 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 17555 14166 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 17473 14166 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 17391 14166 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 17309 14166 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 17227 14166 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 17145 14166 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 17063 14166 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 16981 14166 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 16899 14166 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 16817 14166 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 16735 14166 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 16653 14166 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 16571 14166 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 16472 14162 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 16391 14162 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 16310 14162 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 16229 14162 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 16148 14162 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 16067 14162 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15986 14162 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15905 14162 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15824 14162 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15743 14162 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15662 14162 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15581 14162 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15500 14162 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15419 14162 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15338 14162 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15257 14162 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15176 14162 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15095 14162 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15014 14162 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14933 14162 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14852 14162 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14771 14162 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14690 14162 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14609 14162 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14527 14162 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14445 14162 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14363 14162 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14281 14162 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14199 14162 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14117 14162 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14035 14162 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 13953 14162 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 13871 14162 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 13789 14162 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 13707 14162 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 13625 14162 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 4432 14097 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 4346 14097 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 4260 14097 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 4174 14097 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 4088 14097 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 4002 14097 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 3916 14097 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 3830 14097 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 3744 14097 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 3658 14097 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 3572 14097 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 18539 14084 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 18457 14084 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 18375 14084 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 18293 14084 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 18211 14084 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 18129 14084 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 18047 14084 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 17965 14084 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 17883 14084 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 17801 14084 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 17719 14084 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 17637 14084 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 17555 14084 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 17473 14084 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 17391 14084 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 17309 14084 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 17227 14084 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 17145 14084 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 17063 14084 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 16981 14084 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 16899 14084 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 16817 14084 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 16735 14084 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 16653 14084 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 16571 14084 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 16472 14082 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 16391 14082 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 16310 14082 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 16229 14082 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 16148 14082 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 16067 14082 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15986 14082 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15905 14082 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15824 14082 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15743 14082 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15662 14082 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15581 14082 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15500 14082 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15419 14082 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15338 14082 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15257 14082 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15176 14082 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15095 14082 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15014 14082 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14933 14082 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14852 14082 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14771 14082 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14690 14082 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14609 14082 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14527 14082 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14445 14082 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14363 14082 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14281 14082 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14199 14082 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14117 14082 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14035 14082 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 13953 14082 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 13871 14082 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 13789 14082 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 13707 14082 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 13625 14082 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 4432 14016 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 4346 14016 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 4260 14016 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 4174 14016 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 4088 14016 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 4002 14016 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 3916 14016 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 3830 14016 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 3744 14016 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 3658 14016 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 3572 14016 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 18539 14002 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 18457 14002 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 18375 14002 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 18293 14002 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 18211 14002 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 18129 14002 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 18047 14002 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 17965 14002 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 17883 14002 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 17801 14002 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 17719 14002 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 17637 14002 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 17555 14002 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 17473 14002 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 17391 14002 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 17309 14002 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 17227 14002 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 17145 14002 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 17063 14002 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16981 14002 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16899 14002 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16817 14002 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16735 14002 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16653 14002 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16571 14002 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16472 14002 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16391 14002 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16310 14002 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16229 14002 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16148 14002 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16067 14002 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15986 14002 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15905 14002 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15824 14002 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15743 14002 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15662 14002 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15581 14002 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15500 14002 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15419 14002 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15338 14002 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15257 14002 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15176 14002 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15095 14002 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15014 14002 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14933 14002 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14852 14002 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14771 14002 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14690 14002 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14609 14002 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14527 14002 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14445 14002 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14363 14002 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14281 14002 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14199 14002 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14117 14002 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14035 14002 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 13953 14002 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 13871 14002 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 13789 14002 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 13707 14002 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 13625 14002 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 4432 13935 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 4346 13935 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 4260 13935 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 4174 13935 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 4088 13935 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 4002 13935 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 3916 13935 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 3830 13935 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 3744 13935 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 3658 13935 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 3572 13935 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 16472 13922 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 16391 13922 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 16310 13922 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 16229 13922 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 16148 13922 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 16067 13922 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15986 13922 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15905 13922 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15824 13922 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15743 13922 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15662 13922 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15581 13922 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15500 13922 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15419 13922 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15338 13922 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15257 13922 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15176 13922 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15095 13922 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15014 13922 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14933 13922 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14852 13922 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14771 13922 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14690 13922 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14609 13922 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14527 13922 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14445 13922 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14363 13922 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14281 13922 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14199 13922 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14117 13922 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14035 13922 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 13953 13922 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 13871 13922 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 13789 13922 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 13707 13922 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 13625 13922 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 18539 13920 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 18457 13920 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 18375 13920 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 18293 13920 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 18211 13920 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 18129 13920 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 18047 13920 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 17965 13920 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 17883 13920 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 17801 13920 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 17719 13920 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 17637 13920 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 17555 13920 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 17473 13920 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 17391 13920 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 17309 13920 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 17227 13920 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 17145 13920 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 17063 13920 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 16981 13920 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 16899 13920 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 16817 13920 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 16735 13920 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 16653 13920 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 16571 13920 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 4432 13854 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 4346 13854 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 4260 13854 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 4174 13854 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 4088 13854 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 4002 13854 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 3916 13854 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 3830 13854 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 3744 13854 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 3658 13854 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 3572 13854 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 16472 13842 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 16391 13842 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 16310 13842 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 16229 13842 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 16148 13842 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 16067 13842 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15986 13842 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15905 13842 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15824 13842 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15743 13842 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15662 13842 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15581 13842 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15500 13842 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15419 13842 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15338 13842 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15257 13842 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15176 13842 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15095 13842 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15014 13842 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14933 13842 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14852 13842 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14771 13842 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14690 13842 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14609 13842 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14527 13842 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14445 13842 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14363 13842 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14281 13842 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14199 13842 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14117 13842 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14035 13842 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 13953 13842 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 13871 13842 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 13789 13842 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 13707 13842 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 13625 13842 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 18539 13838 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 18457 13838 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 18375 13838 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 18293 13838 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 18211 13838 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 18129 13838 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 18047 13838 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 17965 13838 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 17883 13838 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 17801 13838 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 17719 13838 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 17637 13838 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 17555 13838 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 17473 13838 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 17391 13838 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 17309 13838 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 17227 13838 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 17145 13838 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 17063 13838 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 16981 13838 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 16899 13838 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 16817 13838 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 16735 13838 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 16653 13838 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 16571 13838 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 4432 13773 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 4346 13773 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 4260 13773 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 4174 13773 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 4088 13773 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 4002 13773 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 3916 13773 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 3830 13773 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 3744 13773 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 3658 13773 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 3572 13773 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 16472 13762 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 16391 13762 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 16310 13762 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 16229 13762 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 16148 13762 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 16067 13762 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15986 13762 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15905 13762 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15824 13762 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15743 13762 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15662 13762 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15581 13762 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15500 13762 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15419 13762 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15338 13762 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15257 13762 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15176 13762 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15095 13762 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15014 13762 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14933 13762 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14852 13762 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14771 13762 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14690 13762 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14609 13762 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14527 13762 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14445 13762 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14363 13762 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14281 13762 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14199 13762 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14117 13762 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14035 13762 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 13953 13762 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 13871 13762 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 13789 13762 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 13707 13762 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 13625 13762 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 18539 13756 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 18457 13756 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 18375 13756 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 18293 13756 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 18211 13756 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 18129 13756 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 18047 13756 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 17965 13756 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 17883 13756 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 17801 13756 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 17719 13756 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 17637 13756 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 17555 13756 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 17473 13756 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 17391 13756 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 17309 13756 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 17227 13756 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 17145 13756 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 17063 13756 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 16981 13756 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 16899 13756 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 16817 13756 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 16735 13756 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 16653 13756 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 16571 13756 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 4432 13692 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 4346 13692 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 4260 13692 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 4174 13692 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 4088 13692 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 4002 13692 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 3916 13692 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 3830 13692 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 3744 13692 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 3658 13692 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 3572 13692 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 16472 13682 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 16391 13682 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 16310 13682 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 16229 13682 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 16148 13682 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 16067 13682 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15986 13682 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15905 13682 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15824 13682 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15743 13682 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15662 13682 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15581 13682 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15500 13682 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15419 13682 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15338 13682 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15257 13682 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15176 13682 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15095 13682 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15014 13682 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14933 13682 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14852 13682 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14771 13682 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14690 13682 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14609 13682 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14527 13682 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14445 13682 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14363 13682 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14281 13682 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14199 13682 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14117 13682 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14035 13682 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 13953 13682 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 13871 13682 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 13789 13682 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 13707 13682 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 13625 13682 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 18539 13674 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 18457 13674 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 18375 13674 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 18293 13674 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 18211 13674 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 18129 13674 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 18047 13674 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 17965 13674 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 17883 13674 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 17801 13674 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 17719 13674 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 17637 13674 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 17555 13674 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 17473 13674 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 17391 13674 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 17309 13674 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 17227 13674 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 17145 13674 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 17063 13674 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 16981 13674 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 16899 13674 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 16817 13674 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 16735 13674 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 16653 13674 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 16571 13674 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 4432 13611 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 4346 13611 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 4260 13611 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 4174 13611 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 4088 13611 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 4002 13611 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 3916 13611 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 3830 13611 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 3744 13611 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 3658 13611 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 3572 13611 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 16472 13602 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 16391 13602 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 16310 13602 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 16229 13602 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 16148 13602 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 16067 13602 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15986 13602 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15905 13602 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15824 13602 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15743 13602 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15662 13602 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15581 13602 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15500 13602 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15419 13602 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15338 13602 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15257 13602 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15176 13602 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15095 13602 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15014 13602 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14933 13602 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14852 13602 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14771 13602 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14690 13602 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14609 13602 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14527 13602 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14445 13602 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14363 13602 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14281 13602 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14199 13602 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14117 13602 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14035 13602 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 13953 13602 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 13871 13602 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 13789 13602 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 13707 13602 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 13625 13602 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 18539 13592 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 18457 13592 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 18375 13592 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 18293 13592 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 18211 13592 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 18129 13592 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 18047 13592 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 17965 13592 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 17883 13592 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 17801 13592 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 17719 13592 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 17637 13592 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 17555 13592 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 17473 13592 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 17391 13592 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 17309 13592 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 17227 13592 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 17145 13592 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 17063 13592 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 16981 13592 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 16899 13592 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 16817 13592 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 16735 13592 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 16653 13592 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 16571 13592 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 4432 13530 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 4346 13530 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 4260 13530 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 4174 13530 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 4088 13530 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 4002 13530 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 3916 13530 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 3830 13530 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 3744 13530 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 3658 13530 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 3572 13530 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 16472 13522 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 16391 13522 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 16310 13522 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 16229 13522 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 16148 13522 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 16067 13522 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15986 13522 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15905 13522 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15824 13522 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15743 13522 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15662 13522 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15581 13522 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15500 13522 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15419 13522 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15338 13522 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15257 13522 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15176 13522 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15095 13522 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15014 13522 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14933 13522 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14852 13522 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14771 13522 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14690 13522 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14609 13522 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14527 13522 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14445 13522 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14363 13522 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14281 13522 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14199 13522 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14117 13522 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14035 13522 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 13953 13522 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 13871 13522 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 13789 13522 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 13707 13522 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 13625 13522 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 18539 13510 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 18457 13510 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 18375 13510 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 18293 13510 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 18211 13510 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 18129 13510 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 18047 13510 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 17965 13510 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 17883 13510 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 17801 13510 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 17719 13510 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 17637 13510 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 17555 13510 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 17473 13510 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 17391 13510 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 17309 13510 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 17227 13510 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 17145 13510 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 17063 13510 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 16981 13510 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 16899 13510 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 16817 13510 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 16735 13510 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 16653 13510 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 16571 13510 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 4432 13449 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 4346 13449 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 4260 13449 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 4174 13449 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 4088 13449 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 4002 13449 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 3916 13449 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 3830 13449 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 3744 13449 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 3658 13449 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 3572 13449 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 16472 13442 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 16391 13442 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 16310 13442 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 16229 13442 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 16148 13442 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 16067 13442 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15986 13442 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15905 13442 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15824 13442 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15743 13442 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15662 13442 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15581 13442 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15500 13442 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15419 13442 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15338 13442 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15257 13442 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15176 13442 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15095 13442 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15014 13442 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14933 13442 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14852 13442 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14771 13442 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14690 13442 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14609 13442 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14527 13442 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14445 13442 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14363 13442 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14281 13442 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14199 13442 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14117 13442 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14035 13442 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 13953 13442 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 13871 13442 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 13789 13442 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 13707 13442 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 13625 13442 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 18539 13428 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 18457 13428 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 18375 13428 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 18293 13428 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 18211 13428 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 18129 13428 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 18047 13428 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 17965 13428 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 17883 13428 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 17801 13428 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 17719 13428 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 17637 13428 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 17555 13428 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 17473 13428 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 17391 13428 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 17309 13428 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 17227 13428 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 17145 13428 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 17063 13428 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 16981 13428 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 16899 13428 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 16817 13428 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 16735 13428 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 16653 13428 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 16571 13428 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 4432 13368 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 4346 13368 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 4260 13368 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 4174 13368 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 4088 13368 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 4002 13368 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 3916 13368 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 3830 13368 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 3744 13368 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 3658 13368 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 3572 13368 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 16472 13362 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 16391 13362 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 16310 13362 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 16229 13362 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 16148 13362 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 16067 13362 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15986 13362 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15905 13362 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15824 13362 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15743 13362 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15662 13362 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15581 13362 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15500 13362 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15419 13362 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15338 13362 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15257 13362 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15176 13362 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15095 13362 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15014 13362 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14933 13362 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14852 13362 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14771 13362 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14690 13362 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14609 13362 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14527 13362 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14445 13362 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14363 13362 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14281 13362 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14199 13362 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14117 13362 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14035 13362 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 13953 13362 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 13871 13362 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 13789 13362 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 13707 13362 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 13625 13362 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 18539 13346 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 18457 13346 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 18375 13346 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 18293 13346 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 18211 13346 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 18129 13346 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 18047 13346 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 17965 13346 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 17883 13346 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 17801 13346 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 17719 13346 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 17637 13346 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 17555 13346 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 17473 13346 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 17391 13346 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 17309 13346 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 17227 13346 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 17145 13346 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 17063 13346 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 16981 13346 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 16899 13346 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 16817 13346 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 16735 13346 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 16653 13346 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 16571 13346 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 4432 13287 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 4346 13287 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 4260 13287 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 4174 13287 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 4088 13287 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 4002 13287 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 3916 13287 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 3830 13287 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 3744 13287 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 3658 13287 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 3572 13287 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 16472 13282 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 16391 13282 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 16310 13282 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 16229 13282 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 16148 13282 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 16067 13282 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15986 13282 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15905 13282 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15824 13282 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15743 13282 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15662 13282 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15581 13282 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15500 13282 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15419 13282 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15338 13282 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15257 13282 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15176 13282 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15095 13282 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15014 13282 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14933 13282 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14852 13282 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14771 13282 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14690 13282 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14609 13282 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14527 13282 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14445 13282 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14363 13282 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14281 13282 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14199 13282 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14117 13282 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14035 13282 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 13953 13282 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 13871 13282 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 13789 13282 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 13707 13282 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 13625 13282 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 18539 13264 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 18457 13264 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 18375 13264 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 18293 13264 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 18211 13264 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 18129 13264 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 18047 13264 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 17965 13264 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 17883 13264 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 17801 13264 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 17719 13264 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 17637 13264 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 17555 13264 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 17473 13264 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 17391 13264 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 17309 13264 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 17227 13264 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 17145 13264 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 17063 13264 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 16981 13264 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 16899 13264 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 16817 13264 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 16735 13264 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 16653 13264 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 16571 13264 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 4432 13206 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 4346 13206 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 4260 13206 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 4174 13206 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 4088 13206 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 4002 13206 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 3916 13206 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 3830 13206 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 3744 13206 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 3658 13206 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 3572 13206 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 16472 13202 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 16391 13202 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 16310 13202 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 16229 13202 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 16148 13202 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 16067 13202 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15986 13202 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15905 13202 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15824 13202 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15743 13202 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15662 13202 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15581 13202 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15500 13202 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15419 13202 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15338 13202 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15257 13202 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15176 13202 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15095 13202 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15014 13202 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14933 13202 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14852 13202 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14771 13202 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14690 13202 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14609 13202 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14527 13202 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14445 13202 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14363 13202 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14281 13202 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14199 13202 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14117 13202 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14035 13202 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 13953 13202 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 13871 13202 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 13789 13202 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 13707 13202 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 13625 13202 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 18539 13182 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 18457 13182 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 18375 13182 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 18293 13182 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 18211 13182 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 18129 13182 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 18047 13182 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 17965 13182 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 17883 13182 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 17801 13182 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 17719 13182 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 17637 13182 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 17555 13182 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 17473 13182 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 17391 13182 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 17309 13182 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 17227 13182 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 17145 13182 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 17063 13182 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 16981 13182 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 16899 13182 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 16817 13182 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 16735 13182 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 16653 13182 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 16571 13182 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 4432 13125 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 4346 13125 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 4260 13125 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 4174 13125 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 4088 13125 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 4002 13125 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 3916 13125 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 3830 13125 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 3744 13125 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 3658 13125 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 3572 13125 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 16472 13122 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 16391 13122 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 16310 13122 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 16229 13122 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 16148 13122 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 16067 13122 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15986 13122 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15905 13122 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15824 13122 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15743 13122 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15662 13122 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15581 13122 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15500 13122 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15419 13122 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15338 13122 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15257 13122 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15176 13122 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15095 13122 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15014 13122 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14933 13122 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14852 13122 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14771 13122 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14690 13122 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14609 13122 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14527 13122 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14445 13122 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14363 13122 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14281 13122 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14199 13122 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14117 13122 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14035 13122 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 13953 13122 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 13871 13122 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 13789 13122 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 13707 13122 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 13625 13122 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 18539 13100 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 18457 13100 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 18375 13100 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 18293 13100 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 18211 13100 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 18129 13100 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 18047 13100 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 17965 13100 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 17883 13100 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 17801 13100 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 17719 13100 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 17637 13100 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 17555 13100 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 17473 13100 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 17391 13100 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 17309 13100 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 17227 13100 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 17145 13100 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 17063 13100 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 16981 13100 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 16899 13100 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 16817 13100 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 16735 13100 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 16653 13100 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 16571 13100 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 4432 13044 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 4346 13044 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 4260 13044 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 4174 13044 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 4088 13044 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 4002 13044 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 3916 13044 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 3830 13044 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 3744 13044 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 3658 13044 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 3572 13044 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 16472 13042 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 16391 13042 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 16310 13042 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 16229 13042 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 16148 13042 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 16067 13042 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15986 13042 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15905 13042 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15824 13042 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15743 13042 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15662 13042 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15581 13042 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15500 13042 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15419 13042 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15338 13042 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15257 13042 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15176 13042 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15095 13042 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15014 13042 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14933 13042 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14852 13042 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14771 13042 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14690 13042 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14609 13042 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14527 13042 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14445 13042 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14363 13042 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14281 13042 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14199 13042 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14117 13042 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14035 13042 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 13953 13042 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 13871 13042 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 13789 13042 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 13707 13042 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 13625 13042 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 18539 13018 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 18457 13018 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 18375 13018 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 18293 13018 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 18211 13018 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 18129 13018 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 18047 13018 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 17965 13018 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 17883 13018 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 17801 13018 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 17719 13018 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 17637 13018 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 17555 13018 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 17473 13018 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 17391 13018 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 17309 13018 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 17227 13018 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 17145 13018 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 17063 13018 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 16981 13018 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 16899 13018 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 16817 13018 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 16735 13018 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 16653 13018 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 16571 13018 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 4432 12963 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 4346 12963 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 4260 12963 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 4174 12963 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 4088 12963 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 4002 12963 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 3916 12963 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 3830 12963 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 3744 12963 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 3658 12963 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 3572 12963 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 16472 12962 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 16391 12962 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 16310 12962 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 16229 12962 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 16148 12962 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 16067 12962 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15986 12962 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15905 12962 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15824 12962 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15743 12962 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15662 12962 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15581 12962 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15500 12962 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15419 12962 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15338 12962 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15257 12962 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15176 12962 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15095 12962 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15014 12962 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14933 12962 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14852 12962 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14771 12962 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14690 12962 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14609 12962 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14527 12962 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14445 12962 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14363 12962 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14281 12962 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14199 12962 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14117 12962 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14035 12962 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 13953 12962 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 13871 12962 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 13789 12962 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 13707 12962 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 13625 12962 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 18539 12936 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 18457 12936 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 18375 12936 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 18293 12936 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 18211 12936 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 18129 12936 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 18047 12936 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 17965 12936 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 17883 12936 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 17801 12936 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 17719 12936 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 17637 12936 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 17555 12936 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 17473 12936 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 17391 12936 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 17309 12936 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 17227 12936 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 17145 12936 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 17063 12936 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 16981 12936 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 16899 12936 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 16817 12936 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 16735 12936 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 16653 12936 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 16571 12936 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 16472 12882 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 16391 12882 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 16310 12882 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 16229 12882 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 16148 12882 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 16067 12882 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15986 12882 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15905 12882 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15824 12882 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15743 12882 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15662 12882 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15581 12882 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15500 12882 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15419 12882 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15338 12882 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15257 12882 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15176 12882 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15095 12882 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15014 12882 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14933 12882 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14852 12882 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14771 12882 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14690 12882 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14609 12882 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14527 12882 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14445 12882 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14363 12882 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14281 12882 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14199 12882 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14117 12882 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14035 12882 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 13953 12882 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 13871 12882 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 13789 12882 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 13707 12882 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 13625 12882 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 4432 12882 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 4346 12882 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 4260 12882 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 4174 12882 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 4088 12882 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 4002 12882 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 3916 12882 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 3830 12882 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 3744 12882 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 3658 12882 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 3572 12882 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 18539 12854 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 18457 12854 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 18375 12854 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 18293 12854 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 18211 12854 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 18129 12854 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 18047 12854 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 17965 12854 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 17883 12854 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 17801 12854 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 17719 12854 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 17637 12854 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 17555 12854 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 17473 12854 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 17391 12854 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 17309 12854 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 17227 12854 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 17145 12854 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 17063 12854 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 16981 12854 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 16899 12854 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 16817 12854 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 16735 12854 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 16653 12854 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 16571 12854 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 16472 12802 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 16391 12802 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 16310 12802 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 16229 12802 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 16148 12802 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 16067 12802 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15986 12802 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15905 12802 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15824 12802 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15743 12802 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15662 12802 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15581 12802 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15500 12802 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15419 12802 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15338 12802 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15257 12802 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15176 12802 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15095 12802 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15014 12802 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14933 12802 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14852 12802 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14771 12802 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14690 12802 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14609 12802 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14527 12802 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14445 12802 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14363 12802 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14281 12802 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14199 12802 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14117 12802 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14035 12802 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 13953 12802 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 13871 12802 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 13789 12802 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 13707 12802 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 13625 12802 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 4432 12801 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 4346 12801 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 4260 12801 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 4174 12801 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 4088 12801 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 4002 12801 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 3916 12801 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 3830 12801 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 3744 12801 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 3658 12801 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 3572 12801 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 18539 12772 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 18457 12772 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 18375 12772 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 18293 12772 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 18211 12772 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 18129 12772 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 18047 12772 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 17965 12772 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 17883 12772 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 17801 12772 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 17719 12772 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 17637 12772 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 17555 12772 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 17473 12772 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 17391 12772 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 17309 12772 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 17227 12772 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 17145 12772 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 17063 12772 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 16981 12772 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 16899 12772 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 16817 12772 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 16735 12772 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 16653 12772 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 16571 12772 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 16472 12722 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 16391 12722 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 16310 12722 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 16229 12722 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 16148 12722 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 16067 12722 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15986 12722 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15905 12722 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15824 12722 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15743 12722 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15662 12722 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15581 12722 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15500 12722 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15419 12722 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15338 12722 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15257 12722 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15176 12722 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15095 12722 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15014 12722 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14933 12722 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14852 12722 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14771 12722 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14690 12722 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14609 12722 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14527 12722 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14445 12722 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14363 12722 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14281 12722 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14199 12722 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14117 12722 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14035 12722 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 13953 12722 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 13871 12722 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 13789 12722 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 13707 12722 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 13625 12722 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 4432 12720 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 4346 12720 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 4260 12720 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 4174 12720 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 4088 12720 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 4002 12720 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 3916 12720 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 3830 12720 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 3744 12720 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 3658 12720 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 3572 12720 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 18539 12690 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 18457 12690 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 18375 12690 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 18293 12690 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 18211 12690 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 18129 12690 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 18047 12690 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 17965 12690 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 17883 12690 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 17801 12690 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 17719 12690 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 17637 12690 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 17555 12690 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 17473 12690 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 17391 12690 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 17309 12690 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 17227 12690 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 17145 12690 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 17063 12690 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 16981 12690 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 16899 12690 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 16817 12690 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 16735 12690 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 16653 12690 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 16571 12690 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 16472 12642 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 16391 12642 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 16310 12642 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 16229 12642 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 16148 12642 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 16067 12642 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15986 12642 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15905 12642 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15824 12642 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15743 12642 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15662 12642 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15581 12642 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15500 12642 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15419 12642 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15338 12642 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15257 12642 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15176 12642 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15095 12642 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15014 12642 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14933 12642 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14852 12642 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14771 12642 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14690 12642 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14609 12642 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14527 12642 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14445 12642 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14363 12642 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14281 12642 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14199 12642 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14117 12642 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14035 12642 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 13953 12642 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 13871 12642 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 13789 12642 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 13707 12642 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 13625 12642 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 4432 12639 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 4346 12639 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 4260 12639 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 4174 12639 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 4088 12639 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 4002 12639 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 3916 12639 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 3830 12639 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 3744 12639 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 3658 12639 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 3572 12639 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 18539 12608 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 18457 12608 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 18375 12608 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 18293 12608 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 18211 12608 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 18129 12608 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 18047 12608 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 17965 12608 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 17883 12608 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 17801 12608 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 17719 12608 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 17637 12608 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 17555 12608 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 17473 12608 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 17391 12608 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 17309 12608 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 17227 12608 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 17145 12608 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 17063 12608 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 16981 12608 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 16899 12608 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 16817 12608 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 16735 12608 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 16653 12608 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 16571 12608 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 16472 12562 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 16391 12562 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 16310 12562 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 16229 12562 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 16148 12562 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 16067 12562 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15986 12562 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15905 12562 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15824 12562 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15743 12562 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15662 12562 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15581 12562 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15500 12562 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15419 12562 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15338 12562 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15257 12562 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15176 12562 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15095 12562 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15014 12562 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14933 12562 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14852 12562 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14771 12562 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14690 12562 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14609 12562 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14527 12562 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14445 12562 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14363 12562 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14281 12562 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14199 12562 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14117 12562 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14035 12562 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 13953 12562 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 13871 12562 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 13789 12562 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 13707 12562 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 13625 12562 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 4432 12558 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 4346 12558 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 4260 12558 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 4174 12558 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 4088 12558 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 4002 12558 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 3916 12558 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 3830 12558 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 3744 12558 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 3658 12558 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 3572 12558 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 18539 12526 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 18457 12526 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 18375 12526 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 18293 12526 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 18211 12526 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 18129 12526 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 18047 12526 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 17965 12526 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 17883 12526 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 17801 12526 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 17719 12526 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 17637 12526 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 17555 12526 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 17473 12526 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 17391 12526 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 17309 12526 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 17227 12526 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 17145 12526 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 17063 12526 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 16981 12526 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 16899 12526 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 16817 12526 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 16735 12526 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 16653 12526 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 16571 12526 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 16472 12482 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 16391 12482 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 16310 12482 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 16229 12482 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 16148 12482 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 16067 12482 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15986 12482 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15905 12482 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15824 12482 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15743 12482 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15662 12482 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15581 12482 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15500 12482 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15419 12482 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15338 12482 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15257 12482 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15176 12482 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15095 12482 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15014 12482 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14933 12482 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14852 12482 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14771 12482 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14690 12482 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14609 12482 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14527 12482 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14445 12482 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14363 12482 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14281 12482 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14199 12482 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14117 12482 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14035 12482 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 13953 12482 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 13871 12482 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 13789 12482 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 13707 12482 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 13625 12482 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 4432 12477 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 4346 12477 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 4260 12477 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 4174 12477 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 4088 12477 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 4002 12477 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 3916 12477 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 3830 12477 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 3744 12477 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 3658 12477 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 3572 12477 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 18539 12445 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 18457 12445 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 18375 12445 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 18293 12445 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 18211 12445 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 18129 12445 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 18047 12445 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 17965 12445 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 17883 12445 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 17801 12445 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 17719 12445 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 17637 12445 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 17555 12445 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 17473 12445 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 17391 12445 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 17309 12445 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 17227 12445 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 17145 12445 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 17063 12445 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 16981 12445 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 16899 12445 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 16817 12445 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 16735 12445 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 16653 12445 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 16571 12445 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 16472 12402 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 16391 12402 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 16310 12402 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 16229 12402 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 16148 12402 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 16067 12402 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15986 12402 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15905 12402 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15824 12402 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15743 12402 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15662 12402 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15581 12402 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15500 12402 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15419 12402 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15338 12402 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15257 12402 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15176 12402 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15095 12402 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15014 12402 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14933 12402 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14852 12402 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14771 12402 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14690 12402 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14609 12402 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14527 12402 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14445 12402 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14363 12402 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14281 12402 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14199 12402 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14117 12402 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14035 12402 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 13953 12402 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 13871 12402 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 13789 12402 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 13707 12402 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 13625 12402 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 4432 12396 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 4346 12396 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 4260 12396 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 4174 12396 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 4088 12396 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 4002 12396 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 3916 12396 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 3830 12396 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 3744 12396 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 3658 12396 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 3572 12396 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 18539 12364 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 18457 12364 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 18375 12364 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 18293 12364 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 18211 12364 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 18129 12364 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 18047 12364 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 17965 12364 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 17883 12364 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 17801 12364 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 17719 12364 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 17637 12364 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 17555 12364 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 17473 12364 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 17391 12364 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 17309 12364 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 17227 12364 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 17145 12364 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 17063 12364 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 16981 12364 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 16899 12364 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 16817 12364 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 16735 12364 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 16653 12364 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 16571 12364 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 16472 12322 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 16391 12322 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 16310 12322 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 16229 12322 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 16148 12322 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 16067 12322 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15986 12322 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15905 12322 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15824 12322 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15743 12322 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15662 12322 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15581 12322 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15500 12322 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15419 12322 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15338 12322 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15257 12322 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15176 12322 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15095 12322 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15014 12322 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14933 12322 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14852 12322 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14771 12322 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14690 12322 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14609 12322 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14527 12322 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14445 12322 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14363 12322 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14281 12322 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14199 12322 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14117 12322 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14035 12322 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 13953 12322 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 13871 12322 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 13789 12322 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 13707 12322 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 13625 12322 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 4432 12315 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 4346 12315 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 4260 12315 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 4174 12315 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 4088 12315 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 4002 12315 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 3916 12315 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 3830 12315 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 3744 12315 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 3658 12315 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 3572 12315 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 18539 12283 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 18457 12283 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 18375 12283 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 18293 12283 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 18211 12283 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 18129 12283 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 18047 12283 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 17965 12283 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 17883 12283 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 17801 12283 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 17719 12283 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 17637 12283 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 17555 12283 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 17473 12283 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 17391 12283 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 17309 12283 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 17227 12283 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 17145 12283 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 17063 12283 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 16981 12283 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 16899 12283 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 16817 12283 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 16735 12283 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 16653 12283 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 16571 12283 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 16472 12242 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 16391 12242 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 16310 12242 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 16229 12242 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 16148 12242 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 16067 12242 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15986 12242 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15905 12242 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15824 12242 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15743 12242 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15662 12242 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15581 12242 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15500 12242 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15419 12242 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15338 12242 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15257 12242 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15176 12242 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15095 12242 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15014 12242 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14933 12242 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14852 12242 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14771 12242 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14690 12242 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14609 12242 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14527 12242 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14445 12242 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14363 12242 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14281 12242 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14199 12242 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14117 12242 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14035 12242 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 13953 12242 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 13871 12242 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 13789 12242 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 13707 12242 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 13625 12242 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 4432 12234 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 4346 12234 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 4260 12234 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 4174 12234 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 4088 12234 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 4002 12234 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 3916 12234 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 3830 12234 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 3744 12234 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 3658 12234 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 3572 12234 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12147 18289 12187 18329 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12147 18203 12187 18243 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12143 18111 12183 18151 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12143 18025 12183 18065 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12143 17939 12183 17979 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12143 17853 12183 17893 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12143 17767 12183 17807 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12143 17682 12183 17722 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 16472 12162 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 16391 12162 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 16310 12162 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 16229 12162 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 16148 12162 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 16067 12162 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15986 12162 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15905 12162 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15824 12162 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15743 12162 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15662 12162 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15581 12162 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15500 12162 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15419 12162 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15338 12162 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15257 12162 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15176 12162 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15095 12162 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15014 12162 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14933 12162 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14852 12162 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14771 12162 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14690 12162 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14609 12162 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14527 12162 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14445 12162 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14363 12162 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14281 12162 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14199 12162 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14117 12162 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14035 12162 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 13953 12162 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 13871 12162 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 13789 12162 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 13707 12162 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 13625 12162 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12118 17575 12158 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12118 17494 12158 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12118 17413 12158 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12118 17332 12158 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12118 17251 12158 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12118 17171 12158 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12118 17091 12158 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12118 17011 12158 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12118 16931 12158 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12118 16851 12158 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12118 16771 12158 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12118 16691 12158 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12118 16611 12158 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 4432 12153 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 4346 12153 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 4260 12153 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 4174 12153 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 4088 12153 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 4002 12153 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 3916 12153 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 3830 12153 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 3744 12153 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 3658 12153 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 3572 12153 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12061 18111 12101 18151 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12061 18025 12101 18065 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12061 17939 12101 17979 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12061 17853 12101 17893 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12061 17767 12101 17807 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12061 17682 12101 17722 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 16472 12082 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 16391 12082 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 16310 12082 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 16229 12082 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 16148 12082 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 16067 12082 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15986 12082 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15905 12082 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15824 12082 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15743 12082 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15662 12082 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15581 12082 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15500 12082 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15419 12082 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15338 12082 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15257 12082 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15176 12082 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15095 12082 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15014 12082 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14933 12082 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14852 12082 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14771 12082 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14690 12082 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14609 12082 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14527 12082 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14445 12082 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14363 12082 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14281 12082 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14199 12082 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14117 12082 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14035 12082 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 13953 12082 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 13871 12082 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 13789 12082 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 13707 12082 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 13625 12082 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12036 17575 12076 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12036 17494 12076 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12036 17413 12076 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12036 17332 12076 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12036 17251 12076 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12036 17171 12076 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12036 17091 12076 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12036 17011 12076 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12036 16931 12076 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12036 16851 12076 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12036 16771 12076 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12036 16691 12076 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12036 16611 12076 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 4432 12072 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 4346 12072 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 4260 12072 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 4174 12072 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 4088 12072 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 4002 12072 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 3916 12072 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 3830 12072 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 3744 12072 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 3658 12072 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 3572 12072 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11991 18289 12031 18329 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11991 18203 12031 18243 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11979 18111 12019 18151 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11979 18025 12019 18065 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11979 17939 12019 17979 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11979 17853 12019 17893 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11979 17767 12019 17807 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11979 17682 12019 17722 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 16472 12002 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 16391 12002 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 16310 12002 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 16229 12002 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 16148 12002 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 16067 12002 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15986 12002 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15905 12002 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15824 12002 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15743 12002 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15662 12002 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15581 12002 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15500 12002 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15419 12002 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15338 12002 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15257 12002 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15176 12002 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15095 12002 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15014 12002 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14933 12002 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14852 12002 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14771 12002 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14690 12002 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14609 12002 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14527 12002 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14445 12002 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14363 12002 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14281 12002 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14199 12002 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14117 12002 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14035 12002 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 13953 12002 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 13871 12002 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 13789 12002 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 13707 12002 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 13625 12002 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11954 17575 11994 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11954 17494 11994 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11954 17413 11994 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11954 17332 11994 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11954 17251 11994 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11954 17171 11994 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11954 17091 11994 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11954 17011 11994 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11954 16931 11994 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11954 16851 11994 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11954 16771 11994 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11954 16691 11994 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11954 16611 11994 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 4432 11991 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 4346 11991 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 4260 11991 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 4174 11991 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 4088 11991 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 4002 11991 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 3916 11991 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 3830 11991 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 3744 11991 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 3658 11991 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 3572 11991 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11897 18111 11937 18151 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11897 18025 11937 18065 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11897 17939 11937 17979 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11897 17853 11937 17893 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11897 17767 11937 17807 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11897 17682 11937 17722 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 16472 11922 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 16391 11922 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 16310 11922 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 16229 11922 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 16148 11922 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 16067 11922 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15986 11922 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15905 11922 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15824 11922 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15743 11922 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15662 11922 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15581 11922 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15500 11922 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15419 11922 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15338 11922 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15257 11922 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15176 11922 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15095 11922 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15014 11922 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14933 11922 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14852 11922 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14771 11922 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14690 11922 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14609 11922 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14527 11922 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14445 11922 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14363 11922 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14281 11922 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14199 11922 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14117 11922 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14035 11922 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 13953 11922 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 13871 11922 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 13789 11922 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 13707 11922 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 13625 11922 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11872 17575 11912 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11872 17494 11912 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11872 17413 11912 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11872 17332 11912 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11872 17251 11912 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11872 17171 11912 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11872 17091 11912 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11872 17011 11912 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11872 16931 11912 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11872 16851 11912 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11872 16771 11912 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11872 16691 11912 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11872 16611 11912 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 4432 11910 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 4346 11910 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 4260 11910 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 4174 11910 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 4088 11910 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 4002 11910 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 3916 11910 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 3830 11910 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 3744 11910 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 3658 11910 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 3572 11910 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11815 18111 11855 18151 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11815 18025 11855 18065 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11815 17939 11855 17979 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11815 17853 11855 17893 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11815 17767 11855 17807 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11815 17682 11855 17722 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 16472 11842 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 16391 11842 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 16310 11842 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 16229 11842 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 16148 11842 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 16067 11842 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15986 11842 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15905 11842 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15824 11842 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15743 11842 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15662 11842 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15581 11842 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15500 11842 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15419 11842 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15338 11842 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15257 11842 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15176 11842 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15095 11842 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15014 11842 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14933 11842 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14852 11842 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14771 11842 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14690 11842 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14609 11842 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14527 11842 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14445 11842 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14363 11842 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14281 11842 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14199 11842 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14117 11842 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14035 11842 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 13953 11842 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 13871 11842 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 13789 11842 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 13707 11842 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 13625 11842 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 17575 11830 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 17494 11830 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 17413 11830 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 17332 11830 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 17251 11830 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 17171 11830 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 17091 11830 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 17011 11830 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 16931 11830 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 16851 11830 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 16771 11830 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 16691 11830 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 16611 11830 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 4432 11829 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 4346 11829 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 4260 11829 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 4174 11829 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 4088 11829 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 4002 11829 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 3916 11829 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 3830 11829 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 3744 11829 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 3658 11829 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 3572 11829 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 16472 11762 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 16391 11762 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 16310 11762 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 16229 11762 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 16148 11762 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 16067 11762 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15986 11762 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15905 11762 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15824 11762 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15743 11762 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15662 11762 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15581 11762 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15500 11762 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15419 11762 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15338 11762 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15257 11762 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15176 11762 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15095 11762 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15014 11762 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14933 11762 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14852 11762 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14771 11762 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14690 11762 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14609 11762 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14527 11762 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14445 11762 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14363 11762 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14281 11762 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14199 11762 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14117 11762 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14035 11762 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 13953 11762 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 13871 11762 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 13789 11762 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 13707 11762 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 13625 11762 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11715 17853 11755 17893 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11715 17769 11755 17809 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11715 17686 11755 17726 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 17575 11748 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 17494 11748 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 17413 11748 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 17332 11748 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 17251 11748 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 17171 11748 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 17091 11748 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 17011 11748 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 16931 11748 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 16851 11748 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 16771 11748 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 16691 11748 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 16611 11748 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 4432 11748 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 4346 11748 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 4260 11748 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 4174 11748 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 4088 11748 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 4002 11748 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 3916 11748 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 3830 11748 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 3744 11748 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 3658 11748 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 3572 11748 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 16472 11682 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 16391 11682 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 16310 11682 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 16229 11682 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 16148 11682 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 16067 11682 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15986 11682 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15905 11682 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15824 11682 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15743 11682 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15662 11682 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15581 11682 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15500 11682 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15419 11682 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15338 11682 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15257 11682 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15176 11682 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15095 11682 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15014 11682 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14933 11682 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14852 11682 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14771 11682 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14690 11682 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14609 11682 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14527 11682 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14445 11682 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14363 11682 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14281 11682 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14199 11682 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14117 11682 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14035 11682 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 13953 11682 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 13871 11682 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 13789 11682 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 13707 11682 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 13625 11682 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 4432 11667 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 4346 11667 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 4260 11667 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 4174 11667 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 4088 11667 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 4002 11667 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 3916 11667 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 3830 11667 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 3744 11667 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 3658 11667 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 3572 11667 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11626 17575 11666 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11626 17494 11666 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11626 17413 11666 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11626 17332 11666 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11626 17251 11666 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11626 17171 11666 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11626 17091 11666 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11626 17011 11666 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11626 16931 11666 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11626 16851 11666 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11626 16771 11666 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11626 16691 11666 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11626 16611 11666 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 16472 11602 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 16391 11602 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 16310 11602 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 16229 11602 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 16148 11602 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 16067 11602 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15986 11602 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15905 11602 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15824 11602 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15743 11602 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15662 11602 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15581 11602 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15500 11602 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15419 11602 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15338 11602 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15257 11602 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15176 11602 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15095 11602 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15014 11602 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14933 11602 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14852 11602 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14771 11602 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14690 11602 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14609 11602 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14527 11602 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14445 11602 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14363 11602 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14281 11602 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14199 11602 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14117 11602 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14035 11602 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 13953 11602 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 13871 11602 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 13789 11602 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 13707 11602 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 13625 11602 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11559 17853 11599 17893 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11559 17769 11599 17809 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11559 17686 11599 17726 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 4432 11586 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 4346 11586 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 4260 11586 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 4174 11586 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 4088 11586 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 4002 11586 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 3916 11586 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 3830 11586 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 3744 11586 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 3658 11586 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 3572 11586 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11544 17575 11584 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11544 17494 11584 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11544 17413 11584 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11544 17332 11584 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11544 17251 11584 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11544 17171 11584 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11544 17091 11584 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11544 17011 11584 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11544 16931 11584 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11544 16851 11584 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11544 16771 11584 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11544 16691 11584 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11544 16611 11584 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 16472 11522 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 16391 11522 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 16310 11522 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 16229 11522 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 16148 11522 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 16067 11522 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15986 11522 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15905 11522 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15824 11522 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15743 11522 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15662 11522 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15581 11522 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15500 11522 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15419 11522 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15338 11522 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15257 11522 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15176 11522 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15095 11522 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15014 11522 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14933 11522 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14852 11522 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14771 11522 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14690 11522 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14609 11522 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14527 11522 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14445 11522 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14363 11522 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14281 11522 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14199 11522 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14117 11522 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14035 11522 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 13953 11522 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 13871 11522 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 13789 11522 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 13707 11522 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 13625 11522 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 4432 11505 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 4346 11505 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 4260 11505 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 4174 11505 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 4088 11505 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 4002 11505 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 3916 11505 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 3830 11505 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 3744 11505 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 3658 11505 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 3572 11505 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11462 17575 11502 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11462 17494 11502 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11462 17413 11502 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11462 17332 11502 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11462 17251 11502 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11462 17171 11502 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11462 17091 11502 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11462 17011 11502 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11462 16931 11502 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11462 16851 11502 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11462 16771 11502 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11462 16691 11502 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11462 16611 11502 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 16472 11442 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 16391 11442 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 16310 11442 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 16229 11442 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 16148 11442 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 16067 11442 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15986 11442 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15905 11442 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15824 11442 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15743 11442 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15662 11442 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15581 11442 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15500 11442 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15419 11442 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15338 11442 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15257 11442 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15176 11442 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15095 11442 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15014 11442 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14933 11442 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14852 11442 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14771 11442 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14690 11442 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14609 11442 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14527 11442 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14445 11442 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14363 11442 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14281 11442 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14199 11442 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14117 11442 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14035 11442 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 13953 11442 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 13871 11442 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 13789 11442 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 13707 11442 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 13625 11442 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 4432 11424 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 4346 11424 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 4260 11424 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 4174 11424 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 4088 11424 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 4002 11424 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 3916 11424 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 3830 11424 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 3744 11424 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 3658 11424 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 3572 11424 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11380 17575 11420 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11380 17494 11420 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11380 17413 11420 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11380 17332 11420 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11380 17251 11420 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11380 17171 11420 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11380 17091 11420 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11380 17011 11420 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11380 16931 11420 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11380 16851 11420 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11380 16771 11420 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11380 16691 11420 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11380 16611 11420 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 16472 11362 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 16391 11362 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 16310 11362 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 16229 11362 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 16148 11362 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 16067 11362 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15986 11362 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15905 11362 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15824 11362 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15743 11362 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15662 11362 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15581 11362 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15500 11362 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15419 11362 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15338 11362 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15257 11362 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15176 11362 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15095 11362 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15014 11362 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14933 11362 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14852 11362 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14771 11362 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14690 11362 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14609 11362 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14527 11362 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14445 11362 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14363 11362 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14281 11362 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14199 11362 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14117 11362 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14035 11362 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 13953 11362 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 13871 11362 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 13789 11362 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 13707 11362 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 13625 11362 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 4432 11343 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 4346 11343 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 4260 11343 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 4174 11343 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 4088 11343 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 4002 11343 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 3916 11343 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 3830 11343 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 3744 11343 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 3658 11343 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 3572 11343 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11298 17575 11338 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11298 17494 11338 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11298 17413 11338 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11298 17332 11338 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11298 17251 11338 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11298 17171 11338 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11298 17091 11338 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11298 17011 11338 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11298 16931 11338 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11298 16851 11338 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11298 16771 11338 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11298 16691 11338 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11298 16611 11338 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 16472 11282 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 16391 11282 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 16310 11282 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 16229 11282 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 16148 11282 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 16067 11282 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15986 11282 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15905 11282 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15824 11282 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15743 11282 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15662 11282 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15581 11282 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15500 11282 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15419 11282 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15338 11282 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15257 11282 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15176 11282 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15095 11282 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15014 11282 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14933 11282 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14852 11282 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14771 11282 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14690 11282 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14609 11282 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14527 11282 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14445 11282 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14363 11282 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14281 11282 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14199 11282 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14117 11282 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14035 11282 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 13953 11282 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 13871 11282 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 13789 11282 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 13707 11282 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 13625 11282 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 4432 11262 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 4346 11262 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 4260 11262 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 4174 11262 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 4088 11262 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 4002 11262 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 3916 11262 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 3830 11262 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 3744 11262 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 3658 11262 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 3572 11262 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11199 17350 11239 17390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11199 17262 11239 17302 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11199 17175 11239 17215 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 16472 11202 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 16391 11202 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 16310 11202 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 16229 11202 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 16148 11202 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 16067 11202 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15986 11202 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15905 11202 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15824 11202 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15743 11202 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15662 11202 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15581 11202 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15500 11202 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15419 11202 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15338 11202 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15257 11202 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15176 11202 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15095 11202 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15014 11202 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14933 11202 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14852 11202 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14771 11202 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14690 11202 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14609 11202 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14527 11202 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14445 11202 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14363 11202 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14281 11202 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14199 11202 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14117 11202 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14035 11202 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 13953 11202 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 13871 11202 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 13789 11202 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 13707 11202 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 13625 11202 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11161 17065 11201 17105 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11161 16972 11201 17012 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11161 16879 11201 16919 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11161 16786 11201 16826 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11161 16694 11201 16734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11161 16602 11201 16642 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 4432 11181 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 4346 11181 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 4260 11181 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 4174 11181 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 4088 11181 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 4002 11181 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 3916 11181 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 3830 11181 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 3744 11181 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 3658 11181 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 3572 11181 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 16472 11122 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 16391 11122 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 16310 11122 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 16229 11122 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 16148 11122 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 16067 11122 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15986 11122 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15905 11122 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15824 11122 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15743 11122 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15662 11122 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15581 11122 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15500 11122 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15419 11122 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15338 11122 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15257 11122 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15176 11122 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15095 11122 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15014 11122 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14933 11122 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14852 11122 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14771 11122 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14690 11122 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14609 11122 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14527 11122 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14445 11122 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14363 11122 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14281 11122 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14199 11122 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14117 11122 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14035 11122 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 13953 11122 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 13871 11122 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 13789 11122 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 13707 11122 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 13625 11122 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11065 17065 11105 17105 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11065 16972 11105 17012 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11065 16879 11105 16919 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11065 16786 11105 16826 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11065 16694 11105 16734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11065 16602 11105 16642 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 4432 11100 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 4346 11100 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 4260 11100 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 4174 11100 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 4088 11100 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 4002 11100 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 3916 11100 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 3830 11100 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 3744 11100 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 3658 11100 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 3572 11100 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11051 17350 11091 17390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11051 17262 11091 17302 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11051 17175 11091 17215 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 16472 11042 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 16391 11042 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 16310 11042 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 16229 11042 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 16148 11042 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 16067 11042 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15986 11042 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15905 11042 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15824 11042 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15743 11042 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15662 11042 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15581 11042 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15500 11042 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15419 11042 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15338 11042 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15257 11042 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15176 11042 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15095 11042 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15014 11042 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14933 11042 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14852 11042 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14771 11042 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14690 11042 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14609 11042 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14527 11042 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14445 11042 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14363 11042 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14281 11042 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14199 11042 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14117 11042 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14035 11042 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 13953 11042 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 13871 11042 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 13789 11042 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 13707 11042 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 13625 11042 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 4432 11019 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 4346 11019 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 4260 11019 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 4174 11019 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 4088 11019 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 4002 11019 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 3916 11019 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 3830 11019 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 3744 11019 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 3658 11019 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 3572 11019 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10969 17065 11009 17105 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10969 16972 11009 17012 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10969 16879 11009 16919 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10969 16786 11009 16826 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10969 16694 11009 16734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10969 16602 11009 16642 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 16472 10962 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 16391 10962 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 16310 10962 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 16229 10962 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 16148 10962 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 16067 10962 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15986 10962 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15905 10962 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15824 10962 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15743 10962 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15662 10962 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15581 10962 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15500 10962 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15419 10962 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15338 10962 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15257 10962 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15176 10962 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15095 10962 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15014 10962 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14933 10962 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14852 10962 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14771 10962 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14690 10962 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14609 10962 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14527 10962 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14445 10962 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14363 10962 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14281 10962 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14199 10962 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14117 10962 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14035 10962 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 13953 10962 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 13871 10962 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 13789 10962 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 13707 10962 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 13625 10962 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 4432 10938 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 4346 10938 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 4260 10938 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 4174 10938 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 4088 10938 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 4002 10938 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 3916 10938 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 3830 10938 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 3744 10938 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 3658 10938 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 3572 10938 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10873 17065 10913 17105 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10873 16972 10913 17012 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10873 16879 10913 16919 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10873 16786 10913 16826 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10873 16694 10913 16734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10873 16602 10913 16642 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 16472 10882 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 16391 10882 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 16310 10882 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 16229 10882 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 16148 10882 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 16067 10882 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15986 10882 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15905 10882 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15824 10882 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15743 10882 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15662 10882 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15581 10882 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15500 10882 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15419 10882 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15338 10882 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15257 10882 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15176 10882 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15095 10882 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15014 10882 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14933 10882 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14852 10882 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14771 10882 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14690 10882 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14609 10882 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14527 10882 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14445 10882 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14363 10882 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14281 10882 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14199 10882 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14117 10882 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14035 10882 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 13953 10882 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 13871 10882 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 13789 10882 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 13707 10882 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 13625 10882 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 4432 10857 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 4346 10857 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 4260 10857 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 4174 10857 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 4088 10857 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 4002 10857 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 3916 10857 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 3830 10857 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 3744 10857 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 3658 10857 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 3572 10857 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10777 17065 10817 17105 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10777 16972 10817 17012 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10777 16879 10817 16919 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10777 16786 10817 16826 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10777 16694 10817 16734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10777 16602 10817 16642 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 16472 10802 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 16391 10802 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 16310 10802 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 16229 10802 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 16148 10802 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 16067 10802 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15986 10802 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15905 10802 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15824 10802 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15743 10802 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15662 10802 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15581 10802 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15500 10802 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15419 10802 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15338 10802 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15257 10802 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15176 10802 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15095 10802 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15014 10802 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14933 10802 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14852 10802 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14771 10802 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14690 10802 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14609 10802 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14527 10802 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14445 10802 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14363 10802 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14281 10802 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14199 10802 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14117 10802 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14035 10802 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 13953 10802 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 13871 10802 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 13789 10802 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 13707 10802 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 13625 10802 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 4432 10776 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 4346 10776 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 4260 10776 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 4174 10776 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 4088 10776 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 4002 10776 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 3916 10776 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 3830 10776 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 3744 10776 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 3658 10776 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 3572 10776 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 16472 10722 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 16391 10722 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 16310 10722 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 16229 10722 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 16148 10722 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 16067 10722 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15986 10722 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15905 10722 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15824 10722 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15743 10722 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15662 10722 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15581 10722 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15500 10722 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15419 10722 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15338 10722 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15257 10722 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15176 10722 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15095 10722 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15014 10722 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14933 10722 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14852 10722 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14771 10722 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14690 10722 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14609 10722 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14527 10722 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14445 10722 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14363 10722 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14281 10722 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14199 10722 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14117 10722 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14035 10722 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 13953 10722 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 13871 10722 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 13789 10722 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 13707 10722 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 13625 10722 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10668 16804 10708 16844 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10668 16694 10708 16734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10668 16584 10708 16624 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 4432 10695 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 4346 10695 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 4260 10695 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 4174 10695 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 4088 10695 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 4002 10695 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 3916 10695 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 3830 10695 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 3744 10695 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 3658 10695 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 3572 10695 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 16472 10642 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 16391 10642 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 16310 10642 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 16229 10642 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 16148 10642 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 16067 10642 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15986 10642 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15905 10642 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15824 10642 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15743 10642 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15662 10642 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15581 10642 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15500 10642 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15419 10642 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15338 10642 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15257 10642 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15176 10642 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15095 10642 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15014 10642 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14933 10642 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14852 10642 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14771 10642 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14690 10642 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14609 10642 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14527 10642 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14445 10642 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14363 10642 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14281 10642 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14199 10642 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14117 10642 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14035 10642 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 13953 10642 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 13871 10642 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 13789 10642 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 13707 10642 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 13625 10642 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 4432 10614 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 4346 10614 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 4260 10614 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 4174 10614 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 4088 10614 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 4002 10614 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 3916 10614 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 3830 10614 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 3744 10614 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 3658 10614 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 3572 10614 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 16472 10562 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 16391 10562 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 16310 10562 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 16229 10562 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 16148 10562 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 16067 10562 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15986 10562 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15905 10562 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15824 10562 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15743 10562 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15662 10562 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15581 10562 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15500 10562 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15419 10562 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15338 10562 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15257 10562 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15176 10562 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15095 10562 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15014 10562 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14933 10562 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14852 10562 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14771 10562 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14690 10562 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14609 10562 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14527 10562 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14445 10562 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14363 10562 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14281 10562 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14199 10562 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14117 10562 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14035 10562 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 13953 10562 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 13871 10562 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 13789 10562 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 13707 10562 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 13625 10562 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 16804 10550 16844 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 16694 10550 16734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 16584 10550 16624 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 4432 10533 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 4346 10533 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 4260 10533 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 4174 10533 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 4088 10533 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 4002 10533 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 3916 10533 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 3830 10533 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 3744 10533 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 3658 10533 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 3572 10533 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 16472 10482 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 16391 10482 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 16310 10482 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 16229 10482 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 16148 10482 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 16067 10482 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15986 10482 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15905 10482 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15824 10482 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15743 10482 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15662 10482 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15581 10482 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15500 10482 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15419 10482 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15338 10482 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15257 10482 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15176 10482 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15095 10482 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15014 10482 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14933 10482 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14852 10482 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14771 10482 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14690 10482 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14609 10482 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14527 10482 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14445 10482 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14363 10482 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14281 10482 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14199 10482 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14117 10482 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14035 10482 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 13953 10482 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 13871 10482 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 13789 10482 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 13707 10482 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 13625 10482 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 4432 10452 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 4346 10452 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 4260 10452 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 4174 10452 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 4088 10452 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 4002 10452 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 3916 10452 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 3830 10452 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 3744 10452 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 3658 10452 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 3572 10452 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 16472 10402 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 16391 10402 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 16310 10402 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 16229 10402 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 16148 10402 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 16067 10402 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15986 10402 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15905 10402 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15824 10402 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15743 10402 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15662 10402 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15581 10402 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15500 10402 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15419 10402 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15338 10402 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15257 10402 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15176 10402 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15095 10402 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15014 10402 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14933 10402 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14852 10402 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14771 10402 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14690 10402 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14609 10402 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14527 10402 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14445 10402 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14363 10402 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14281 10402 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14199 10402 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14117 10402 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14035 10402 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 13953 10402 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 13871 10402 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 13789 10402 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 13707 10402 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 13625 10402 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 4432 10371 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 4346 10371 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 4260 10371 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 4174 10371 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 4088 10371 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 4002 10371 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 3916 10371 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 3830 10371 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 3744 10371 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 3658 10371 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 3572 10371 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 16472 10322 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 16391 10322 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 16310 10322 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 16229 10322 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 16148 10322 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 16067 10322 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15986 10322 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15905 10322 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15824 10322 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15743 10322 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15662 10322 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15581 10322 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15500 10322 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15419 10322 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15338 10322 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15257 10322 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15176 10322 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15095 10322 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15014 10322 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14933 10322 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14852 10322 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14771 10322 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14690 10322 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14609 10322 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14527 10322 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14445 10322 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14363 10322 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14281 10322 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14199 10322 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14117 10322 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14035 10322 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 13953 10322 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 13871 10322 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 13789 10322 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 13707 10322 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 13625 10322 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 4432 10290 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 4346 10290 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 4260 10290 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 4174 10290 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 4088 10290 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 4002 10290 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 3916 10290 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 3830 10290 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 3744 10290 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 3658 10290 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 3572 10290 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 16472 10242 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 16391 10242 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 16310 10242 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 16229 10242 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 16148 10242 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 16067 10242 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15986 10242 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15905 10242 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15824 10242 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15743 10242 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15662 10242 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15581 10242 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15500 10242 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15419 10242 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15338 10242 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15257 10242 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15176 10242 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15095 10242 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15014 10242 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14933 10242 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14852 10242 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14771 10242 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14690 10242 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14609 10242 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14527 10242 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14445 10242 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14363 10242 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14281 10242 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14199 10242 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14117 10242 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14035 10242 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 13953 10242 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 13871 10242 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 13789 10242 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 13707 10242 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 13625 10242 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 4432 10209 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 4346 10209 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 4260 10209 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 4174 10209 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 4088 10209 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 4002 10209 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 3916 10209 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 3830 10209 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 3744 10209 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 3658 10209 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 3572 10209 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 4432 4882 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 4346 4882 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 4260 4882 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 4174 4882 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 4088 4882 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 4002 4882 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 3916 4882 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 3830 4882 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 3744 4882 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 3658 4882 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 3572 4882 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 16460 4861 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 16379 4861 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 16298 4861 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 16217 4861 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 16136 4861 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 16055 4861 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15974 4861 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15893 4861 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15812 4861 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15731 4861 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15650 4861 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15569 4861 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15488 4861 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15407 4861 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15326 4861 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15245 4861 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15164 4861 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15083 4861 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 15002 4861 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14921 4861 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14840 4861 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14759 4861 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14678 4861 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14597 4861 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14515 4861 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14433 4861 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14351 4861 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14269 4861 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14187 4861 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14105 4861 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 14023 4861 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 13941 4861 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 13859 4861 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 13777 4861 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 13695 4861 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4797 13613 4861 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 4432 4800 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 4346 4800 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 4260 4800 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 4174 4800 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 4088 4800 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 4002 4800 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 3916 4800 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 3830 4800 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 3744 4800 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 3658 4800 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 3572 4800 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 16460 4781 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 16379 4781 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 16298 4781 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 16217 4781 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 16136 4781 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 16055 4781 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15974 4781 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15893 4781 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15812 4781 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15731 4781 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15650 4781 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15569 4781 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15488 4781 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15407 4781 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15326 4781 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15245 4781 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15164 4781 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15083 4781 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 15002 4781 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14921 4781 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14840 4781 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14759 4781 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14678 4781 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14597 4781 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14515 4781 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14433 4781 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14351 4781 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14269 4781 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14187 4781 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14105 4781 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 14023 4781 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 13941 4781 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 13859 4781 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 13777 4781 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 13695 4781 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4717 13613 4781 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 4432 4718 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 4346 4718 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 4260 4718 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 4174 4718 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 4088 4718 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 4002 4718 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 3916 4718 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 3830 4718 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 3744 4718 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 3658 4718 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 3572 4718 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 16460 4701 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 16379 4701 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 16298 4701 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 16217 4701 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 16136 4701 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 16055 4701 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15974 4701 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15893 4701 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15812 4701 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15731 4701 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15650 4701 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15569 4701 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15488 4701 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15407 4701 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15326 4701 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15245 4701 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15164 4701 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15083 4701 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 15002 4701 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14921 4701 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14840 4701 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14759 4701 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14678 4701 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14597 4701 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14515 4701 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14433 4701 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14351 4701 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14269 4701 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14187 4701 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14105 4701 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 14023 4701 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 13941 4701 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 13859 4701 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 13777 4701 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 13695 4701 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4637 13613 4701 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 4432 4636 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 4346 4636 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 4260 4636 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 4174 4636 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 4088 4636 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 4002 4636 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 3916 4636 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 3830 4636 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 3744 4636 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 3658 4636 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 3572 4636 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 16460 4621 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 16379 4621 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 16298 4621 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 16217 4621 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 16136 4621 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 16055 4621 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15974 4621 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15893 4621 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15812 4621 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15731 4621 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15650 4621 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15569 4621 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15488 4621 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15407 4621 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15326 4621 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15245 4621 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15164 4621 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15083 4621 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 15002 4621 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14921 4621 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14840 4621 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14759 4621 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14678 4621 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14597 4621 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14515 4621 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14433 4621 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14351 4621 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14269 4621 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14187 4621 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14105 4621 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 14023 4621 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 13941 4621 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 13859 4621 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 13777 4621 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 13695 4621 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4557 13613 4621 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 4432 4554 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 4346 4554 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 4260 4554 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 4174 4554 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 4088 4554 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 4002 4554 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 3916 4554 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 3830 4554 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 3744 4554 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 3658 4554 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 3572 4554 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 16792 4553 16856 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 16682 4553 16746 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 16572 4553 16636 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 16460 4541 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 16379 4541 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 16298 4541 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 16217 4541 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 16136 4541 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 16055 4541 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15974 4541 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15893 4541 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15812 4541 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15731 4541 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15650 4541 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15569 4541 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15488 4541 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15407 4541 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15326 4541 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15245 4541 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15164 4541 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15083 4541 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 15002 4541 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14921 4541 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14840 4541 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14759 4541 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14678 4541 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14597 4541 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14515 4541 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14433 4541 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14351 4541 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14269 4541 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14187 4541 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14105 4541 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 14023 4541 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 13941 4541 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 13859 4541 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 13777 4541 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 13695 4541 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4477 13613 4541 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 4432 4472 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 4346 4472 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 4260 4472 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 4174 4472 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 4088 4472 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 4002 4472 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 3916 4472 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 3830 4472 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 3744 4472 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 3658 4472 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 3572 4472 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 16460 4461 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 16379 4461 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 16298 4461 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 16217 4461 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 16136 4461 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 16055 4461 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15974 4461 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15893 4461 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15812 4461 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15731 4461 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15650 4461 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15569 4461 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15488 4461 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15407 4461 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15326 4461 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15245 4461 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15164 4461 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15083 4461 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 15002 4461 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14921 4461 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14840 4461 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14759 4461 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14678 4461 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14597 4461 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14515 4461 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14433 4461 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14351 4461 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14269 4461 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14187 4461 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14105 4461 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 14023 4461 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 13941 4461 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 13859 4461 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 13777 4461 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 13695 4461 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4397 13613 4461 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 4432 4390 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 4346 4390 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 4260 4390 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 4174 4390 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 4088 4390 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 4002 4390 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 3916 4390 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 3830 4390 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 3744 4390 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 3658 4390 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 3572 4390 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4331 16792 4395 16856 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4331 16682 4395 16746 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4331 16572 4395 16636 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 16460 4381 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 16379 4381 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 16298 4381 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 16217 4381 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 16136 4381 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 16055 4381 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15974 4381 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15893 4381 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15812 4381 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15731 4381 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15650 4381 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15569 4381 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15488 4381 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15407 4381 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15326 4381 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15245 4381 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15164 4381 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15083 4381 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 15002 4381 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14921 4381 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14840 4381 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14759 4381 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14678 4381 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14597 4381 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14515 4381 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14433 4381 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14351 4381 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14269 4381 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14187 4381 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14105 4381 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 14023 4381 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 13941 4381 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 13859 4381 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 13777 4381 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 13695 4381 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4317 13613 4381 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 4432 4309 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 4346 4309 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 4260 4309 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 4174 4309 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 4088 4309 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 4002 4309 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 3916 4309 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 3830 4309 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 3744 4309 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 3658 4309 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 3572 4309 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 16460 4301 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 16379 4301 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 16298 4301 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 16217 4301 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 16136 4301 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 16055 4301 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15974 4301 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15893 4301 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15812 4301 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15731 4301 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15650 4301 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15569 4301 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15488 4301 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15407 4301 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15326 4301 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15245 4301 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15164 4301 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15083 4301 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 15002 4301 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14921 4301 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14840 4301 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14759 4301 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14678 4301 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14597 4301 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14515 4301 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14433 4301 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14351 4301 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14269 4301 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14187 4301 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14105 4301 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 14023 4301 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 13941 4301 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 13859 4301 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 13777 4301 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 13695 4301 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4237 13613 4301 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4222 17053 4286 17117 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4222 16960 4286 17024 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4222 16867 4286 16931 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4222 16774 4286 16838 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4222 16682 4286 16746 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4222 16590 4286 16654 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 4432 4228 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 4346 4228 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 4260 4228 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 4174 4228 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 4088 4228 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 4002 4228 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 3916 4228 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 3830 4228 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 3744 4228 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 3658 4228 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 3572 4228 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 16460 4221 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 16379 4221 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 16298 4221 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 16217 4221 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 16136 4221 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 16055 4221 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15974 4221 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15893 4221 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15812 4221 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15731 4221 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15650 4221 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15569 4221 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15488 4221 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15407 4221 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15326 4221 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15245 4221 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15164 4221 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15083 4221 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 15002 4221 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14921 4221 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14840 4221 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14759 4221 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14678 4221 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14597 4221 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14515 4221 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14433 4221 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14351 4221 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14269 4221 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14187 4221 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14105 4221 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 14023 4221 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 13941 4221 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 13859 4221 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 13777 4221 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 13695 4221 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4157 13613 4221 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4126 17053 4190 17117 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4126 16960 4190 17024 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4126 16867 4190 16931 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4126 16774 4190 16838 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4126 16682 4190 16746 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4126 16590 4190 16654 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 4432 4147 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 4346 4147 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 4260 4147 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 4174 4147 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 4088 4147 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 4002 4147 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 3916 4147 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 3830 4147 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 3744 4147 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 3658 4147 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 3572 4147 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 16460 4141 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 16379 4141 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 16298 4141 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 16217 4141 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 16136 4141 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 16055 4141 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15974 4141 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15893 4141 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15812 4141 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15731 4141 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15650 4141 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15569 4141 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15488 4141 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15407 4141 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15326 4141 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15245 4141 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15164 4141 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15083 4141 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 15002 4141 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14921 4141 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14840 4141 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14759 4141 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14678 4141 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14597 4141 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14515 4141 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14433 4141 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14351 4141 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14269 4141 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14187 4141 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14105 4141 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 14023 4141 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 13941 4141 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 13859 4141 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 13777 4141 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 13695 4141 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4077 13613 4141 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4030 17053 4094 17117 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4030 16960 4094 17024 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4030 16867 4094 16931 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4030 16774 4094 16838 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4030 16682 4094 16746 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4030 16590 4094 16654 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 4432 4066 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 4346 4066 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 4260 4066 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 4174 4066 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 4088 4066 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 4002 4066 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 3916 4066 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 3830 4066 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 3744 4066 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 3658 4066 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 3572 4066 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 16460 4061 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 16379 4061 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 16298 4061 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 16217 4061 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 16136 4061 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 16055 4061 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15974 4061 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15893 4061 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15812 4061 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15731 4061 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15650 4061 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15569 4061 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15488 4061 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15407 4061 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15326 4061 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15245 4061 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15164 4061 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15083 4061 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 15002 4061 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14921 4061 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14840 4061 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14759 4061 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14678 4061 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14597 4061 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14515 4061 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14433 4061 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14351 4061 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14269 4061 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14187 4061 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14105 4061 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 14023 4061 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 13941 4061 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 13859 4061 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 13777 4061 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 13695 4061 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3997 13613 4061 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3948 17338 4012 17402 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3948 17250 4012 17314 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3948 17163 4012 17227 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3934 17053 3998 17117 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3934 16960 3998 17024 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3934 16867 3998 16931 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3934 16774 3998 16838 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3934 16682 3998 16746 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3934 16590 3998 16654 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 4432 3985 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 4346 3985 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 4260 3985 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 4174 3985 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 4088 3985 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 4002 3985 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 3916 3985 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 3830 3985 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 3744 3985 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 3658 3985 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 3572 3985 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 16460 3981 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 16379 3981 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 16298 3981 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 16217 3981 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 16136 3981 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 16055 3981 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15974 3981 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15893 3981 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15812 3981 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15731 3981 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15650 3981 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15569 3981 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15488 3981 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15407 3981 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15326 3981 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15245 3981 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15164 3981 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15083 3981 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 15002 3981 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14921 3981 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14840 3981 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14759 3981 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14678 3981 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14597 3981 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14515 3981 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14433 3981 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14351 3981 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14269 3981 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14187 3981 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14105 3981 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 14023 3981 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 13941 3981 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 13859 3981 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 13777 3981 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 13695 3981 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3917 13613 3981 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 4432 3904 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 4346 3904 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 4260 3904 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 4174 3904 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 4088 3904 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 4002 3904 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 3916 3904 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 3830 3904 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 3744 3904 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 3658 3904 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 3572 3904 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3838 17053 3902 17117 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3838 16960 3902 17024 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3838 16867 3902 16931 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3838 16774 3902 16838 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3838 16682 3902 16746 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3838 16590 3902 16654 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 16460 3901 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 16379 3901 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 16298 3901 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 16217 3901 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 16136 3901 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 16055 3901 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15974 3901 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15893 3901 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15812 3901 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15731 3901 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15650 3901 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15569 3901 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15488 3901 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15407 3901 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15326 3901 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15245 3901 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15164 3901 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15083 3901 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 15002 3901 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14921 3901 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14840 3901 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14759 3901 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14678 3901 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14597 3901 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14515 3901 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14433 3901 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14351 3901 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14269 3901 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14187 3901 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14105 3901 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 14023 3901 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 13941 3901 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 13859 3901 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 13777 3901 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 13695 3901 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3837 13613 3901 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3800 17338 3864 17402 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3800 17250 3864 17314 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3800 17163 3864 17227 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 4432 3823 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 4346 3823 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 4260 3823 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 4174 3823 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 4088 3823 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 4002 3823 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 3916 3823 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 3830 3823 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 3744 3823 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 3658 3823 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 3572 3823 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 16460 3821 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 16379 3821 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 16298 3821 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 16217 3821 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 16136 3821 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 16055 3821 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15974 3821 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15893 3821 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15812 3821 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15731 3821 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15650 3821 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15569 3821 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15488 3821 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15407 3821 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15326 3821 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15245 3821 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15164 3821 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15083 3821 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 15002 3821 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14921 3821 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14840 3821 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14759 3821 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14678 3821 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14597 3821 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14515 3821 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14433 3821 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14351 3821 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14269 3821 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14187 3821 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14105 3821 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 14023 3821 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 13941 3821 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 13859 3821 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 13777 3821 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 13695 3821 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3757 13613 3821 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 17563 3765 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 17482 3765 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 17401 3765 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 17320 3765 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 17239 3765 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 17159 3765 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 17079 3765 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 16999 3765 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 16919 3765 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 16839 3765 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 16759 3765 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 16679 3765 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3701 16599 3765 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 4432 3742 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 4346 3742 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 4260 3742 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 4174 3742 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 4088 3742 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 4002 3742 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 3916 3742 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 3830 3742 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 3744 3742 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 3658 3742 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 3572 3742 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 16460 3741 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 16379 3741 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 16298 3741 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 16217 3741 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 16136 3741 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 16055 3741 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15974 3741 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15893 3741 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15812 3741 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15731 3741 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15650 3741 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15569 3741 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15488 3741 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15407 3741 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15326 3741 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15245 3741 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15164 3741 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15083 3741 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 15002 3741 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14921 3741 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14840 3741 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14759 3741 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14678 3741 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14597 3741 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14515 3741 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14433 3741 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14351 3741 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14269 3741 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14187 3741 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14105 3741 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 14023 3741 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 13941 3741 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 13859 3741 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 13777 3741 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 13695 3741 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3677 13613 3741 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 17563 3683 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 17482 3683 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 17401 3683 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 17320 3683 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 17239 3683 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 17159 3683 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 17079 3683 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 16999 3683 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 16919 3683 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 16839 3683 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 16759 3683 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 16679 3683 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3619 16599 3683 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 4432 3661 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 4346 3661 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 4260 3661 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 4174 3661 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 4088 3661 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 4002 3661 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 3916 3661 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 3830 3661 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 3744 3661 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 3658 3661 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 3572 3661 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 16460 3661 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 16379 3661 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 16298 3661 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 16217 3661 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 16136 3661 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 16055 3661 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15974 3661 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15893 3661 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15812 3661 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15731 3661 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15650 3661 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15569 3661 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15488 3661 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15407 3661 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15326 3661 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15245 3661 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15164 3661 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15083 3661 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 15002 3661 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14921 3661 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14840 3661 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14759 3661 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14678 3661 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14597 3661 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14515 3661 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14433 3661 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14351 3661 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14269 3661 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14187 3661 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14105 3661 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 14023 3661 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 13941 3661 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 13859 3661 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 13777 3661 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 13695 3661 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3597 13613 3661 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 17563 3601 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 17482 3601 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 17401 3601 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 17320 3601 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 17239 3601 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 17159 3601 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 17079 3601 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 16999 3601 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 16919 3601 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 16839 3601 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 16759 3601 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 16679 3601 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3537 16599 3601 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 4432 3580 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 4346 3580 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 4260 3580 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 4174 3580 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 4088 3580 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 4002 3580 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 3916 3580 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 3830 3580 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 3744 3580 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 3658 3580 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 3572 3580 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 16460 3581 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 16379 3581 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 16298 3581 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 16217 3581 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 16136 3581 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 16055 3581 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15974 3581 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15893 3581 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15812 3581 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15731 3581 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15650 3581 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15569 3581 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15488 3581 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15407 3581 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15326 3581 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15245 3581 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15164 3581 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15083 3581 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 15002 3581 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14921 3581 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14840 3581 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14759 3581 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14678 3581 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14597 3581 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14515 3581 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14433 3581 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14351 3581 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14269 3581 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14187 3581 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14105 3581 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 14023 3581 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 13941 3581 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 13859 3581 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 13777 3581 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 13695 3581 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3517 13613 3581 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 17563 3519 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 17482 3519 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 17401 3519 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 17320 3519 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 17239 3519 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 17159 3519 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 17079 3519 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 16999 3519 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 16919 3519 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 16839 3519 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 16759 3519 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 16679 3519 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3455 16599 3519 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 4432 3499 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 4346 3499 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 4260 3499 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 4174 3499 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 4088 3499 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 4002 3499 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 3916 3499 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 3830 3499 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 3744 3499 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 3658 3499 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 3572 3499 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3440 17841 3504 17905 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3440 17757 3504 17821 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3440 17674 3504 17738 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 16460 3501 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 16379 3501 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 16298 3501 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 16217 3501 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 16136 3501 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 16055 3501 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15974 3501 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15893 3501 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15812 3501 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15731 3501 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15650 3501 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15569 3501 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15488 3501 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15407 3501 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15326 3501 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15245 3501 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15164 3501 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15083 3501 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 15002 3501 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14921 3501 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14840 3501 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14759 3501 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14678 3501 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14597 3501 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14515 3501 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14433 3501 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14351 3501 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14269 3501 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14187 3501 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14105 3501 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 14023 3501 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 13941 3501 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 13859 3501 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 13777 3501 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 13695 3501 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3437 13613 3501 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 17563 3437 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 17482 3437 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 17401 3437 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 17320 3437 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 17239 3437 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 17159 3437 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 17079 3437 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 16999 3437 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 16919 3437 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 16839 3437 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 16759 3437 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 16679 3437 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3373 16599 3437 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 4432 3418 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 4346 3418 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 4260 3418 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 4174 3418 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 4088 3418 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 4002 3418 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 3916 3418 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 3830 3418 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 3744 3418 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 3658 3418 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 3572 3418 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 16460 3421 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 16379 3421 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 16298 3421 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 16217 3421 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 16136 3421 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 16055 3421 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15974 3421 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15893 3421 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15812 3421 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15731 3421 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15650 3421 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15569 3421 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15488 3421 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15407 3421 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15326 3421 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15245 3421 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15164 3421 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15083 3421 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 15002 3421 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14921 3421 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14840 3421 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14759 3421 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14678 3421 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14597 3421 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14515 3421 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14433 3421 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14351 3421 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14269 3421 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14187 3421 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14105 3421 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 14023 3421 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 13941 3421 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 13859 3421 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 13777 3421 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 13695 3421 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3357 13613 3421 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 17563 3355 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 17482 3355 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 17401 3355 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 17320 3355 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 17239 3355 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 17159 3355 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 17079 3355 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 16999 3355 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 16919 3355 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 16839 3355 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 16759 3355 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 16679 3355 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3291 16599 3355 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 4432 3337 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 4346 3337 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 4260 3337 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 4174 3337 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 4088 3337 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 4002 3337 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 3916 3337 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 3830 3337 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 3744 3337 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 3658 3337 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 3572 3337 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3284 17841 3348 17905 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3284 17757 3348 17821 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3284 17674 3348 17738 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 16460 3341 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 16379 3341 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 16298 3341 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 16217 3341 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 16136 3341 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 16055 3341 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15974 3341 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15893 3341 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15812 3341 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15731 3341 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15650 3341 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15569 3341 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15488 3341 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15407 3341 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15326 3341 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15245 3341 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15164 3341 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15083 3341 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 15002 3341 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14921 3341 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14840 3341 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14759 3341 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14678 3341 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14597 3341 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14515 3341 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14433 3341 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14351 3341 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14269 3341 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14187 3341 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14105 3341 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 14023 3341 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 13941 3341 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 13859 3341 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 13777 3341 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 13695 3341 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3277 13613 3341 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 17563 3273 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 17482 3273 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 17401 3273 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 17320 3273 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 17239 3273 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 17159 3273 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 17079 3273 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 16999 3273 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 16919 3273 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 16839 3273 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 16759 3273 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 16679 3273 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 16599 3273 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 4432 3256 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 4346 3256 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 4260 3256 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 4174 3256 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 4088 3256 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 4002 3256 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 3916 3256 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 3830 3256 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 3744 3256 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 3658 3256 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 3572 3256 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 16460 3261 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 16379 3261 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 16298 3261 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 16217 3261 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 16136 3261 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 16055 3261 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15974 3261 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15893 3261 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15812 3261 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15731 3261 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15650 3261 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15569 3261 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15488 3261 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15407 3261 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15326 3261 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15245 3261 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15164 3261 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15083 3261 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 15002 3261 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14921 3261 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14840 3261 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14759 3261 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14678 3261 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14597 3261 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14515 3261 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14433 3261 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14351 3261 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14269 3261 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14187 3261 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14105 3261 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 14023 3261 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 13941 3261 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 13859 3261 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 13777 3261 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 13695 3261 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3197 13613 3261 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3184 18099 3248 18163 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3184 18013 3248 18077 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3184 17927 3248 17991 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3184 17841 3248 17905 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3184 17755 3248 17819 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3184 17670 3248 17734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 17563 3191 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 17482 3191 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 17401 3191 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 17320 3191 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 17239 3191 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 17159 3191 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 17079 3191 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 16999 3191 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 16919 3191 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 16839 3191 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 16759 3191 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 16679 3191 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3127 16599 3191 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 4432 3175 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 4346 3175 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 4260 3175 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 4174 3175 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 4088 3175 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 4002 3175 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 3916 3175 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 3830 3175 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 3744 3175 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 3658 3175 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 3572 3175 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 16460 3181 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 16379 3181 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 16298 3181 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 16217 3181 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 16136 3181 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 16055 3181 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15974 3181 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15893 3181 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15812 3181 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15731 3181 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15650 3181 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15569 3181 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15488 3181 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15407 3181 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15326 3181 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15245 3181 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15164 3181 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15083 3181 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 15002 3181 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14921 3181 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14840 3181 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14759 3181 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14678 3181 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14597 3181 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14515 3181 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14433 3181 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14351 3181 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14269 3181 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14187 3181 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14105 3181 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 14023 3181 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 13941 3181 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 13859 3181 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 13777 3181 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 13695 3181 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3117 13613 3181 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3102 18099 3166 18163 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3102 18013 3166 18077 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3102 17927 3166 17991 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3102 17841 3166 17905 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3102 17755 3166 17819 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3102 17670 3166 17734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 17563 3109 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 17482 3109 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 17401 3109 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 17320 3109 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 17239 3109 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 17159 3109 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 17079 3109 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 16999 3109 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 16919 3109 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 16839 3109 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 16759 3109 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 16679 3109 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3045 16599 3109 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 4432 3094 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 4346 3094 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 4260 3094 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 4174 3094 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 4088 3094 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 4002 3094 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 3916 3094 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 3830 3094 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 3744 3094 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 3658 3094 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 3572 3094 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 16460 3101 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 16379 3101 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 16298 3101 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 16217 3101 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 16136 3101 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 16055 3101 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15974 3101 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15893 3101 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15812 3101 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15731 3101 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15650 3101 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15569 3101 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15488 3101 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15407 3101 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15326 3101 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15245 3101 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15164 3101 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15083 3101 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 15002 3101 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14921 3101 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14840 3101 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14759 3101 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14678 3101 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14597 3101 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14515 3101 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14433 3101 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14351 3101 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14269 3101 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14187 3101 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14105 3101 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 14023 3101 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 13941 3101 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 13859 3101 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 13777 3101 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 13695 3101 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3037 13613 3101 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3020 18099 3084 18163 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3020 18013 3084 18077 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3020 17927 3084 17991 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3020 17841 3084 17905 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3020 17755 3084 17819 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3020 17670 3084 17734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3008 18277 3072 18341 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3008 18191 3072 18255 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 17563 3027 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 17482 3027 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 17401 3027 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 17320 3027 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 17239 3027 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 17159 3027 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 17079 3027 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 16999 3027 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 16919 3027 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 16839 3027 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 16759 3027 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 16679 3027 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2963 16599 3027 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 4432 3013 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 4346 3013 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 4260 3013 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 4174 3013 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 4088 3013 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 4002 3013 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 3916 3013 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 3830 3013 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 3744 3013 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 3658 3013 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 3572 3013 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 16460 3021 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 16379 3021 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 16298 3021 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 16217 3021 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 16136 3021 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 16055 3021 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15974 3021 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15893 3021 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15812 3021 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15731 3021 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15650 3021 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15569 3021 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15488 3021 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15407 3021 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15326 3021 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15245 3021 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15164 3021 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15083 3021 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 15002 3021 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14921 3021 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14840 3021 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14759 3021 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14678 3021 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14597 3021 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14515 3021 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14433 3021 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14351 3021 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14269 3021 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14187 3021 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14105 3021 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 14023 3021 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 13941 3021 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 13859 3021 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 13777 3021 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 13695 3021 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2957 13613 3021 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2938 18099 3002 18163 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2938 18013 3002 18077 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2938 17927 3002 17991 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2938 17841 3002 17905 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2938 17755 3002 17819 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2938 17670 3002 17734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 17563 2945 17627 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 17482 2945 17546 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 17401 2945 17465 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 17320 2945 17384 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 17239 2945 17303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 17159 2945 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 17079 2945 17143 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 16999 2945 17063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 16919 2945 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 16839 2945 16903 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 16759 2945 16823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 16679 2945 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2881 16599 2945 16663 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 4432 2932 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 4346 2932 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 4260 2932 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 4174 2932 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 4088 2932 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 4002 2932 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 3916 2932 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 3830 2932 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 3744 2932 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 3658 2932 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 3572 2932 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 16460 2941 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 16379 2941 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 16298 2941 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 16217 2941 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 16136 2941 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 16055 2941 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15974 2941 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15893 2941 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15812 2941 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15731 2941 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15650 2941 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15569 2941 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15488 2941 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15407 2941 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15326 2941 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15245 2941 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15164 2941 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15083 2941 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 15002 2941 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14921 2941 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14840 2941 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14759 2941 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14678 2941 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14597 2941 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14515 2941 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14433 2941 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14351 2941 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14269 2941 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14187 2941 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14105 2941 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 14023 2941 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 13941 2941 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 13859 2941 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 13777 2941 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 13695 2941 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2877 13613 2941 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2856 18099 2920 18163 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2856 18013 2920 18077 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2856 17927 2920 17991 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2856 17841 2920 17905 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2856 17755 2920 17819 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2856 17670 2920 17734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2852 18277 2916 18341 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2852 18191 2916 18255 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 4432 2851 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 4346 2851 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 4260 2851 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 4174 2851 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 4088 2851 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 4002 2851 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 3916 2851 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 3830 2851 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 3744 2851 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 3658 2851 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 3572 2851 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 16460 2861 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 16379 2861 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 16298 2861 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 16217 2861 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 16136 2861 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 16055 2861 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15974 2861 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15893 2861 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15812 2861 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15731 2861 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15650 2861 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15569 2861 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15488 2861 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15407 2861 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15326 2861 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15245 2861 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15164 2861 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15083 2861 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 15002 2861 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14921 2861 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14840 2861 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14759 2861 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14678 2861 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14597 2861 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14515 2861 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14433 2861 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14351 2861 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14269 2861 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14187 2861 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14105 2861 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 14023 2861 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 13941 2861 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 13859 2861 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 13777 2861 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 13695 2861 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2797 13613 2861 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 18527 2820 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 18445 2820 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 18363 2820 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 18281 2820 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 18199 2820 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 18117 2820 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 18035 2820 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17953 2820 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17871 2820 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17789 2820 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17707 2820 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17625 2820 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17543 2820 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17461 2820 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17379 2820 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17297 2820 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17215 2820 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17133 2820 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 17051 2820 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 16969 2820 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 16887 2820 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 16805 2820 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 16723 2820 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 16641 2820 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2756 16559 2820 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 4432 2770 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 4346 2770 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 4260 2770 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 4174 2770 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 4088 2770 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 4002 2770 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 3916 2770 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 3830 2770 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 3744 2770 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 3658 2770 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 3572 2770 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 16460 2781 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 16379 2781 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 16298 2781 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 16217 2781 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 16136 2781 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 16055 2781 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15974 2781 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15893 2781 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15812 2781 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15731 2781 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15650 2781 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15569 2781 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15488 2781 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15407 2781 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15326 2781 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15245 2781 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15164 2781 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15083 2781 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 15002 2781 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14921 2781 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14840 2781 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14759 2781 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14678 2781 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14597 2781 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14515 2781 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14433 2781 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14351 2781 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14269 2781 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14187 2781 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14105 2781 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 14023 2781 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 13941 2781 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 13859 2781 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 13777 2781 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 13695 2781 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2717 13613 2781 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 18527 2739 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 18445 2739 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 18363 2739 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 18281 2739 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 18199 2739 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 18117 2739 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 18035 2739 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17953 2739 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17871 2739 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17789 2739 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17707 2739 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17625 2739 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17543 2739 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17461 2739 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17379 2739 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17297 2739 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17215 2739 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17133 2739 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 17051 2739 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 16969 2739 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 16887 2739 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 16805 2739 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 16723 2739 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 16641 2739 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2675 16559 2739 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 16460 2701 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 16379 2701 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 16298 2701 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 16217 2701 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 16136 2701 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 16055 2701 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15974 2701 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15893 2701 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15812 2701 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15731 2701 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15650 2701 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15569 2701 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15488 2701 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15407 2701 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15326 2701 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15245 2701 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15164 2701 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15083 2701 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 15002 2701 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14921 2701 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14840 2701 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14759 2701 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14678 2701 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14597 2701 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14515 2701 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14433 2701 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14351 2701 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14269 2701 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14187 2701 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14105 2701 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 14023 2701 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 13941 2701 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 13859 2701 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 13777 2701 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 13695 2701 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2637 13613 2701 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 4432 2689 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 4346 2689 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 4260 2689 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 4174 2689 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 4088 2689 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 4002 2689 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 3916 2689 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 3830 2689 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 3744 2689 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 3658 2689 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 3572 2689 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 18527 2658 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 18445 2658 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 18363 2658 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 18281 2658 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 18199 2658 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 18117 2658 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 18035 2658 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17953 2658 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17871 2658 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17789 2658 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17707 2658 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17625 2658 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17543 2658 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17461 2658 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17379 2658 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17297 2658 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17215 2658 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17133 2658 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 17051 2658 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 16969 2658 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 16887 2658 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 16805 2658 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 16723 2658 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 16641 2658 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2594 16559 2658 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 16460 2621 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 16379 2621 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 16298 2621 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 16217 2621 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 16136 2621 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 16055 2621 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15974 2621 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15893 2621 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15812 2621 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15731 2621 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15650 2621 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15569 2621 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15488 2621 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15407 2621 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15326 2621 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15245 2621 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15164 2621 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15083 2621 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 15002 2621 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14921 2621 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14840 2621 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14759 2621 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14678 2621 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14597 2621 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14515 2621 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14433 2621 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14351 2621 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14269 2621 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14187 2621 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14105 2621 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 14023 2621 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 13941 2621 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 13859 2621 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 13777 2621 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 13695 2621 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2557 13613 2621 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 4432 2608 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 4346 2608 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 4260 2608 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 4174 2608 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 4088 2608 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 4002 2608 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 3916 2608 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 3830 2608 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 3744 2608 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 3658 2608 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 3572 2608 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 18527 2577 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 18445 2577 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 18363 2577 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 18281 2577 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 18199 2577 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 18117 2577 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 18035 2577 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17953 2577 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17871 2577 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17789 2577 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17707 2577 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17625 2577 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17543 2577 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17461 2577 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17379 2577 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17297 2577 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17215 2577 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17133 2577 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 17051 2577 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 16969 2577 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 16887 2577 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 16805 2577 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 16723 2577 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 16641 2577 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2513 16559 2577 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 16460 2541 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 16379 2541 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 16298 2541 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 16217 2541 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 16136 2541 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 16055 2541 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15974 2541 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15893 2541 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15812 2541 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15731 2541 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15650 2541 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15569 2541 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15488 2541 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15407 2541 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15326 2541 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15245 2541 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15164 2541 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15083 2541 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 15002 2541 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14921 2541 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14840 2541 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14759 2541 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14678 2541 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14597 2541 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14515 2541 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14433 2541 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14351 2541 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14269 2541 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14187 2541 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14105 2541 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 14023 2541 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 13941 2541 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 13859 2541 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 13777 2541 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 13695 2541 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2477 13613 2541 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 4432 2527 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 4346 2527 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 4260 2527 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 4174 2527 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 4088 2527 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 4002 2527 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 3916 2527 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 3830 2527 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 3744 2527 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 3658 2527 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 3572 2527 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 18527 2495 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 18445 2495 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 18363 2495 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 18281 2495 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 18199 2495 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 18117 2495 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 18035 2495 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17953 2495 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17871 2495 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17789 2495 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17707 2495 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17625 2495 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17543 2495 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17461 2495 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17379 2495 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17297 2495 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17215 2495 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17133 2495 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 17051 2495 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 16969 2495 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 16887 2495 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 16805 2495 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 16723 2495 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 16641 2495 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2431 16559 2495 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 16460 2461 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 16379 2461 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 16298 2461 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 16217 2461 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 16136 2461 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 16055 2461 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15974 2461 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15893 2461 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15812 2461 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15731 2461 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15650 2461 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15569 2461 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15488 2461 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15407 2461 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15326 2461 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15245 2461 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15164 2461 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15083 2461 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 15002 2461 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14921 2461 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14840 2461 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14759 2461 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14678 2461 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14597 2461 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14515 2461 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14433 2461 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14351 2461 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14269 2461 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14187 2461 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14105 2461 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 14023 2461 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 13941 2461 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 13859 2461 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 13777 2461 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 13695 2461 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2397 13613 2461 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 4432 2446 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 4346 2446 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 4260 2446 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 4174 2446 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 4088 2446 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 4002 2446 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 3916 2446 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 3830 2446 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 3744 2446 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 3658 2446 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 3572 2446 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 18527 2413 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 18445 2413 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 18363 2413 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 18281 2413 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 18199 2413 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 18117 2413 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 18035 2413 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17953 2413 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17871 2413 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17789 2413 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17707 2413 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17625 2413 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17543 2413 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17461 2413 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17379 2413 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17297 2413 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17215 2413 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17133 2413 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 17051 2413 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 16969 2413 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 16887 2413 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 16805 2413 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 16723 2413 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 16641 2413 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2349 16559 2413 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 16460 2381 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 16379 2381 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 16298 2381 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 16217 2381 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 16136 2381 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 16055 2381 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15974 2381 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15893 2381 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15812 2381 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15731 2381 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15650 2381 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15569 2381 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15488 2381 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15407 2381 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15326 2381 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15245 2381 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15164 2381 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15083 2381 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 15002 2381 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14921 2381 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14840 2381 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14759 2381 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14678 2381 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14597 2381 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14515 2381 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14433 2381 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14351 2381 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14269 2381 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14187 2381 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14105 2381 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 14023 2381 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 13941 2381 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 13859 2381 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 13777 2381 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 13695 2381 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2317 13613 2381 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 4432 2365 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 4346 2365 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 4260 2365 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 4174 2365 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 4088 2365 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 4002 2365 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 3916 2365 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 3830 2365 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 3744 2365 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 3658 2365 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 3572 2365 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 18527 2331 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 18445 2331 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 18363 2331 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 18281 2331 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 18199 2331 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 18117 2331 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 18035 2331 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17953 2331 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17871 2331 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17789 2331 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17707 2331 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17625 2331 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17543 2331 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17461 2331 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17379 2331 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17297 2331 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17215 2331 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17133 2331 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 17051 2331 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 16969 2331 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 16887 2331 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 16805 2331 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 16723 2331 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 16641 2331 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2267 16559 2331 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 16460 2301 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 16379 2301 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 16298 2301 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 16217 2301 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 16136 2301 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 16055 2301 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15974 2301 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15893 2301 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15812 2301 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15731 2301 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15650 2301 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15569 2301 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15488 2301 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15407 2301 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15326 2301 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15245 2301 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15164 2301 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15083 2301 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 15002 2301 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14921 2301 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14840 2301 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14759 2301 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14678 2301 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14597 2301 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14515 2301 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14433 2301 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14351 2301 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14269 2301 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14187 2301 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14105 2301 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 14023 2301 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 13941 2301 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 13859 2301 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 13777 2301 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 13695 2301 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2237 13613 2301 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 4432 2284 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 4346 2284 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 4260 2284 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 4174 2284 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 4088 2284 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 4002 2284 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 3916 2284 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 3830 2284 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 3744 2284 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 3658 2284 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 3572 2284 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 18527 2249 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 18445 2249 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 18363 2249 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 18281 2249 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 18199 2249 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 18117 2249 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 18035 2249 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17953 2249 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17871 2249 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17789 2249 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17707 2249 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17625 2249 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17543 2249 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17461 2249 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17379 2249 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17297 2249 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17215 2249 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17133 2249 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 17051 2249 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 16969 2249 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 16887 2249 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 16805 2249 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 16723 2249 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 16641 2249 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2185 16559 2249 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 16460 2221 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 16379 2221 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 16298 2221 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 16217 2221 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 16136 2221 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 16055 2221 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15974 2221 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15893 2221 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15812 2221 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15731 2221 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15650 2221 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15569 2221 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15488 2221 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15407 2221 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15326 2221 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15245 2221 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15164 2221 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15083 2221 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 15002 2221 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14921 2221 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14840 2221 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14759 2221 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14678 2221 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14597 2221 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14515 2221 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14433 2221 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14351 2221 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14269 2221 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14187 2221 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14105 2221 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 14023 2221 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 13941 2221 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 13859 2221 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 13777 2221 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 13695 2221 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2157 13613 2221 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 4432 2203 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 4346 2203 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 4260 2203 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 4174 2203 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 4088 2203 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 4002 2203 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 3916 2203 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 3830 2203 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 3744 2203 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 3658 2203 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 3572 2203 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 18527 2167 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 18445 2167 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 18363 2167 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 18281 2167 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 18199 2167 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 18117 2167 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 18035 2167 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17953 2167 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17871 2167 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17789 2167 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17707 2167 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17625 2167 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17543 2167 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17461 2167 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17379 2167 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17297 2167 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17215 2167 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17133 2167 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 17051 2167 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 16969 2167 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 16887 2167 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 16805 2167 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 16723 2167 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 16641 2167 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2103 16559 2167 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 16460 2141 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 16379 2141 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 16298 2141 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 16217 2141 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 16136 2141 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 16055 2141 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15974 2141 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15893 2141 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15812 2141 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15731 2141 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15650 2141 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15569 2141 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15488 2141 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15407 2141 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15326 2141 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15245 2141 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15164 2141 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15083 2141 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 15002 2141 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14921 2141 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14840 2141 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14759 2141 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14678 2141 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14597 2141 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14515 2141 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14433 2141 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14351 2141 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14269 2141 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14187 2141 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14105 2141 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 14023 2141 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 13941 2141 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 13859 2141 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 13777 2141 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 13695 2141 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2077 13613 2141 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 4432 2122 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 4346 2122 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 4260 2122 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 4174 2122 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 4088 2122 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 4002 2122 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 3916 2122 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 3830 2122 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 3744 2122 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 3658 2122 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 3572 2122 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 18527 2085 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 18445 2085 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 18363 2085 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 18281 2085 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 18199 2085 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 18117 2085 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 18035 2085 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17953 2085 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17871 2085 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17789 2085 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17707 2085 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17625 2085 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17543 2085 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17461 2085 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17379 2085 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17297 2085 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17215 2085 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17133 2085 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 17051 2085 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 16969 2085 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 16887 2085 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 16805 2085 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 16723 2085 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 16641 2085 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2021 16559 2085 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 16460 2061 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 16379 2061 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 16298 2061 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 16217 2061 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 16136 2061 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 16055 2061 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15974 2061 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15893 2061 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15812 2061 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15731 2061 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15650 2061 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15569 2061 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15488 2061 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15407 2061 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15326 2061 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15245 2061 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15164 2061 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15083 2061 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 15002 2061 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14921 2061 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14840 2061 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14759 2061 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14678 2061 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14597 2061 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14515 2061 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14433 2061 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14351 2061 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14269 2061 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14187 2061 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14105 2061 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 14023 2061 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 13941 2061 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 13859 2061 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 13777 2061 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 13695 2061 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1997 13613 2061 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 4432 2041 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 4346 2041 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 4260 2041 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 4174 2041 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 4088 2041 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 4002 2041 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 3916 2041 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 3830 2041 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 3744 2041 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 3658 2041 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 3572 2041 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 18527 2003 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 18445 2003 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 18363 2003 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 18281 2003 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 18199 2003 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 18117 2003 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 18035 2003 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17953 2003 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17871 2003 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17789 2003 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17707 2003 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17625 2003 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17543 2003 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17461 2003 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17379 2003 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17297 2003 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17215 2003 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17133 2003 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 17051 2003 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 16969 2003 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 16887 2003 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 16805 2003 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 16723 2003 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 16641 2003 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1939 16559 2003 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 16460 1981 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 16379 1981 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 16298 1981 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 16217 1981 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 16136 1981 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 16055 1981 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15974 1981 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15893 1981 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15812 1981 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15731 1981 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15650 1981 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15569 1981 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15488 1981 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15407 1981 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15326 1981 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15245 1981 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15164 1981 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15083 1981 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 15002 1981 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14921 1981 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14840 1981 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14759 1981 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14678 1981 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14597 1981 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14515 1981 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14433 1981 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14351 1981 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14269 1981 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14187 1981 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14105 1981 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 14023 1981 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 13941 1981 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 13859 1981 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 13777 1981 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 13695 1981 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1917 13613 1981 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 4432 1960 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 4346 1960 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 4260 1960 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 4174 1960 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 4088 1960 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 4002 1960 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 3916 1960 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 3830 1960 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 3744 1960 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 3658 1960 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 3572 1960 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 18527 1921 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 18445 1921 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 18363 1921 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 18281 1921 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 18199 1921 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 18117 1921 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 18035 1921 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17953 1921 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17871 1921 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17789 1921 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17707 1921 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17625 1921 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17543 1921 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17461 1921 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17379 1921 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17297 1921 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17215 1921 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17133 1921 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 17051 1921 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 16969 1921 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 16887 1921 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 16805 1921 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 16723 1921 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 16641 1921 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1857 16559 1921 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 16460 1901 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 16379 1901 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 16298 1901 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 16217 1901 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 16136 1901 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 16055 1901 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15974 1901 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15893 1901 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15812 1901 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15731 1901 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15650 1901 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15569 1901 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15488 1901 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15407 1901 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15326 1901 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15245 1901 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15164 1901 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15083 1901 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 15002 1901 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14921 1901 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14840 1901 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14759 1901 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14678 1901 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14597 1901 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14515 1901 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14433 1901 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14351 1901 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14269 1901 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14187 1901 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14105 1901 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 14023 1901 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 13941 1901 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 13859 1901 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 13777 1901 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 13695 1901 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1837 13613 1901 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 4432 1879 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 4346 1879 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 4260 1879 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 4174 1879 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 4088 1879 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 4002 1879 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 3916 1879 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 3830 1879 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 3744 1879 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 3658 1879 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 3572 1879 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 18527 1839 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 18445 1839 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 18363 1839 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 18281 1839 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 18199 1839 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 18117 1839 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 18035 1839 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17953 1839 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17871 1839 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17789 1839 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17707 1839 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17625 1839 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17543 1839 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17461 1839 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17379 1839 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17297 1839 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17215 1839 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17133 1839 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 17051 1839 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 16969 1839 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 16887 1839 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 16805 1839 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 16723 1839 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 16641 1839 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1775 16559 1839 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 16460 1821 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 16379 1821 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 16298 1821 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 16217 1821 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 16136 1821 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 16055 1821 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15974 1821 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15893 1821 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15812 1821 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15731 1821 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15650 1821 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15569 1821 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15488 1821 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15407 1821 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15326 1821 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15245 1821 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15164 1821 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15083 1821 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 15002 1821 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14921 1821 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14840 1821 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14759 1821 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14678 1821 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14597 1821 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14515 1821 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14433 1821 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14351 1821 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14269 1821 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14187 1821 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14105 1821 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 14023 1821 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 13941 1821 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 13859 1821 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 13777 1821 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 13695 1821 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1757 13613 1821 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 4432 1798 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 4346 1798 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 4260 1798 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 4174 1798 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 4088 1798 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 4002 1798 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 3916 1798 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 3830 1798 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 3744 1798 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 3658 1798 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 3572 1798 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 18527 1757 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 18445 1757 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 18363 1757 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 18281 1757 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 18199 1757 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 18117 1757 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 18035 1757 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17953 1757 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17871 1757 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17789 1757 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17707 1757 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17625 1757 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17543 1757 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17461 1757 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17379 1757 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17297 1757 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17215 1757 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17133 1757 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 17051 1757 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 16969 1757 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 16887 1757 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 16805 1757 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 16723 1757 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 16641 1757 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1693 16559 1757 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 16460 1741 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 16379 1741 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 16298 1741 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 16217 1741 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 16136 1741 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 16055 1741 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15974 1741 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15893 1741 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15812 1741 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15731 1741 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15650 1741 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15569 1741 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15488 1741 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15407 1741 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15326 1741 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15245 1741 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15164 1741 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15083 1741 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 15002 1741 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14921 1741 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14840 1741 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14759 1741 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14678 1741 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14597 1741 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14515 1741 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14433 1741 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14351 1741 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14269 1741 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14187 1741 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14105 1741 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 14023 1741 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 13941 1741 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 13859 1741 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 13777 1741 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 13695 1741 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 13613 1741 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 4432 1717 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 4346 1717 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 4260 1717 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 4174 1717 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 4088 1717 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 4002 1717 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 3916 1717 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 3830 1717 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 3744 1717 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 3658 1717 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 3572 1717 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 18527 1675 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 18445 1675 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 18363 1675 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 18281 1675 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 18199 1675 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 18117 1675 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 18035 1675 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17953 1675 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17871 1675 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17789 1675 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17707 1675 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17625 1675 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17543 1675 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17461 1675 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17379 1675 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17297 1675 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17215 1675 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17133 1675 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 17051 1675 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 16969 1675 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 16887 1675 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 16805 1675 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 16723 1675 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 16641 1675 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1611 16559 1675 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 16460 1661 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 16379 1661 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 16298 1661 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 16217 1661 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 16136 1661 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 16055 1661 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15974 1661 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15893 1661 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15812 1661 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15731 1661 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15650 1661 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15569 1661 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15488 1661 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15407 1661 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15326 1661 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15245 1661 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15164 1661 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15083 1661 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 15002 1661 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14921 1661 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14840 1661 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14759 1661 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14678 1661 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14597 1661 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14515 1661 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14433 1661 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14351 1661 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14269 1661 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14187 1661 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14105 1661 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 14023 1661 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 13941 1661 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 13859 1661 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 13777 1661 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 13695 1661 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1597 13613 1661 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 4432 1636 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 4346 1636 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 4260 1636 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 4174 1636 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 4088 1636 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 4002 1636 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 3916 1636 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 3830 1636 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 3744 1636 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 3658 1636 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 3572 1636 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 18527 1593 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 18445 1593 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 18363 1593 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 18281 1593 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 18199 1593 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 18117 1593 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 18035 1593 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17953 1593 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17871 1593 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17789 1593 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17707 1593 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17625 1593 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17543 1593 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17461 1593 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17379 1593 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17297 1593 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17215 1593 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17133 1593 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 17051 1593 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 16969 1593 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 16887 1593 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 16805 1593 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 16723 1593 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 16641 1593 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 16559 1593 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 16460 1581 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 16379 1581 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 16298 1581 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 16217 1581 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 16136 1581 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 16055 1581 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15974 1581 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15893 1581 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15812 1581 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15731 1581 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15650 1581 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15569 1581 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15488 1581 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15407 1581 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15326 1581 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15245 1581 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15164 1581 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15083 1581 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 15002 1581 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14921 1581 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14840 1581 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14759 1581 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14678 1581 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14597 1581 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14515 1581 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14433 1581 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14351 1581 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14269 1581 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14187 1581 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14105 1581 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 14023 1581 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 13941 1581 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 13859 1581 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 13777 1581 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 13695 1581 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1517 13613 1581 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 4432 1555 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 4346 1555 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 4260 1555 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 4174 1555 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 4088 1555 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 4002 1555 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 3916 1555 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 3830 1555 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 3744 1555 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 3658 1555 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 3572 1555 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 18527 1511 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 18445 1511 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 18363 1511 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 18281 1511 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 18199 1511 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 18117 1511 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 18035 1511 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17953 1511 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17871 1511 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17789 1511 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17707 1511 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17625 1511 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17543 1511 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17461 1511 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17379 1511 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17297 1511 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17215 1511 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17133 1511 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 17051 1511 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 16969 1511 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 16887 1511 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 16805 1511 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 16723 1511 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 16641 1511 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1447 16559 1511 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 16460 1501 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 16379 1501 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 16298 1501 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 16217 1501 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 16136 1501 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 16055 1501 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15974 1501 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15893 1501 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15812 1501 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15731 1501 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15650 1501 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15569 1501 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15488 1501 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15407 1501 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15326 1501 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15245 1501 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15164 1501 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15083 1501 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 15002 1501 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14921 1501 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14840 1501 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14759 1501 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14678 1501 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14597 1501 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14515 1501 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14433 1501 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14351 1501 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14269 1501 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14187 1501 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14105 1501 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 14023 1501 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 13941 1501 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 13859 1501 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 13777 1501 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 13695 1501 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1437 13613 1501 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 4432 1474 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 4346 1474 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 4260 1474 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 4174 1474 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 4088 1474 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 4002 1474 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 3916 1474 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 3830 1474 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 3744 1474 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 3658 1474 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 3572 1474 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 18527 1429 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 18445 1429 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 18363 1429 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 18281 1429 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 18199 1429 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 18117 1429 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 18035 1429 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17953 1429 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17871 1429 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17789 1429 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17707 1429 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17625 1429 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17543 1429 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17461 1429 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17379 1429 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17297 1429 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17215 1429 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17133 1429 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 17051 1429 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 16969 1429 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 16887 1429 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 16805 1429 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 16723 1429 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 16641 1429 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1365 16559 1429 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 16460 1421 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 16379 1421 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 16298 1421 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 16217 1421 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 16136 1421 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 16055 1421 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15974 1421 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15893 1421 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15812 1421 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15731 1421 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15650 1421 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15569 1421 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15488 1421 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15407 1421 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15326 1421 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15245 1421 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15164 1421 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15083 1421 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 15002 1421 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14921 1421 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14840 1421 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14759 1421 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14678 1421 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14597 1421 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14515 1421 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14433 1421 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14351 1421 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14269 1421 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14187 1421 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14105 1421 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 14023 1421 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 13941 1421 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 13859 1421 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 13777 1421 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 13695 1421 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1357 13613 1421 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 4432 1393 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 4346 1393 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 4260 1393 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 4174 1393 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 4088 1393 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 4002 1393 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 3916 1393 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 3830 1393 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 3744 1393 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 3658 1393 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 3572 1393 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 18527 1347 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 18445 1347 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 18363 1347 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 18281 1347 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 18199 1347 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 18117 1347 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 18035 1347 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17953 1347 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17871 1347 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17789 1347 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17707 1347 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17625 1347 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17543 1347 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17461 1347 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17379 1347 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17297 1347 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17215 1347 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17133 1347 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 17051 1347 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 16969 1347 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 16887 1347 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 16805 1347 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 16723 1347 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 16641 1347 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1283 16559 1347 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 16460 1341 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 16379 1341 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 16298 1341 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 16217 1341 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 16136 1341 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 16055 1341 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15974 1341 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15893 1341 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15812 1341 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15731 1341 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15650 1341 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15569 1341 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15488 1341 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15407 1341 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15326 1341 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15245 1341 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15164 1341 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15083 1341 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 15002 1341 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14921 1341 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14840 1341 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14759 1341 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14678 1341 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14597 1341 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14515 1341 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14433 1341 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14351 1341 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14269 1341 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14187 1341 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14105 1341 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 14023 1341 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 13941 1341 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 13859 1341 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 13777 1341 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 13695 1341 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1277 13613 1341 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 4432 1312 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 4346 1312 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 4260 1312 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 4174 1312 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 4088 1312 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 4002 1312 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 3916 1312 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 3830 1312 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 3744 1312 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 3658 1312 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 3572 1312 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 18527 1265 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 18445 1265 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 18363 1265 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 18281 1265 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 18199 1265 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 18117 1265 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 18035 1265 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17953 1265 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17871 1265 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17789 1265 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17707 1265 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17625 1265 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17543 1265 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17461 1265 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17379 1265 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17297 1265 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17215 1265 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17133 1265 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 17051 1265 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 16969 1265 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 16887 1265 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 16805 1265 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 16723 1265 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 16641 1265 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1201 16559 1265 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 16460 1261 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 16379 1261 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 16298 1261 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 16217 1261 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 16136 1261 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 16055 1261 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15974 1261 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15893 1261 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15812 1261 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15731 1261 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15650 1261 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15569 1261 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15488 1261 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15407 1261 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15326 1261 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15245 1261 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15164 1261 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15083 1261 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 15002 1261 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14921 1261 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14840 1261 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14759 1261 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14678 1261 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14597 1261 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14515 1261 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14433 1261 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14351 1261 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14269 1261 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14187 1261 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14105 1261 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 14023 1261 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 13941 1261 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 13859 1261 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 13777 1261 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 13695 1261 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1197 13613 1261 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 4432 1231 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 4346 1231 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 4260 1231 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 4174 1231 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 4088 1231 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 4002 1231 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 3916 1231 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 3830 1231 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 3744 1231 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 3658 1231 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 3572 1231 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 18527 1183 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 18445 1183 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 18363 1183 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 18281 1183 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 18199 1183 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 18117 1183 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 18035 1183 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17953 1183 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17871 1183 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17789 1183 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17707 1183 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17625 1183 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17543 1183 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17461 1183 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17379 1183 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17297 1183 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17215 1183 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17133 1183 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 17051 1183 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 16969 1183 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 16887 1183 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 16805 1183 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 16723 1183 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 16641 1183 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1119 16559 1183 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 16460 1181 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 16379 1181 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 16298 1181 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 16217 1181 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 16136 1181 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 16055 1181 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15974 1181 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15893 1181 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15812 1181 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15731 1181 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15650 1181 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15569 1181 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15488 1181 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15407 1181 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15326 1181 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15245 1181 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15164 1181 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15083 1181 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 15002 1181 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14921 1181 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14840 1181 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14759 1181 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14678 1181 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14597 1181 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14515 1181 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14433 1181 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14351 1181 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14269 1181 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14187 1181 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14105 1181 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 14023 1181 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 13941 1181 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 13859 1181 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 13777 1181 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 13695 1181 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1117 13613 1181 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 4432 1150 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 4346 1150 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 4260 1150 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 4174 1150 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 4088 1150 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 4002 1150 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 3916 1150 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 3830 1150 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 3744 1150 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 3658 1150 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 3572 1150 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 18527 1101 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 18445 1101 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 18363 1101 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 18281 1101 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 18199 1101 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 18117 1101 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 18035 1101 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17953 1101 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17871 1101 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17789 1101 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17707 1101 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17625 1101 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17543 1101 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17461 1101 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17379 1101 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17297 1101 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17215 1101 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17133 1101 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 17051 1101 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16969 1101 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16887 1101 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16805 1101 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16723 1101 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16641 1101 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16559 1101 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16460 1101 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16379 1101 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16298 1101 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16217 1101 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16136 1101 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 16055 1101 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15974 1101 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15893 1101 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15812 1101 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15731 1101 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15650 1101 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15569 1101 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15488 1101 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15407 1101 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15326 1101 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15245 1101 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15164 1101 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15083 1101 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 15002 1101 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14921 1101 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14840 1101 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14759 1101 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14678 1101 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14597 1101 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14515 1101 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14433 1101 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14351 1101 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14269 1101 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14187 1101 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14105 1101 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 14023 1101 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 13941 1101 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 13859 1101 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 13777 1101 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 13695 1101 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1037 13613 1101 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 4432 1069 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 4346 1069 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 4260 1069 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 4174 1069 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 4088 1069 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 4002 1069 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 3916 1069 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 3830 1069 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 3744 1069 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 3658 1069 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 3572 1069 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 16460 1021 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 16379 1021 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 16298 1021 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 16217 1021 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 16136 1021 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 16055 1021 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15974 1021 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15893 1021 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15812 1021 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15731 1021 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15650 1021 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15569 1021 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15488 1021 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15407 1021 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15326 1021 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15245 1021 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15164 1021 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15083 1021 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 15002 1021 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14921 1021 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14840 1021 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14759 1021 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14678 1021 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14597 1021 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14515 1021 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14433 1021 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14351 1021 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14269 1021 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14187 1021 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14105 1021 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 14023 1021 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 13941 1021 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 13859 1021 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 13777 1021 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 13695 1021 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 957 13613 1021 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 18527 1019 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 18445 1019 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 18363 1019 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 18281 1019 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 18199 1019 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 18117 1019 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 18035 1019 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17953 1019 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17871 1019 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17789 1019 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17707 1019 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17625 1019 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17543 1019 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17461 1019 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17379 1019 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17297 1019 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17215 1019 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17133 1019 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 17051 1019 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 16969 1019 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 16887 1019 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 16805 1019 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 16723 1019 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 16641 1019 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 955 16559 1019 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 4432 988 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 4346 988 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 4260 988 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 4174 988 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 4088 988 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 4002 988 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 3916 988 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 3830 988 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 3744 988 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 3658 988 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 3572 988 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 16460 941 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 16379 941 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 16298 941 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 16217 941 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 16136 941 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 16055 941 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15974 941 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15893 941 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15812 941 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15731 941 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15650 941 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15569 941 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15488 941 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15407 941 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15326 941 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15245 941 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15164 941 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15083 941 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 15002 941 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14921 941 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14840 941 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14759 941 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14678 941 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14597 941 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14515 941 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14433 941 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14351 941 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14269 941 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14187 941 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14105 941 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 14023 941 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 13941 941 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 13859 941 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 13777 941 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 13695 941 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 877 13613 941 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 18527 937 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 18445 937 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 18363 937 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 18281 937 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 18199 937 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 18117 937 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 18035 937 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17953 937 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17871 937 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17789 937 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17707 937 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17625 937 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17543 937 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17461 937 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17379 937 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17297 937 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17215 937 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17133 937 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 17051 937 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 16969 937 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 16887 937 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 16805 937 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 16723 937 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 16641 937 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 873 16559 937 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 4432 907 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 4346 907 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 4260 907 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 4174 907 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 4088 907 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 4002 907 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 3916 907 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 3830 907 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 3744 907 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 3658 907 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 3572 907 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 16460 861 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 16379 861 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 16298 861 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 16217 861 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 16136 861 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 16055 861 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15974 861 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15893 861 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15812 861 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15731 861 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15650 861 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15569 861 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15488 861 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15407 861 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15326 861 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15245 861 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15164 861 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15083 861 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 15002 861 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14921 861 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14840 861 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14759 861 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14678 861 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14597 861 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14515 861 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14433 861 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14351 861 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14269 861 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14187 861 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14105 861 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 14023 861 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 13941 861 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 13859 861 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 13777 861 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 13695 861 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 797 13613 861 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 18527 855 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 18445 855 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 18363 855 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 18281 855 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 18199 855 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 18117 855 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 18035 855 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17953 855 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17871 855 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17789 855 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17707 855 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17625 855 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17543 855 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17461 855 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17379 855 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17297 855 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17215 855 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17133 855 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 17051 855 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 16969 855 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 16887 855 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 16805 855 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 16723 855 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 16641 855 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 791 16559 855 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 4432 826 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 4346 826 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 4260 826 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 4174 826 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 4088 826 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 4002 826 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 3916 826 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 3830 826 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 3744 826 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 3658 826 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 3572 826 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 16460 781 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 16379 781 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 16298 781 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 16217 781 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 16136 781 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 16055 781 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15974 781 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15893 781 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15812 781 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15731 781 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15650 781 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15569 781 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15488 781 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15407 781 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15326 781 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15245 781 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15164 781 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15083 781 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 15002 781 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14921 781 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14840 781 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14759 781 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14678 781 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14597 781 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14515 781 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14433 781 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14351 781 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14269 781 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14187 781 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14105 781 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 14023 781 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 13941 781 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 13859 781 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 13777 781 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 13695 781 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 717 13613 781 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 18527 773 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 18445 773 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 18363 773 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 18281 773 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 18199 773 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 18117 773 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 18035 773 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17953 773 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17871 773 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17789 773 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17707 773 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17625 773 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17543 773 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17461 773 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17379 773 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17297 773 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17215 773 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17133 773 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 17051 773 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 16969 773 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 16887 773 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 16805 773 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 16723 773 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 16641 773 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 709 16559 773 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 4432 745 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 4346 745 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 4260 745 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 4174 745 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 4088 745 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 4002 745 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 3916 745 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 3830 745 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 3744 745 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 3658 745 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 3572 745 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 16460 701 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 16379 701 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 16298 701 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 16217 701 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 16136 701 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 16055 701 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15974 701 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15893 701 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15812 701 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15731 701 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15650 701 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15569 701 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15488 701 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15407 701 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15326 701 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15245 701 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15164 701 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15083 701 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 15002 701 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14921 701 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14840 701 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14759 701 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14678 701 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14597 701 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14515 701 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14433 701 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14351 701 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14269 701 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14187 701 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14105 701 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 14023 701 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 13941 701 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 13859 701 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 13777 701 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 13695 701 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 637 13613 701 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 18527 691 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 18445 691 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 18363 691 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 18281 691 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 18199 691 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 18117 691 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 18035 691 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17953 691 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17871 691 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17789 691 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17707 691 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17625 691 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17543 691 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17461 691 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17379 691 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17297 691 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17215 691 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17133 691 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 17051 691 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 16969 691 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 16887 691 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 16805 691 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 16723 691 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 16641 691 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 627 16559 691 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 4432 664 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 4346 664 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 4260 664 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 4174 664 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 4088 664 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 4002 664 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 3916 664 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 3830 664 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 3744 664 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 3658 664 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 3572 664 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 16460 621 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 16379 621 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 16298 621 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 16217 621 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 16136 621 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 16055 621 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15974 621 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15893 621 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15812 621 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15731 621 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15650 621 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15569 621 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15488 621 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15407 621 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15326 621 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15245 621 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15164 621 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15083 621 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 15002 621 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14921 621 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14840 621 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14759 621 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14678 621 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14597 621 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14515 621 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14433 621 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14351 621 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14269 621 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14187 621 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14105 621 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 14023 621 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 13941 621 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 13859 621 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 13777 621 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 13695 621 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 13613 621 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 18527 609 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 18445 609 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 18363 609 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 18281 609 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 18199 609 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 18117 609 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 18035 609 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17953 609 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17871 609 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17789 609 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17707 609 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17625 609 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17543 609 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17461 609 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17379 609 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17297 609 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17215 609 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17133 609 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 17051 609 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 16969 609 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 16887 609 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 16805 609 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 16723 609 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 16641 609 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 545 16559 609 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 4432 583 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 4346 583 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 4260 583 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 4174 583 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 4088 583 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 4002 583 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 3916 583 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 3830 583 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 3744 583 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 3658 583 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 3572 583 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 16460 541 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 16379 541 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 16298 541 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 16217 541 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 16136 541 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 16055 541 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15974 541 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15893 541 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15812 541 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15731 541 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15650 541 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15569 541 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15488 541 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15407 541 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15326 541 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15245 541 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15164 541 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15083 541 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 15002 541 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14921 541 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14840 541 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14759 541 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14678 541 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14597 541 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14515 541 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14433 541 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14351 541 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14269 541 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14187 541 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14105 541 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 14023 541 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 13941 541 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 13859 541 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 13777 541 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 13695 541 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 477 13613 541 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 18527 527 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 18445 527 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 18363 527 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 18281 527 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 18199 527 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 18117 527 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 18035 527 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17953 527 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17871 527 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17789 527 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17707 527 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17625 527 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17543 527 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17461 527 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17379 527 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17297 527 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17215 527 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17133 527 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 17051 527 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 16969 527 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 16887 527 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 16805 527 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 16723 527 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 16641 527 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 463 16559 527 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 4432 502 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 4346 502 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 4260 502 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 4174 502 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 4088 502 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 4002 502 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 3916 502 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 3830 502 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 3744 502 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 3658 502 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 3572 502 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 16460 461 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 16379 461 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 16298 461 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 16217 461 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 16136 461 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 16055 461 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15974 461 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15893 461 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15812 461 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15731 461 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15650 461 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15569 461 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15488 461 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15407 461 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15326 461 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15245 461 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15164 461 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15083 461 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 15002 461 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14921 461 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14840 461 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14759 461 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14678 461 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14597 461 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14515 461 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14433 461 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14351 461 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14269 461 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14187 461 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14105 461 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 14023 461 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 13941 461 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 13859 461 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 13777 461 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 13695 461 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 397 13613 461 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 18527 445 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 18445 445 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 18363 445 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 18281 445 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 18199 445 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 18117 445 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 18035 445 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17953 445 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17871 445 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17789 445 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17707 445 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17625 445 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17543 445 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17461 445 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17379 445 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17297 445 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17215 445 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17133 445 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 17051 445 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 16969 445 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 16887 445 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 16805 445 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 16723 445 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 16641 445 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 16559 445 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 4432 421 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 4346 421 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 4260 421 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 4174 421 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 4088 421 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 4002 421 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 3916 421 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 3830 421 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 3744 421 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 3658 421 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 3572 421 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 16460 381 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 16379 381 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 16298 381 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 16217 381 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 16136 381 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 16055 381 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15974 381 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15893 381 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15812 381 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15731 381 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15650 381 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15569 381 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15488 381 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15407 381 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15326 381 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15245 381 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15164 381 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15083 381 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 15002 381 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14921 381 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14840 381 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14759 381 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14678 381 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14597 381 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14515 381 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14433 381 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14351 381 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14269 381 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14187 381 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14105 381 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 14023 381 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 13941 381 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 13859 381 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 13777 381 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 13695 381 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 317 13613 381 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 18527 363 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 18445 363 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 18363 363 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 18281 363 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 18199 363 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 18117 363 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 18035 363 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17953 363 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17871 363 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17789 363 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17707 363 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17625 363 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17543 363 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17461 363 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17379 363 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17297 363 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17215 363 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17133 363 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 17051 363 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 16969 363 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 16887 363 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 16805 363 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 16723 363 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 16641 363 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 299 16559 363 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 4432 340 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 4346 340 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 4260 340 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 4174 340 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 4088 340 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 4002 340 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 3916 340 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 3830 340 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 3744 340 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 3658 340 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 3572 340 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 16460 301 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 16379 301 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 16298 301 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 16217 301 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 16136 301 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 16055 301 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15974 301 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15893 301 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15812 301 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15731 301 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15650 301 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15569 301 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15488 301 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15407 301 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15326 301 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15245 301 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15164 301 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15083 301 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 15002 301 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14921 301 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14840 301 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14759 301 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14678 301 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14597 301 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14515 301 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14433 301 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14351 301 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14269 301 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14187 301 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14105 301 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 14023 301 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 13941 301 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 13859 301 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 13777 301 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 13695 301 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 237 13613 301 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 18527 281 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 18445 281 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 18363 281 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 18281 281 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 18199 281 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 18117 281 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 18035 281 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17953 281 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17871 281 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17789 281 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17707 281 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17625 281 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17543 281 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17461 281 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17379 281 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17297 281 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17215 281 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17133 281 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 17051 281 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 16969 281 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 16887 281 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 16805 281 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 16723 281 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 16641 281 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 217 16559 281 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 4432 259 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 4346 259 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 4260 259 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 4174 259 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 4088 259 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 4002 259 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 3916 259 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 3830 259 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 3744 259 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 3658 259 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 3572 259 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 16460 221 16524 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 16379 221 16443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 16298 221 16362 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 16217 221 16281 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 16136 221 16200 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 16055 221 16119 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15974 221 16038 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15893 221 15957 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15812 221 15876 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15731 221 15795 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15650 221 15714 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15569 221 15633 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15488 221 15552 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15407 221 15471 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15326 221 15390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15245 221 15309 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15164 221 15228 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15083 221 15147 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 15002 221 15066 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14921 221 14985 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14840 221 14904 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14759 221 14823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14678 221 14742 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14597 221 14661 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14515 221 14579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14433 221 14497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14351 221 14415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14269 221 14333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14187 221 14251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14105 221 14169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 14023 221 14087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 13941 221 14005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 13859 221 13923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 13777 221 13841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 13695 221 13759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 157 13613 221 13677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 18527 199 18591 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 18445 199 18509 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 18363 199 18427 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 18281 199 18345 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 18199 199 18263 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 18117 199 18181 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 18035 199 18099 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17953 199 18017 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17871 199 17935 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17789 199 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17707 199 17771 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17625 199 17689 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17543 199 17607 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17461 199 17525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17379 199 17443 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17297 199 17361 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17215 199 17279 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17133 199 17197 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 17051 199 17115 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 16969 199 17033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 16887 199 16951 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 16805 199 16869 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 16723 199 16787 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 16641 199 16705 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 135 16559 199 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 4432 178 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 4346 178 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 4260 178 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 4174 178 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 4088 178 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 4002 178 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 3916 178 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 3830 178 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 3744 178 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 3658 178 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 3572 178 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 120 3558 4900 4486 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10151 3558 14931 4486 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12211 18573 14932 18592 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12192 18543 14932 18573 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12162 18513 14932 18543 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12132 18483 14932 18513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12102 18453 14932 18483 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12072 18423 14932 18453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 18393 14932 18423 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12012 18363 14932 18393 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11982 18333 14932 18363 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11952 18303 14932 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11922 18273 14932 18303 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11892 18243 14932 18273 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11862 18213 14932 18243 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11832 18183 14932 18213 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 18153 14932 18183 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11772 18123 14932 18153 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11742 18093 14932 18123 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11712 18063 14932 18093 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11682 18033 14932 18063 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11652 18003 14932 18033 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11622 17973 14932 18003 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11592 17943 14932 17973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 17913 14932 17943 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11532 17883 14932 17913 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11502 17853 14932 17883 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11472 17823 14932 17853 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11442 17793 14932 17823 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11412 17763 14932 17793 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11382 17733 14932 17763 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11352 17703 14932 17733 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 17673 14932 17703 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11292 17643 14932 17673 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11262 17613 14932 17643 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11232 17583 14932 17613 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11202 17553 14932 17583 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11172 17523 14932 17553 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11142 17493 14932 17523 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11112 17463 14932 17493 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 17433 14932 17463 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11052 17403 14932 17433 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11022 17373 14932 17403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10992 17343 14932 17373 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10962 17313 14932 17343 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10932 17283 14932 17313 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10902 17253 14932 17283 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10872 17223 14932 17253 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 17193 14932 17223 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10812 17163 14932 17193 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10782 17133 14932 17163 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10752 17103 14932 17133 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10722 17073 14932 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10692 17043 14932 17073 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10662 17013 14932 17043 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10632 16983 14932 17013 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 16953 14932 16983 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10572 16923 14932 16953 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10542 16893 14932 16923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10512 16863 14932 16893 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10482 16833 14932 16863 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10452 16803 14932 16833 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10422 16773 14932 16803 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10392 16743 14932 16773 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 16713 14932 16743 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10332 16683 14932 16713 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10302 16653 14932 16683 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10272 16623 14932 16653 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10242 16593 14932 16623 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10212 16563 14932 16593 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10182 16533 14932 16563 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10152 13607 14932 16533 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 0 3557 4895 4487 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 0 18592 254 18600 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 0 16558 2821 18592 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 0 16525 254 16558 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 0 13612 4900 16525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 0 13607 254 13612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2851 18190 3073 18342 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2854 17669 3250 18164 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 2875 16598 3771 17628 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3283 17673 3505 17906 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3799 17162 4013 17403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 3834 16589 4290 17118 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 4330 16571 4554 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14746 18593 15000 18600 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14746 16525 15000 16557 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 14746 13607 15000 13612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 12230 16557 15000 18593 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10151 13612 15000 16525 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10156 3557 15000 4487 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10497 16571 10721 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 10761 16589 11217 17118 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11038 17162 11252 17403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11280 16598 12176 17628 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11546 17673 11768 17906 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11801 17669 12197 18164 6 VDDIO
port 7 nsew power bidirectional
rlabel metal4 s 11978 18190 12200 18342 6 VDDIO
port 7 nsew power bidirectional
rlabel metal5 s 0 3577 254 4467 6 VDDIO
port 7 nsew power bidirectional
rlabel metal5 s 0 13607 254 18597 6 VDDIO
port 7 nsew power bidirectional
rlabel metal5 s 14746 3577 15000 4467 6 VDDIO
port 7 nsew power bidirectional
rlabel metal5 s 14746 13607 15000 18597 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 4432 14913 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 4346 14913 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 4260 14913 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 4174 14913 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 4088 14913 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 4002 14913 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 3916 14913 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 3830 14913 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 3744 14913 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 3658 14913 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14873 3572 14913 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 18539 14904 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 18457 14904 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 18375 14904 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 18293 14904 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 18211 14904 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 18129 14904 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 18047 14904 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 17965 14904 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 17883 14904 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 17801 14904 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 17719 14904 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 17637 14904 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 17555 14904 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 17473 14904 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 17391 14904 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 17309 14904 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 17227 14904 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 17145 14904 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 17063 14904 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 16981 14904 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 16899 14904 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 16817 14904 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 16735 14904 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 16653 14904 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14864 16571 14904 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 16472 14882 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 16391 14882 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 16310 14882 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 16229 14882 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 16148 14882 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 16067 14882 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15986 14882 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15905 14882 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15824 14882 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15743 14882 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15662 14882 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15581 14882 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15500 14882 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15419 14882 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15338 14882 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15257 14882 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15176 14882 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15095 14882 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 15014 14882 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14933 14882 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14852 14882 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14771 14882 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14690 14882 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14609 14882 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14527 14882 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14445 14882 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14363 14882 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14281 14882 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14199 14882 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14117 14882 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 14035 14882 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 13953 14882 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 13871 14882 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 13789 14882 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 13707 14882 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14842 13625 14882 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 4432 14831 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 4346 14831 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 4260 14831 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 4174 14831 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 4088 14831 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 4002 14831 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 3916 14831 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 3830 14831 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 3744 14831 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 3658 14831 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14791 3572 14831 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 18539 14822 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 18457 14822 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 18375 14822 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 18293 14822 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 18211 14822 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 18129 14822 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 18047 14822 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 17965 14822 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 17883 14822 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 17801 14822 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 17719 14822 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 17637 14822 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 17555 14822 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 17473 14822 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 17391 14822 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 17309 14822 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 17227 14822 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 17145 14822 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 17063 14822 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 16981 14822 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 16899 14822 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 16817 14822 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 16735 14822 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 16653 14822 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14782 16571 14822 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 16472 14802 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 16391 14802 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 16310 14802 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 16229 14802 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 16148 14802 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 16067 14802 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15986 14802 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15905 14802 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15824 14802 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15743 14802 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15662 14802 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15581 14802 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15500 14802 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15419 14802 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15338 14802 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15257 14802 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15176 14802 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15095 14802 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 15014 14802 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14933 14802 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14852 14802 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14771 14802 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14690 14802 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14609 14802 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14527 14802 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14445 14802 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14363 14802 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14281 14802 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14199 14802 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14117 14802 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 14035 14802 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 13953 14802 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 13871 14802 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 13789 14802 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 13707 14802 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14762 13625 14802 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 4432 14749 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 4346 14749 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 4260 14749 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 4174 14749 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 4088 14749 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 4002 14749 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 3916 14749 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 3830 14749 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 3744 14749 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 3658 14749 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14709 3572 14749 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 18539 14740 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 18457 14740 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 18375 14740 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 18293 14740 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 18211 14740 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 18129 14740 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 18047 14740 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 17965 14740 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 17883 14740 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 17801 14740 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 17719 14740 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 17637 14740 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 17555 14740 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 17473 14740 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 17391 14740 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 17309 14740 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 17227 14740 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 17145 14740 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 17063 14740 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 16981 14740 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 16899 14740 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 16817 14740 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 16735 14740 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 16653 14740 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14700 16571 14740 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 16472 14722 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 16391 14722 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 16310 14722 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 16229 14722 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 16148 14722 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 16067 14722 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15986 14722 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15905 14722 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15824 14722 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15743 14722 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15662 14722 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15581 14722 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15500 14722 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15419 14722 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15338 14722 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15257 14722 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15176 14722 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15095 14722 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 15014 14722 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14933 14722 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14852 14722 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14771 14722 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14690 14722 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14609 14722 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14527 14722 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14445 14722 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14363 14722 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14281 14722 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14199 14722 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14117 14722 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 14035 14722 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 13953 14722 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 13871 14722 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 13789 14722 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 13707 14722 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14682 13625 14722 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 4432 14667 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 4346 14667 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 4260 14667 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 4174 14667 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 4088 14667 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 4002 14667 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 3916 14667 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 3830 14667 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 3744 14667 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 3658 14667 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14627 3572 14667 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 18539 14658 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 18457 14658 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 18375 14658 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 18293 14658 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 18211 14658 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 18129 14658 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 18047 14658 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 17965 14658 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 17883 14658 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 17801 14658 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 17719 14658 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 17637 14658 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 17555 14658 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 17473 14658 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 17391 14658 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 17309 14658 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 17227 14658 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 17145 14658 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 17063 14658 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 16981 14658 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 16899 14658 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 16817 14658 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 16735 14658 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 16653 14658 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14618 16571 14658 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 16472 14642 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 16391 14642 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 16310 14642 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 16229 14642 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 16148 14642 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 16067 14642 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15986 14642 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15905 14642 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15824 14642 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15743 14642 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15662 14642 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15581 14642 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15500 14642 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15419 14642 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15338 14642 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15257 14642 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15176 14642 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15095 14642 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 15014 14642 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14933 14642 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14852 14642 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14771 14642 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14690 14642 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14609 14642 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14527 14642 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14445 14642 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14363 14642 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14281 14642 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14199 14642 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14117 14642 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 14035 14642 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 13953 14642 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 13871 14642 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 13789 14642 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 13707 14642 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14602 13625 14642 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 4432 14585 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 4346 14585 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 4260 14585 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 4174 14585 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 4088 14585 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 4002 14585 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 3916 14585 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 3830 14585 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 3744 14585 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 3658 14585 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14545 3572 14585 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 18539 14576 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 18457 14576 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 18375 14576 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 18293 14576 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 18211 14576 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 18129 14576 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 18047 14576 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 17965 14576 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 17883 14576 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 17801 14576 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 17719 14576 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 17637 14576 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 17555 14576 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 17473 14576 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 17391 14576 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 17309 14576 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 17227 14576 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 17145 14576 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 17063 14576 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 16981 14576 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 16899 14576 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 16817 14576 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 16735 14576 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 16653 14576 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14536 16571 14576 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 16472 14562 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 16391 14562 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 16310 14562 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 16229 14562 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 16148 14562 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 16067 14562 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15986 14562 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15905 14562 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15824 14562 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15743 14562 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15662 14562 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15581 14562 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15500 14562 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15419 14562 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15338 14562 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15257 14562 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15176 14562 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15095 14562 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 15014 14562 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14933 14562 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14852 14562 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14771 14562 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14690 14562 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14609 14562 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14527 14562 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14445 14562 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14363 14562 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14281 14562 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14199 14562 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14117 14562 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 14035 14562 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 13953 14562 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 13871 14562 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 13789 14562 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 13707 14562 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14522 13625 14562 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 4432 14503 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 4346 14503 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 4260 14503 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 4174 14503 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 4088 14503 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 4002 14503 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 3916 14503 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 3830 14503 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 3744 14503 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 3658 14503 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14463 3572 14503 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 18539 14494 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 18457 14494 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 18375 14494 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 18293 14494 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 18211 14494 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 18129 14494 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 18047 14494 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 17965 14494 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 17883 14494 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 17801 14494 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 17719 14494 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 17637 14494 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 17555 14494 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 17473 14494 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 17391 14494 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 17309 14494 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 17227 14494 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 17145 14494 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 17063 14494 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 16981 14494 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 16899 14494 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 16817 14494 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 16735 14494 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 16653 14494 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14454 16571 14494 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16472 14482 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16391 14482 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16310 14482 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16229 14482 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16148 14482 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 16067 14482 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15986 14482 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15905 14482 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15824 14482 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15743 14482 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15662 14482 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15581 14482 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15500 14482 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15419 14482 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15338 14482 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15257 14482 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15176 14482 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15095 14482 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 15014 14482 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14933 14482 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14852 14482 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14771 14482 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14690 14482 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14609 14482 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14527 14482 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14445 14482 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14363 14482 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14281 14482 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14199 14482 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14117 14482 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 14035 14482 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 13953 14482 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 13871 14482 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 13789 14482 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 13707 14482 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14442 13625 14482 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 4432 14421 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 4346 14421 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 4260 14421 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 4174 14421 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 4088 14421 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 4002 14421 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 3916 14421 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 3830 14421 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 3744 14421 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 3658 14421 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14381 3572 14421 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 18539 14412 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 18457 14412 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 18375 14412 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 18293 14412 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 18211 14412 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 18129 14412 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 18047 14412 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 17965 14412 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 17883 14412 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 17801 14412 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 17719 14412 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 17637 14412 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 17555 14412 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 17473 14412 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 17391 14412 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 17309 14412 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 17227 14412 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 17145 14412 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 17063 14412 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 16981 14412 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 16899 14412 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 16817 14412 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 16735 14412 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 16653 14412 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14372 16571 14412 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 16472 14402 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 16391 14402 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 16310 14402 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 16229 14402 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 16148 14402 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 16067 14402 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15986 14402 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15905 14402 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15824 14402 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15743 14402 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15662 14402 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15581 14402 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15500 14402 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15419 14402 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15338 14402 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15257 14402 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15176 14402 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15095 14402 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 15014 14402 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14933 14402 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14852 14402 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14771 14402 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14690 14402 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14609 14402 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14527 14402 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14445 14402 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14363 14402 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14281 14402 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14199 14402 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14117 14402 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 14035 14402 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 13953 14402 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 13871 14402 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 13789 14402 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 13707 14402 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14362 13625 14402 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 4432 14340 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 4346 14340 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 4260 14340 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 4174 14340 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 4088 14340 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 4002 14340 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 3916 14340 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 3830 14340 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 3744 14340 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 3658 14340 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14300 3572 14340 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 18539 14330 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 18457 14330 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 18375 14330 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 18293 14330 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 18211 14330 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 18129 14330 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 18047 14330 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 17965 14330 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 17883 14330 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 17801 14330 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 17719 14330 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 17637 14330 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 17555 14330 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 17473 14330 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 17391 14330 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 17309 14330 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 17227 14330 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 17145 14330 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 17063 14330 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 16981 14330 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 16899 14330 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 16817 14330 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 16735 14330 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 16653 14330 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14290 16571 14330 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 16472 14322 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 16391 14322 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 16310 14322 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 16229 14322 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 16148 14322 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 16067 14322 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15986 14322 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15905 14322 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15824 14322 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15743 14322 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15662 14322 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15581 14322 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15500 14322 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15419 14322 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15338 14322 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15257 14322 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15176 14322 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15095 14322 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 15014 14322 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14933 14322 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14852 14322 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14771 14322 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14690 14322 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14609 14322 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14527 14322 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14445 14322 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14363 14322 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14281 14322 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14199 14322 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14117 14322 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 14035 14322 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 13953 14322 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 13871 14322 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 13789 14322 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 13707 14322 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14282 13625 14322 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 4432 14259 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 4346 14259 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 4260 14259 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 4174 14259 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 4088 14259 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 4002 14259 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 3916 14259 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 3830 14259 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 3744 14259 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 3658 14259 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14219 3572 14259 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 18539 14248 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 18457 14248 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 18375 14248 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 18293 14248 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 18211 14248 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 18129 14248 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 18047 14248 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 17965 14248 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 17883 14248 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 17801 14248 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 17719 14248 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 17637 14248 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 17555 14248 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 17473 14248 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 17391 14248 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 17309 14248 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 17227 14248 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 17145 14248 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 17063 14248 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 16981 14248 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 16899 14248 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 16817 14248 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 16735 14248 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 16653 14248 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14208 16571 14248 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 16472 14242 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 16391 14242 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 16310 14242 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 16229 14242 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 16148 14242 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 16067 14242 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15986 14242 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15905 14242 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15824 14242 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15743 14242 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15662 14242 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15581 14242 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15500 14242 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15419 14242 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15338 14242 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15257 14242 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15176 14242 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15095 14242 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 15014 14242 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14933 14242 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14852 14242 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14771 14242 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14690 14242 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14609 14242 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14527 14242 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14445 14242 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14363 14242 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14281 14242 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14199 14242 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14117 14242 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 14035 14242 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 13953 14242 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 13871 14242 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 13789 14242 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 13707 14242 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14202 13625 14242 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 4432 14178 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 4346 14178 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 4260 14178 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 4174 14178 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 4088 14178 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 4002 14178 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 3916 14178 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 3830 14178 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 3744 14178 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 3658 14178 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14138 3572 14178 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 18539 14166 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 18457 14166 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 18375 14166 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 18293 14166 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 18211 14166 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 18129 14166 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 18047 14166 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 17965 14166 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 17883 14166 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 17801 14166 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 17719 14166 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 17637 14166 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 17555 14166 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 17473 14166 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 17391 14166 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 17309 14166 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 17227 14166 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 17145 14166 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 17063 14166 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 16981 14166 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 16899 14166 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 16817 14166 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 16735 14166 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 16653 14166 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14126 16571 14166 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 16472 14162 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 16391 14162 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 16310 14162 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 16229 14162 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 16148 14162 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 16067 14162 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15986 14162 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15905 14162 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15824 14162 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15743 14162 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15662 14162 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15581 14162 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15500 14162 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15419 14162 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15338 14162 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15257 14162 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15176 14162 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15095 14162 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 15014 14162 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14933 14162 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14852 14162 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14771 14162 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14690 14162 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14609 14162 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14527 14162 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14445 14162 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14363 14162 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14281 14162 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14199 14162 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14117 14162 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 14035 14162 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 13953 14162 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 13871 14162 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 13789 14162 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 13707 14162 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14122 13625 14162 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 4432 14097 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 4346 14097 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 4260 14097 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 4174 14097 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 4088 14097 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 4002 14097 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 3916 14097 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 3830 14097 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 3744 14097 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 3658 14097 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14057 3572 14097 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 18539 14084 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 18457 14084 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 18375 14084 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 18293 14084 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 18211 14084 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 18129 14084 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 18047 14084 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 17965 14084 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 17883 14084 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 17801 14084 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 17719 14084 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 17637 14084 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 17555 14084 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 17473 14084 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 17391 14084 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 17309 14084 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 17227 14084 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 17145 14084 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 17063 14084 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 16981 14084 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 16899 14084 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 16817 14084 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 16735 14084 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 16653 14084 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14044 16571 14084 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 16472 14082 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 16391 14082 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 16310 14082 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 16229 14082 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 16148 14082 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 16067 14082 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15986 14082 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15905 14082 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15824 14082 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15743 14082 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15662 14082 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15581 14082 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15500 14082 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15419 14082 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15338 14082 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15257 14082 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15176 14082 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15095 14082 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 15014 14082 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14933 14082 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14852 14082 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14771 14082 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14690 14082 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14609 14082 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14527 14082 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14445 14082 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14363 14082 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14281 14082 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14199 14082 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14117 14082 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 14035 14082 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 13953 14082 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 13871 14082 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 13789 14082 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 13707 14082 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 14042 13625 14082 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 4432 14016 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 4346 14016 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 4260 14016 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 4174 14016 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 4088 14016 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 4002 14016 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 3916 14016 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 3830 14016 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 3744 14016 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 3658 14016 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13976 3572 14016 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 18539 14002 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 18457 14002 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 18375 14002 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 18293 14002 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 18211 14002 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 18129 14002 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 18047 14002 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 17965 14002 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 17883 14002 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 17801 14002 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 17719 14002 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 17637 14002 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 17555 14002 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 17473 14002 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 17391 14002 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 17309 14002 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 17227 14002 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 17145 14002 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 17063 14002 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16981 14002 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16899 14002 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16817 14002 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16735 14002 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16653 14002 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16571 14002 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16472 14002 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16391 14002 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16310 14002 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16229 14002 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16148 14002 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 16067 14002 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15986 14002 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15905 14002 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15824 14002 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15743 14002 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15662 14002 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15581 14002 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15500 14002 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15419 14002 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15338 14002 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15257 14002 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15176 14002 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15095 14002 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 15014 14002 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14933 14002 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14852 14002 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14771 14002 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14690 14002 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14609 14002 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14527 14002 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14445 14002 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14363 14002 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14281 14002 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14199 14002 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14117 14002 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 14035 14002 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 13953 14002 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 13871 14002 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 13789 14002 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 13707 14002 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13962 13625 14002 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 4432 13935 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 4346 13935 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 4260 13935 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 4174 13935 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 4088 13935 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 4002 13935 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 3916 13935 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 3830 13935 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 3744 13935 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 3658 13935 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13895 3572 13935 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 16472 13922 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 16391 13922 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 16310 13922 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 16229 13922 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 16148 13922 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 16067 13922 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15986 13922 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15905 13922 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15824 13922 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15743 13922 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15662 13922 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15581 13922 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15500 13922 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15419 13922 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15338 13922 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15257 13922 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15176 13922 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15095 13922 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 15014 13922 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14933 13922 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14852 13922 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14771 13922 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14690 13922 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14609 13922 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14527 13922 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14445 13922 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14363 13922 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14281 13922 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14199 13922 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14117 13922 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 14035 13922 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 13953 13922 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 13871 13922 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 13789 13922 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 13707 13922 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13882 13625 13922 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 18539 13920 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 18457 13920 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 18375 13920 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 18293 13920 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 18211 13920 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 18129 13920 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 18047 13920 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 17965 13920 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 17883 13920 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 17801 13920 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 17719 13920 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 17637 13920 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 17555 13920 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 17473 13920 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 17391 13920 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 17309 13920 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 17227 13920 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 17145 13920 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 17063 13920 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 16981 13920 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 16899 13920 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 16817 13920 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 16735 13920 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 16653 13920 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13880 16571 13920 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 4432 13854 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 4346 13854 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 4260 13854 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 4174 13854 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 4088 13854 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 4002 13854 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 3916 13854 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 3830 13854 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 3744 13854 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 3658 13854 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13814 3572 13854 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 16472 13842 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 16391 13842 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 16310 13842 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 16229 13842 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 16148 13842 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 16067 13842 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15986 13842 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15905 13842 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15824 13842 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15743 13842 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15662 13842 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15581 13842 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15500 13842 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15419 13842 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15338 13842 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15257 13842 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15176 13842 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15095 13842 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 15014 13842 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14933 13842 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14852 13842 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14771 13842 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14690 13842 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14609 13842 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14527 13842 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14445 13842 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14363 13842 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14281 13842 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14199 13842 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14117 13842 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 14035 13842 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 13953 13842 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 13871 13842 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 13789 13842 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 13707 13842 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13802 13625 13842 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 18539 13838 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 18457 13838 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 18375 13838 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 18293 13838 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 18211 13838 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 18129 13838 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 18047 13838 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 17965 13838 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 17883 13838 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 17801 13838 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 17719 13838 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 17637 13838 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 17555 13838 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 17473 13838 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 17391 13838 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 17309 13838 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 17227 13838 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 17145 13838 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 17063 13838 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 16981 13838 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 16899 13838 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 16817 13838 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 16735 13838 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 16653 13838 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13798 16571 13838 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 4432 13773 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 4346 13773 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 4260 13773 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 4174 13773 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 4088 13773 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 4002 13773 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 3916 13773 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 3830 13773 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 3744 13773 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 3658 13773 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13733 3572 13773 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 16472 13762 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 16391 13762 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 16310 13762 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 16229 13762 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 16148 13762 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 16067 13762 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15986 13762 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15905 13762 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15824 13762 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15743 13762 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15662 13762 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15581 13762 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15500 13762 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15419 13762 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15338 13762 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15257 13762 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15176 13762 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15095 13762 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 15014 13762 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14933 13762 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14852 13762 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14771 13762 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14690 13762 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14609 13762 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14527 13762 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14445 13762 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14363 13762 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14281 13762 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14199 13762 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14117 13762 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 14035 13762 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 13953 13762 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 13871 13762 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 13789 13762 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 13707 13762 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13722 13625 13762 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 18539 13756 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 18457 13756 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 18375 13756 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 18293 13756 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 18211 13756 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 18129 13756 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 18047 13756 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 17965 13756 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 17883 13756 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 17801 13756 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 17719 13756 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 17637 13756 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 17555 13756 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 17473 13756 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 17391 13756 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 17309 13756 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 17227 13756 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 17145 13756 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 17063 13756 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 16981 13756 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 16899 13756 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 16817 13756 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 16735 13756 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 16653 13756 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13716 16571 13756 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 4432 13692 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 4346 13692 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 4260 13692 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 4174 13692 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 4088 13692 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 4002 13692 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 3916 13692 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 3830 13692 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 3744 13692 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 3658 13692 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13652 3572 13692 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 16472 13682 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 16391 13682 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 16310 13682 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 16229 13682 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 16148 13682 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 16067 13682 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15986 13682 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15905 13682 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15824 13682 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15743 13682 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15662 13682 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15581 13682 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15500 13682 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15419 13682 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15338 13682 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15257 13682 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15176 13682 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15095 13682 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 15014 13682 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14933 13682 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14852 13682 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14771 13682 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14690 13682 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14609 13682 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14527 13682 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14445 13682 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14363 13682 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14281 13682 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14199 13682 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14117 13682 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 14035 13682 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 13953 13682 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 13871 13682 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 13789 13682 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 13707 13682 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13642 13625 13682 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 18539 13674 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 18457 13674 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 18375 13674 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 18293 13674 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 18211 13674 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 18129 13674 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 18047 13674 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 17965 13674 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 17883 13674 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 17801 13674 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 17719 13674 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 17637 13674 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 17555 13674 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 17473 13674 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 17391 13674 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 17309 13674 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 17227 13674 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 17145 13674 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 17063 13674 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 16981 13674 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 16899 13674 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 16817 13674 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 16735 13674 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 16653 13674 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13634 16571 13674 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 4432 13611 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 4346 13611 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 4260 13611 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 4174 13611 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 4088 13611 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 4002 13611 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 3916 13611 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 3830 13611 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 3744 13611 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 3658 13611 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13571 3572 13611 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 16472 13602 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 16391 13602 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 16310 13602 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 16229 13602 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 16148 13602 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 16067 13602 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15986 13602 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15905 13602 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15824 13602 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15743 13602 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15662 13602 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15581 13602 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15500 13602 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15419 13602 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15338 13602 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15257 13602 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15176 13602 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15095 13602 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 15014 13602 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14933 13602 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14852 13602 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14771 13602 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14690 13602 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14609 13602 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14527 13602 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14445 13602 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14363 13602 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14281 13602 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14199 13602 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14117 13602 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 14035 13602 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 13953 13602 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 13871 13602 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 13789 13602 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 13707 13602 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13562 13625 13602 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 18539 13592 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 18457 13592 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 18375 13592 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 18293 13592 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 18211 13592 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 18129 13592 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 18047 13592 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 17965 13592 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 17883 13592 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 17801 13592 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 17719 13592 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 17637 13592 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 17555 13592 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 17473 13592 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 17391 13592 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 17309 13592 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 17227 13592 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 17145 13592 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 17063 13592 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 16981 13592 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 16899 13592 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 16817 13592 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 16735 13592 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 16653 13592 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13552 16571 13592 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 4432 13530 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 4346 13530 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 4260 13530 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 4174 13530 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 4088 13530 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 4002 13530 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 3916 13530 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 3830 13530 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 3744 13530 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 3658 13530 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13490 3572 13530 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 16472 13522 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 16391 13522 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 16310 13522 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 16229 13522 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 16148 13522 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 16067 13522 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15986 13522 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15905 13522 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15824 13522 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15743 13522 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15662 13522 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15581 13522 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15500 13522 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15419 13522 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15338 13522 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15257 13522 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15176 13522 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15095 13522 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 15014 13522 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14933 13522 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14852 13522 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14771 13522 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14690 13522 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14609 13522 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14527 13522 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14445 13522 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14363 13522 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14281 13522 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14199 13522 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14117 13522 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 14035 13522 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 13953 13522 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 13871 13522 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 13789 13522 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 13707 13522 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13482 13625 13522 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 18539 13510 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 18457 13510 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 18375 13510 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 18293 13510 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 18211 13510 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 18129 13510 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 18047 13510 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 17965 13510 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 17883 13510 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 17801 13510 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 17719 13510 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 17637 13510 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 17555 13510 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 17473 13510 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 17391 13510 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 17309 13510 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 17227 13510 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 17145 13510 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 17063 13510 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 16981 13510 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 16899 13510 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 16817 13510 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 16735 13510 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 16653 13510 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13470 16571 13510 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 4432 13449 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 4346 13449 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 4260 13449 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 4174 13449 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 4088 13449 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 4002 13449 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 3916 13449 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 3830 13449 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 3744 13449 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 3658 13449 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13409 3572 13449 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 16472 13442 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 16391 13442 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 16310 13442 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 16229 13442 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 16148 13442 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 16067 13442 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15986 13442 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15905 13442 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15824 13442 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15743 13442 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15662 13442 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15581 13442 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15500 13442 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15419 13442 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15338 13442 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15257 13442 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15176 13442 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15095 13442 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 15014 13442 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14933 13442 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14852 13442 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14771 13442 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14690 13442 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14609 13442 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14527 13442 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14445 13442 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14363 13442 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14281 13442 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14199 13442 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14117 13442 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 14035 13442 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 13953 13442 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 13871 13442 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 13789 13442 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 13707 13442 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13402 13625 13442 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 18539 13428 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 18457 13428 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 18375 13428 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 18293 13428 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 18211 13428 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 18129 13428 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 18047 13428 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 17965 13428 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 17883 13428 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 17801 13428 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 17719 13428 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 17637 13428 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 17555 13428 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 17473 13428 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 17391 13428 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 17309 13428 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 17227 13428 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 17145 13428 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 17063 13428 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 16981 13428 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 16899 13428 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 16817 13428 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 16735 13428 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 16653 13428 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13388 16571 13428 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 4432 13368 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 4346 13368 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 4260 13368 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 4174 13368 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 4088 13368 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 4002 13368 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 3916 13368 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 3830 13368 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 3744 13368 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 3658 13368 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13328 3572 13368 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 16472 13362 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 16391 13362 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 16310 13362 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 16229 13362 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 16148 13362 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 16067 13362 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15986 13362 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15905 13362 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15824 13362 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15743 13362 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15662 13362 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15581 13362 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15500 13362 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15419 13362 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15338 13362 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15257 13362 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15176 13362 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15095 13362 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 15014 13362 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14933 13362 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14852 13362 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14771 13362 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14690 13362 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14609 13362 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14527 13362 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14445 13362 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14363 13362 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14281 13362 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14199 13362 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14117 13362 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 14035 13362 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 13953 13362 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 13871 13362 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 13789 13362 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 13707 13362 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13322 13625 13362 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 18539 13346 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 18457 13346 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 18375 13346 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 18293 13346 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 18211 13346 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 18129 13346 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 18047 13346 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 17965 13346 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 17883 13346 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 17801 13346 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 17719 13346 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 17637 13346 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 17555 13346 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 17473 13346 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 17391 13346 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 17309 13346 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 17227 13346 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 17145 13346 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 17063 13346 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 16981 13346 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 16899 13346 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 16817 13346 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 16735 13346 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 16653 13346 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13306 16571 13346 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 4432 13287 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 4346 13287 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 4260 13287 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 4174 13287 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 4088 13287 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 4002 13287 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 3916 13287 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 3830 13287 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 3744 13287 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 3658 13287 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13247 3572 13287 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 16472 13282 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 16391 13282 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 16310 13282 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 16229 13282 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 16148 13282 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 16067 13282 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15986 13282 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15905 13282 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15824 13282 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15743 13282 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15662 13282 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15581 13282 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15500 13282 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15419 13282 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15338 13282 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15257 13282 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15176 13282 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15095 13282 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 15014 13282 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14933 13282 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14852 13282 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14771 13282 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14690 13282 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14609 13282 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14527 13282 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14445 13282 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14363 13282 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14281 13282 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14199 13282 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14117 13282 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 14035 13282 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 13953 13282 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 13871 13282 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 13789 13282 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 13707 13282 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13242 13625 13282 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 18539 13264 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 18457 13264 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 18375 13264 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 18293 13264 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 18211 13264 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 18129 13264 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 18047 13264 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 17965 13264 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 17883 13264 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 17801 13264 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 17719 13264 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 17637 13264 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 17555 13264 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 17473 13264 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 17391 13264 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 17309 13264 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 17227 13264 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 17145 13264 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 17063 13264 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 16981 13264 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 16899 13264 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 16817 13264 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 16735 13264 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 16653 13264 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13224 16571 13264 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 4432 13206 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 4346 13206 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 4260 13206 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 4174 13206 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 4088 13206 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 4002 13206 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 3916 13206 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 3830 13206 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 3744 13206 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 3658 13206 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13166 3572 13206 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 16472 13202 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 16391 13202 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 16310 13202 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 16229 13202 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 16148 13202 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 16067 13202 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15986 13202 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15905 13202 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15824 13202 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15743 13202 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15662 13202 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15581 13202 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15500 13202 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15419 13202 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15338 13202 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15257 13202 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15176 13202 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15095 13202 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 15014 13202 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14933 13202 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14852 13202 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14771 13202 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14690 13202 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14609 13202 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14527 13202 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14445 13202 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14363 13202 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14281 13202 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14199 13202 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14117 13202 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 14035 13202 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 13953 13202 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 13871 13202 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 13789 13202 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 13707 13202 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13162 13625 13202 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 18539 13182 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 18457 13182 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 18375 13182 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 18293 13182 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 18211 13182 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 18129 13182 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 18047 13182 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 17965 13182 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 17883 13182 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 17801 13182 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 17719 13182 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 17637 13182 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 17555 13182 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 17473 13182 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 17391 13182 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 17309 13182 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 17227 13182 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 17145 13182 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 17063 13182 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 16981 13182 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 16899 13182 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 16817 13182 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 16735 13182 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 16653 13182 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13142 16571 13182 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 4432 13125 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 4346 13125 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 4260 13125 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 4174 13125 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 4088 13125 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 4002 13125 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 3916 13125 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 3830 13125 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 3744 13125 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 3658 13125 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13085 3572 13125 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 16472 13122 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 16391 13122 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 16310 13122 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 16229 13122 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 16148 13122 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 16067 13122 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15986 13122 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15905 13122 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15824 13122 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15743 13122 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15662 13122 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15581 13122 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15500 13122 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15419 13122 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15338 13122 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15257 13122 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15176 13122 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15095 13122 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 15014 13122 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14933 13122 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14852 13122 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14771 13122 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14690 13122 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14609 13122 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14527 13122 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14445 13122 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14363 13122 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14281 13122 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14199 13122 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14117 13122 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 14035 13122 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 13953 13122 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 13871 13122 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 13789 13122 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 13707 13122 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13082 13625 13122 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 18539 13100 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 18457 13100 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 18375 13100 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 18293 13100 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 18211 13100 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 18129 13100 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 18047 13100 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 17965 13100 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 17883 13100 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 17801 13100 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 17719 13100 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 17637 13100 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 17555 13100 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 17473 13100 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 17391 13100 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 17309 13100 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 17227 13100 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 17145 13100 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 17063 13100 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 16981 13100 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 16899 13100 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 16817 13100 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 16735 13100 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 16653 13100 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13060 16571 13100 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 4432 13044 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 4346 13044 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 4260 13044 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 4174 13044 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 4088 13044 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 4002 13044 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 3916 13044 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 3830 13044 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 3744 13044 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 3658 13044 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13004 3572 13044 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 16472 13042 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 16391 13042 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 16310 13042 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 16229 13042 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 16148 13042 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 16067 13042 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15986 13042 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15905 13042 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15824 13042 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15743 13042 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15662 13042 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15581 13042 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15500 13042 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15419 13042 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15338 13042 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15257 13042 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15176 13042 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15095 13042 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 15014 13042 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14933 13042 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14852 13042 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14771 13042 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14690 13042 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14609 13042 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14527 13042 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14445 13042 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14363 13042 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14281 13042 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14199 13042 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14117 13042 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 14035 13042 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 13953 13042 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 13871 13042 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 13789 13042 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 13707 13042 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 13002 13625 13042 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 18539 13018 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 18457 13018 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 18375 13018 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 18293 13018 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 18211 13018 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 18129 13018 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 18047 13018 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 17965 13018 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 17883 13018 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 17801 13018 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 17719 13018 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 17637 13018 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 17555 13018 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 17473 13018 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 17391 13018 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 17309 13018 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 17227 13018 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 17145 13018 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 17063 13018 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 16981 13018 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 16899 13018 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 16817 13018 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 16735 13018 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 16653 13018 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12978 16571 13018 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 4432 12963 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 4346 12963 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 4260 12963 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 4174 12963 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 4088 12963 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 4002 12963 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 3916 12963 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 3830 12963 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 3744 12963 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 3658 12963 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12923 3572 12963 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 16472 12962 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 16391 12962 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 16310 12962 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 16229 12962 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 16148 12962 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 16067 12962 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15986 12962 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15905 12962 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15824 12962 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15743 12962 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15662 12962 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15581 12962 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15500 12962 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15419 12962 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15338 12962 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15257 12962 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15176 12962 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15095 12962 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 15014 12962 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14933 12962 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14852 12962 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14771 12962 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14690 12962 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14609 12962 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14527 12962 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14445 12962 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14363 12962 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14281 12962 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14199 12962 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14117 12962 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 14035 12962 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 13953 12962 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 13871 12962 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 13789 12962 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 13707 12962 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12922 13625 12962 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 18539 12936 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 18457 12936 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 18375 12936 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 18293 12936 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 18211 12936 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 18129 12936 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 18047 12936 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 17965 12936 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 17883 12936 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 17801 12936 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 17719 12936 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 17637 12936 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 17555 12936 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 17473 12936 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 17391 12936 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 17309 12936 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 17227 12936 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 17145 12936 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 17063 12936 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 16981 12936 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 16899 12936 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 16817 12936 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 16735 12936 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 16653 12936 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12896 16571 12936 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 16472 12882 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 16391 12882 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 16310 12882 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 16229 12882 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 16148 12882 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 16067 12882 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15986 12882 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15905 12882 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15824 12882 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15743 12882 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15662 12882 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15581 12882 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15500 12882 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15419 12882 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15338 12882 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15257 12882 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15176 12882 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15095 12882 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 15014 12882 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14933 12882 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14852 12882 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14771 12882 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14690 12882 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14609 12882 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14527 12882 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14445 12882 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14363 12882 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14281 12882 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14199 12882 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14117 12882 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 14035 12882 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 13953 12882 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 13871 12882 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 13789 12882 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 13707 12882 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 13625 12882 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 4432 12882 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 4346 12882 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 4260 12882 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 4174 12882 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 4088 12882 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 4002 12882 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 3916 12882 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 3830 12882 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 3744 12882 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 3658 12882 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12842 3572 12882 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 18539 12854 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 18457 12854 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 18375 12854 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 18293 12854 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 18211 12854 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 18129 12854 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 18047 12854 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 17965 12854 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 17883 12854 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 17801 12854 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 17719 12854 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 17637 12854 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 17555 12854 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 17473 12854 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 17391 12854 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 17309 12854 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 17227 12854 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 17145 12854 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 17063 12854 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 16981 12854 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 16899 12854 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 16817 12854 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 16735 12854 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 16653 12854 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12814 16571 12854 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 16472 12802 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 16391 12802 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 16310 12802 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 16229 12802 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 16148 12802 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 16067 12802 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15986 12802 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15905 12802 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15824 12802 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15743 12802 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15662 12802 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15581 12802 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15500 12802 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15419 12802 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15338 12802 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15257 12802 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15176 12802 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15095 12802 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 15014 12802 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14933 12802 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14852 12802 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14771 12802 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14690 12802 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14609 12802 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14527 12802 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14445 12802 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14363 12802 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14281 12802 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14199 12802 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14117 12802 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 14035 12802 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 13953 12802 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 13871 12802 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 13789 12802 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 13707 12802 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12762 13625 12802 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 4432 12801 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 4346 12801 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 4260 12801 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 4174 12801 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 4088 12801 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 4002 12801 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 3916 12801 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 3830 12801 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 3744 12801 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 3658 12801 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12761 3572 12801 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 18539 12772 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 18457 12772 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 18375 12772 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 18293 12772 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 18211 12772 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 18129 12772 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 18047 12772 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 17965 12772 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 17883 12772 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 17801 12772 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 17719 12772 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 17637 12772 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 17555 12772 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 17473 12772 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 17391 12772 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 17309 12772 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 17227 12772 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 17145 12772 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 17063 12772 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 16981 12772 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 16899 12772 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 16817 12772 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 16735 12772 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 16653 12772 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12732 16571 12772 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 16472 12722 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 16391 12722 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 16310 12722 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 16229 12722 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 16148 12722 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 16067 12722 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15986 12722 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15905 12722 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15824 12722 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15743 12722 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15662 12722 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15581 12722 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15500 12722 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15419 12722 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15338 12722 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15257 12722 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15176 12722 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15095 12722 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 15014 12722 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14933 12722 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14852 12722 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14771 12722 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14690 12722 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14609 12722 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14527 12722 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14445 12722 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14363 12722 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14281 12722 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14199 12722 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14117 12722 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 14035 12722 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 13953 12722 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 13871 12722 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 13789 12722 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 13707 12722 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12682 13625 12722 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 4432 12720 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 4346 12720 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 4260 12720 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 4174 12720 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 4088 12720 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 4002 12720 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 3916 12720 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 3830 12720 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 3744 12720 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 3658 12720 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12680 3572 12720 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 18539 12690 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 18457 12690 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 18375 12690 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 18293 12690 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 18211 12690 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 18129 12690 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 18047 12690 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 17965 12690 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 17883 12690 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 17801 12690 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 17719 12690 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 17637 12690 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 17555 12690 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 17473 12690 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 17391 12690 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 17309 12690 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 17227 12690 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 17145 12690 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 17063 12690 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 16981 12690 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 16899 12690 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 16817 12690 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 16735 12690 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 16653 12690 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12650 16571 12690 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 16472 12642 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 16391 12642 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 16310 12642 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 16229 12642 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 16148 12642 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 16067 12642 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15986 12642 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15905 12642 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15824 12642 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15743 12642 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15662 12642 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15581 12642 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15500 12642 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15419 12642 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15338 12642 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15257 12642 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15176 12642 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15095 12642 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 15014 12642 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14933 12642 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14852 12642 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14771 12642 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14690 12642 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14609 12642 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14527 12642 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14445 12642 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14363 12642 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14281 12642 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14199 12642 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14117 12642 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 14035 12642 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 13953 12642 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 13871 12642 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 13789 12642 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 13707 12642 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12602 13625 12642 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 4432 12639 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 4346 12639 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 4260 12639 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 4174 12639 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 4088 12639 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 4002 12639 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 3916 12639 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 3830 12639 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 3744 12639 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 3658 12639 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12599 3572 12639 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 18539 12608 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 18457 12608 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 18375 12608 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 18293 12608 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 18211 12608 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 18129 12608 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 18047 12608 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 17965 12608 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 17883 12608 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 17801 12608 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 17719 12608 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 17637 12608 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 17555 12608 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 17473 12608 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 17391 12608 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 17309 12608 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 17227 12608 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 17145 12608 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 17063 12608 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 16981 12608 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 16899 12608 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 16817 12608 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 16735 12608 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 16653 12608 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12568 16571 12608 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 16472 12562 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 16391 12562 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 16310 12562 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 16229 12562 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 16148 12562 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 16067 12562 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15986 12562 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15905 12562 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15824 12562 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15743 12562 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15662 12562 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15581 12562 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15500 12562 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15419 12562 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15338 12562 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15257 12562 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15176 12562 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15095 12562 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 15014 12562 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14933 12562 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14852 12562 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14771 12562 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14690 12562 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14609 12562 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14527 12562 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14445 12562 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14363 12562 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14281 12562 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14199 12562 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14117 12562 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 14035 12562 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 13953 12562 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 13871 12562 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 13789 12562 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 13707 12562 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12522 13625 12562 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 4432 12558 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 4346 12558 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 4260 12558 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 4174 12558 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 4088 12558 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 4002 12558 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 3916 12558 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 3830 12558 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 3744 12558 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 3658 12558 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12518 3572 12558 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 18539 12526 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 18457 12526 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 18375 12526 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 18293 12526 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 18211 12526 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 18129 12526 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 18047 12526 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 17965 12526 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 17883 12526 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 17801 12526 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 17719 12526 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 17637 12526 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 17555 12526 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 17473 12526 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 17391 12526 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 17309 12526 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 17227 12526 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 17145 12526 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 17063 12526 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 16981 12526 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 16899 12526 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 16817 12526 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 16735 12526 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 16653 12526 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12486 16571 12526 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 16472 12482 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 16391 12482 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 16310 12482 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 16229 12482 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 16148 12482 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 16067 12482 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15986 12482 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15905 12482 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15824 12482 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15743 12482 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15662 12482 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15581 12482 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15500 12482 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15419 12482 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15338 12482 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15257 12482 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15176 12482 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15095 12482 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 15014 12482 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14933 12482 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14852 12482 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14771 12482 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14690 12482 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14609 12482 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14527 12482 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14445 12482 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14363 12482 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14281 12482 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14199 12482 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14117 12482 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 14035 12482 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 13953 12482 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 13871 12482 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 13789 12482 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 13707 12482 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12442 13625 12482 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 4432 12477 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 4346 12477 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 4260 12477 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 4174 12477 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 4088 12477 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 4002 12477 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 3916 12477 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 3830 12477 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 3744 12477 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 3658 12477 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12437 3572 12477 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 18539 12445 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 18457 12445 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 18375 12445 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 18293 12445 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 18211 12445 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 18129 12445 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 18047 12445 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 17965 12445 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 17883 12445 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 17801 12445 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 17719 12445 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 17637 12445 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 17555 12445 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 17473 12445 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 17391 12445 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 17309 12445 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 17227 12445 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 17145 12445 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 17063 12445 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 16981 12445 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 16899 12445 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 16817 12445 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 16735 12445 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 16653 12445 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12405 16571 12445 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 16472 12402 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 16391 12402 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 16310 12402 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 16229 12402 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 16148 12402 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 16067 12402 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15986 12402 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15905 12402 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15824 12402 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15743 12402 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15662 12402 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15581 12402 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15500 12402 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15419 12402 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15338 12402 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15257 12402 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15176 12402 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15095 12402 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 15014 12402 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14933 12402 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14852 12402 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14771 12402 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14690 12402 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14609 12402 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14527 12402 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14445 12402 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14363 12402 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14281 12402 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14199 12402 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14117 12402 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 14035 12402 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 13953 12402 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 13871 12402 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 13789 12402 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 13707 12402 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12362 13625 12402 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 4432 12396 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 4346 12396 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 4260 12396 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 4174 12396 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 4088 12396 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 4002 12396 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 3916 12396 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 3830 12396 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 3744 12396 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 3658 12396 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12356 3572 12396 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 18539 12364 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 18457 12364 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 18375 12364 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 18293 12364 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 18211 12364 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 18129 12364 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 18047 12364 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 17965 12364 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 17883 12364 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 17801 12364 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 17719 12364 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 17637 12364 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 17555 12364 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 17473 12364 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 17391 12364 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 17309 12364 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 17227 12364 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 17145 12364 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 17063 12364 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 16981 12364 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 16899 12364 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 16817 12364 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 16735 12364 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 16653 12364 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12324 16571 12364 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 16472 12322 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 16391 12322 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 16310 12322 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 16229 12322 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 16148 12322 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 16067 12322 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15986 12322 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15905 12322 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15824 12322 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15743 12322 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15662 12322 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15581 12322 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15500 12322 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15419 12322 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15338 12322 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15257 12322 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15176 12322 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15095 12322 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 15014 12322 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14933 12322 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14852 12322 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14771 12322 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14690 12322 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14609 12322 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14527 12322 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14445 12322 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14363 12322 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14281 12322 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14199 12322 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14117 12322 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 14035 12322 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 13953 12322 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 13871 12322 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 13789 12322 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 13707 12322 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12282 13625 12322 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 4432 12315 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 4346 12315 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 4260 12315 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 4174 12315 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 4088 12315 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 4002 12315 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 3916 12315 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 3830 12315 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 3744 12315 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 3658 12315 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12275 3572 12315 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 18539 12283 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 18457 12283 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 18375 12283 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 18293 12283 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 18211 12283 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 18129 12283 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 18047 12283 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 17965 12283 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 17883 12283 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 17801 12283 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 17719 12283 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 17637 12283 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 17555 12283 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 17473 12283 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 17391 12283 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 17309 12283 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 17227 12283 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 17145 12283 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 17063 12283 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 16981 12283 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 16899 12283 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 16817 12283 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 16735 12283 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 16653 12283 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12243 16571 12283 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 16472 12242 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 16391 12242 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 16310 12242 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 16229 12242 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 16148 12242 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 16067 12242 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15986 12242 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15905 12242 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15824 12242 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15743 12242 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15662 12242 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15581 12242 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15500 12242 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15419 12242 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15338 12242 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15257 12242 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15176 12242 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15095 12242 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 15014 12242 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14933 12242 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14852 12242 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14771 12242 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14690 12242 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14609 12242 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14527 12242 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14445 12242 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14363 12242 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14281 12242 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14199 12242 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14117 12242 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 14035 12242 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 13953 12242 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 13871 12242 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 13789 12242 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 13707 12242 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12202 13625 12242 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 4432 12234 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 4346 12234 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 4260 12234 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 4174 12234 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 4088 12234 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 4002 12234 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 3916 12234 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 3830 12234 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 3744 12234 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 3658 12234 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12194 3572 12234 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12147 18289 12187 18329 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12147 18203 12187 18243 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12143 18111 12183 18151 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12143 18025 12183 18065 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12143 17939 12183 17979 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12143 17853 12183 17893 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12143 17767 12183 17807 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12143 17682 12183 17722 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 16472 12162 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 16391 12162 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 16310 12162 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 16229 12162 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 16148 12162 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 16067 12162 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15986 12162 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15905 12162 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15824 12162 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15743 12162 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15662 12162 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15581 12162 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15500 12162 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15419 12162 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15338 12162 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15257 12162 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15176 12162 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15095 12162 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 15014 12162 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14933 12162 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14852 12162 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14771 12162 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14690 12162 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14609 12162 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14527 12162 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14445 12162 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14363 12162 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14281 12162 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14199 12162 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14117 12162 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 14035 12162 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 13953 12162 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 13871 12162 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 13789 12162 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 13707 12162 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12122 13625 12162 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12118 17575 12158 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12118 17494 12158 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12118 17413 12158 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12118 17332 12158 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12118 17251 12158 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12118 17171 12158 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12118 17091 12158 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12118 17011 12158 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12118 16931 12158 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12118 16851 12158 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12118 16771 12158 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12118 16691 12158 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12118 16611 12158 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 4432 12153 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 4346 12153 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 4260 12153 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 4174 12153 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 4088 12153 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 4002 12153 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 3916 12153 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 3830 12153 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 3744 12153 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 3658 12153 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12113 3572 12153 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12061 18111 12101 18151 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12061 18025 12101 18065 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12061 17939 12101 17979 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12061 17853 12101 17893 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12061 17767 12101 17807 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12061 17682 12101 17722 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 16472 12082 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 16391 12082 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 16310 12082 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 16229 12082 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 16148 12082 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 16067 12082 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15986 12082 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15905 12082 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15824 12082 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15743 12082 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15662 12082 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15581 12082 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15500 12082 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15419 12082 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15338 12082 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15257 12082 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15176 12082 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15095 12082 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 15014 12082 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14933 12082 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14852 12082 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14771 12082 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14690 12082 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14609 12082 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14527 12082 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14445 12082 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14363 12082 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14281 12082 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14199 12082 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14117 12082 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 14035 12082 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 13953 12082 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 13871 12082 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 13789 12082 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 13707 12082 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12042 13625 12082 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12036 17575 12076 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12036 17494 12076 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12036 17413 12076 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12036 17332 12076 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12036 17251 12076 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12036 17171 12076 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12036 17091 12076 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12036 17011 12076 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12036 16931 12076 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12036 16851 12076 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12036 16771 12076 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12036 16691 12076 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12036 16611 12076 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 4432 12072 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 4346 12072 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 4260 12072 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 4174 12072 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 4088 12072 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 4002 12072 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 3916 12072 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 3830 12072 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 3744 12072 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 3658 12072 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 12032 3572 12072 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11991 18289 12031 18329 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11991 18203 12031 18243 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11979 18111 12019 18151 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11979 18025 12019 18065 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11979 17939 12019 17979 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11979 17853 12019 17893 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11979 17767 12019 17807 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11979 17682 12019 17722 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 16472 12002 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 16391 12002 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 16310 12002 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 16229 12002 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 16148 12002 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 16067 12002 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15986 12002 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15905 12002 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15824 12002 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15743 12002 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15662 12002 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15581 12002 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15500 12002 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15419 12002 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15338 12002 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15257 12002 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15176 12002 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15095 12002 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 15014 12002 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14933 12002 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14852 12002 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14771 12002 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14690 12002 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14609 12002 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14527 12002 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14445 12002 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14363 12002 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14281 12002 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14199 12002 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14117 12002 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 14035 12002 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 13953 12002 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 13871 12002 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 13789 12002 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 13707 12002 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11962 13625 12002 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11954 17575 11994 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11954 17494 11994 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11954 17413 11994 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11954 17332 11994 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11954 17251 11994 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11954 17171 11994 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11954 17091 11994 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11954 17011 11994 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11954 16931 11994 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11954 16851 11994 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11954 16771 11994 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11954 16691 11994 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11954 16611 11994 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 4432 11991 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 4346 11991 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 4260 11991 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 4174 11991 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 4088 11991 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 4002 11991 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 3916 11991 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 3830 11991 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 3744 11991 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 3658 11991 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11951 3572 11991 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11897 18111 11937 18151 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11897 18025 11937 18065 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11897 17939 11937 17979 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11897 17853 11937 17893 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11897 17767 11937 17807 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11897 17682 11937 17722 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 16472 11922 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 16391 11922 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 16310 11922 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 16229 11922 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 16148 11922 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 16067 11922 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15986 11922 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15905 11922 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15824 11922 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15743 11922 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15662 11922 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15581 11922 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15500 11922 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15419 11922 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15338 11922 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15257 11922 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15176 11922 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15095 11922 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 15014 11922 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14933 11922 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14852 11922 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14771 11922 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14690 11922 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14609 11922 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14527 11922 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14445 11922 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14363 11922 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14281 11922 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14199 11922 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14117 11922 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 14035 11922 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 13953 11922 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 13871 11922 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 13789 11922 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 13707 11922 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11882 13625 11922 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11872 17575 11912 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11872 17494 11912 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11872 17413 11912 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11872 17332 11912 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11872 17251 11912 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11872 17171 11912 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11872 17091 11912 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11872 17011 11912 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11872 16931 11912 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11872 16851 11912 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11872 16771 11912 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11872 16691 11912 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11872 16611 11912 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 4432 11910 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 4346 11910 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 4260 11910 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 4174 11910 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 4088 11910 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 4002 11910 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 3916 11910 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 3830 11910 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 3744 11910 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 3658 11910 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11870 3572 11910 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11815 18111 11855 18151 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11815 18025 11855 18065 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11815 17939 11855 17979 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11815 17853 11855 17893 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11815 17767 11855 17807 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11815 17682 11855 17722 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 16472 11842 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 16391 11842 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 16310 11842 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 16229 11842 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 16148 11842 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 16067 11842 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15986 11842 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15905 11842 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15824 11842 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15743 11842 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15662 11842 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15581 11842 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15500 11842 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15419 11842 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15338 11842 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15257 11842 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15176 11842 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15095 11842 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 15014 11842 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14933 11842 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14852 11842 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14771 11842 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14690 11842 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14609 11842 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14527 11842 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14445 11842 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14363 11842 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14281 11842 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14199 11842 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14117 11842 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 14035 11842 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 13953 11842 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 13871 11842 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 13789 11842 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 13707 11842 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11802 13625 11842 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 17575 11830 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 17494 11830 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 17413 11830 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 17332 11830 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 17251 11830 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 17171 11830 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 17091 11830 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 17011 11830 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 16931 11830 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 16851 11830 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 16771 11830 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 16691 11830 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11790 16611 11830 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 4432 11829 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 4346 11829 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 4260 11829 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 4174 11829 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 4088 11829 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 4002 11829 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 3916 11829 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 3830 11829 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 3744 11829 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 3658 11829 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11789 3572 11829 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 16472 11762 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 16391 11762 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 16310 11762 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 16229 11762 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 16148 11762 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 16067 11762 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15986 11762 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15905 11762 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15824 11762 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15743 11762 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15662 11762 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15581 11762 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15500 11762 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15419 11762 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15338 11762 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15257 11762 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15176 11762 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15095 11762 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 15014 11762 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14933 11762 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14852 11762 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14771 11762 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14690 11762 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14609 11762 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14527 11762 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14445 11762 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14363 11762 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14281 11762 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14199 11762 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14117 11762 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 14035 11762 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 13953 11762 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 13871 11762 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 13789 11762 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 13707 11762 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11722 13625 11762 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11715 17853 11755 17893 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11715 17769 11755 17809 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11715 17686 11755 17726 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 17575 11748 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 17494 11748 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 17413 11748 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 17332 11748 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 17251 11748 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 17171 11748 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 17091 11748 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 17011 11748 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 16931 11748 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 16851 11748 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 16771 11748 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 16691 11748 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 16611 11748 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 4432 11748 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 4346 11748 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 4260 11748 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 4174 11748 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 4088 11748 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 4002 11748 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 3916 11748 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 3830 11748 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 3744 11748 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 3658 11748 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11708 3572 11748 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 16472 11682 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 16391 11682 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 16310 11682 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 16229 11682 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 16148 11682 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 16067 11682 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15986 11682 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15905 11682 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15824 11682 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15743 11682 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15662 11682 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15581 11682 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15500 11682 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15419 11682 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15338 11682 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15257 11682 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15176 11682 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15095 11682 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 15014 11682 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14933 11682 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14852 11682 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14771 11682 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14690 11682 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14609 11682 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14527 11682 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14445 11682 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14363 11682 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14281 11682 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14199 11682 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14117 11682 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 14035 11682 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 13953 11682 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 13871 11682 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 13789 11682 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 13707 11682 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11642 13625 11682 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 4432 11667 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 4346 11667 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 4260 11667 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 4174 11667 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 4088 11667 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 4002 11667 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 3916 11667 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 3830 11667 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 3744 11667 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 3658 11667 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11627 3572 11667 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11626 17575 11666 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11626 17494 11666 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11626 17413 11666 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11626 17332 11666 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11626 17251 11666 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11626 17171 11666 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11626 17091 11666 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11626 17011 11666 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11626 16931 11666 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11626 16851 11666 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11626 16771 11666 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11626 16691 11666 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11626 16611 11666 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 16472 11602 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 16391 11602 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 16310 11602 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 16229 11602 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 16148 11602 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 16067 11602 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15986 11602 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15905 11602 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15824 11602 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15743 11602 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15662 11602 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15581 11602 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15500 11602 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15419 11602 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15338 11602 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15257 11602 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15176 11602 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15095 11602 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 15014 11602 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14933 11602 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14852 11602 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14771 11602 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14690 11602 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14609 11602 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14527 11602 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14445 11602 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14363 11602 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14281 11602 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14199 11602 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14117 11602 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 14035 11602 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 13953 11602 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 13871 11602 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 13789 11602 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 13707 11602 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11562 13625 11602 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11559 17853 11599 17893 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11559 17769 11599 17809 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11559 17686 11599 17726 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 4432 11586 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 4346 11586 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 4260 11586 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 4174 11586 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 4088 11586 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 4002 11586 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 3916 11586 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 3830 11586 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 3744 11586 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 3658 11586 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11546 3572 11586 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11544 17575 11584 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11544 17494 11584 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11544 17413 11584 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11544 17332 11584 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11544 17251 11584 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11544 17171 11584 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11544 17091 11584 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11544 17011 11584 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11544 16931 11584 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11544 16851 11584 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11544 16771 11584 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11544 16691 11584 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11544 16611 11584 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 16472 11522 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 16391 11522 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 16310 11522 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 16229 11522 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 16148 11522 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 16067 11522 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15986 11522 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15905 11522 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15824 11522 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15743 11522 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15662 11522 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15581 11522 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15500 11522 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15419 11522 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15338 11522 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15257 11522 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15176 11522 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15095 11522 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 15014 11522 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14933 11522 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14852 11522 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14771 11522 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14690 11522 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14609 11522 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14527 11522 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14445 11522 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14363 11522 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14281 11522 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14199 11522 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14117 11522 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 14035 11522 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 13953 11522 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 13871 11522 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 13789 11522 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 13707 11522 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11482 13625 11522 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 4432 11505 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 4346 11505 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 4260 11505 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 4174 11505 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 4088 11505 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 4002 11505 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 3916 11505 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 3830 11505 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 3744 11505 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 3658 11505 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11465 3572 11505 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11462 17575 11502 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11462 17494 11502 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11462 17413 11502 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11462 17332 11502 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11462 17251 11502 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11462 17171 11502 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11462 17091 11502 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11462 17011 11502 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11462 16931 11502 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11462 16851 11502 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11462 16771 11502 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11462 16691 11502 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11462 16611 11502 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 16472 11442 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 16391 11442 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 16310 11442 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 16229 11442 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 16148 11442 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 16067 11442 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15986 11442 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15905 11442 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15824 11442 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15743 11442 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15662 11442 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15581 11442 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15500 11442 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15419 11442 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15338 11442 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15257 11442 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15176 11442 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15095 11442 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 15014 11442 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14933 11442 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14852 11442 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14771 11442 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14690 11442 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14609 11442 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14527 11442 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14445 11442 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14363 11442 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14281 11442 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14199 11442 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14117 11442 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 14035 11442 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 13953 11442 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 13871 11442 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 13789 11442 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 13707 11442 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11402 13625 11442 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 4432 11424 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 4346 11424 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 4260 11424 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 4174 11424 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 4088 11424 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 4002 11424 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 3916 11424 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 3830 11424 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 3744 11424 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 3658 11424 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11384 3572 11424 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11380 17575 11420 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11380 17494 11420 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11380 17413 11420 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11380 17332 11420 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11380 17251 11420 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11380 17171 11420 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11380 17091 11420 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11380 17011 11420 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11380 16931 11420 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11380 16851 11420 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11380 16771 11420 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11380 16691 11420 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11380 16611 11420 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 16472 11362 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 16391 11362 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 16310 11362 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 16229 11362 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 16148 11362 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 16067 11362 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15986 11362 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15905 11362 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15824 11362 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15743 11362 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15662 11362 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15581 11362 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15500 11362 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15419 11362 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15338 11362 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15257 11362 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15176 11362 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15095 11362 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 15014 11362 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14933 11362 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14852 11362 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14771 11362 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14690 11362 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14609 11362 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14527 11362 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14445 11362 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14363 11362 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14281 11362 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14199 11362 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14117 11362 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 14035 11362 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 13953 11362 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 13871 11362 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 13789 11362 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 13707 11362 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11322 13625 11362 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 4432 11343 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 4346 11343 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 4260 11343 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 4174 11343 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 4088 11343 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 4002 11343 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 3916 11343 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 3830 11343 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 3744 11343 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 3658 11343 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11303 3572 11343 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11298 17575 11338 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11298 17494 11338 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11298 17413 11338 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11298 17332 11338 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11298 17251 11338 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11298 17171 11338 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11298 17091 11338 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11298 17011 11338 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11298 16931 11338 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11298 16851 11338 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11298 16771 11338 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11298 16691 11338 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11298 16611 11338 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 16472 11282 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 16391 11282 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 16310 11282 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 16229 11282 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 16148 11282 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 16067 11282 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15986 11282 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15905 11282 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15824 11282 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15743 11282 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15662 11282 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15581 11282 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15500 11282 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15419 11282 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15338 11282 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15257 11282 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15176 11282 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15095 11282 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 15014 11282 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14933 11282 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14852 11282 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14771 11282 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14690 11282 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14609 11282 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14527 11282 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14445 11282 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14363 11282 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14281 11282 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14199 11282 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14117 11282 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 14035 11282 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 13953 11282 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 13871 11282 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 13789 11282 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 13707 11282 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11242 13625 11282 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 4432 11262 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 4346 11262 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 4260 11262 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 4174 11262 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 4088 11262 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 4002 11262 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 3916 11262 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 3830 11262 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 3744 11262 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 3658 11262 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11222 3572 11262 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11199 17350 11239 17390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11199 17262 11239 17302 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11199 17175 11239 17215 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 16472 11202 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 16391 11202 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 16310 11202 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 16229 11202 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 16148 11202 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 16067 11202 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15986 11202 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15905 11202 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15824 11202 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15743 11202 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15662 11202 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15581 11202 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15500 11202 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15419 11202 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15338 11202 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15257 11202 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15176 11202 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15095 11202 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 15014 11202 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14933 11202 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14852 11202 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14771 11202 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14690 11202 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14609 11202 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14527 11202 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14445 11202 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14363 11202 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14281 11202 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14199 11202 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14117 11202 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 14035 11202 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 13953 11202 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 13871 11202 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 13789 11202 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 13707 11202 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11162 13625 11202 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11161 17065 11201 17105 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11161 16972 11201 17012 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11161 16879 11201 16919 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11161 16786 11201 16826 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11161 16694 11201 16734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11161 16602 11201 16642 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 4432 11181 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 4346 11181 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 4260 11181 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 4174 11181 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 4088 11181 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 4002 11181 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 3916 11181 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 3830 11181 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 3744 11181 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 3658 11181 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11141 3572 11181 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 16472 11122 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 16391 11122 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 16310 11122 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 16229 11122 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 16148 11122 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 16067 11122 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15986 11122 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15905 11122 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15824 11122 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15743 11122 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15662 11122 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15581 11122 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15500 11122 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15419 11122 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15338 11122 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15257 11122 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15176 11122 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15095 11122 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 15014 11122 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14933 11122 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14852 11122 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14771 11122 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14690 11122 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14609 11122 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14527 11122 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14445 11122 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14363 11122 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14281 11122 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14199 11122 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14117 11122 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 14035 11122 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 13953 11122 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 13871 11122 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 13789 11122 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 13707 11122 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11082 13625 11122 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11065 17065 11105 17105 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11065 16972 11105 17012 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11065 16879 11105 16919 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11065 16786 11105 16826 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11065 16694 11105 16734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11065 16602 11105 16642 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 4432 11100 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 4346 11100 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 4260 11100 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 4174 11100 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 4088 11100 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 4002 11100 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 3916 11100 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 3830 11100 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 3744 11100 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 3658 11100 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11060 3572 11100 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11051 17350 11091 17390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11051 17262 11091 17302 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11051 17175 11091 17215 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 16472 11042 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 16391 11042 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 16310 11042 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 16229 11042 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 16148 11042 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 16067 11042 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15986 11042 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15905 11042 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15824 11042 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15743 11042 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15662 11042 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15581 11042 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15500 11042 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15419 11042 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15338 11042 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15257 11042 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15176 11042 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15095 11042 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 15014 11042 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14933 11042 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14852 11042 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14771 11042 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14690 11042 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14609 11042 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14527 11042 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14445 11042 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14363 11042 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14281 11042 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14199 11042 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14117 11042 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 14035 11042 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 13953 11042 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 13871 11042 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 13789 11042 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 13707 11042 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 11002 13625 11042 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 4432 11019 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 4346 11019 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 4260 11019 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 4174 11019 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 4088 11019 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 4002 11019 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 3916 11019 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 3830 11019 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 3744 11019 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 3658 11019 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10979 3572 11019 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10969 17065 11009 17105 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10969 16972 11009 17012 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10969 16879 11009 16919 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10969 16786 11009 16826 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10969 16694 11009 16734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10969 16602 11009 16642 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 16472 10962 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 16391 10962 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 16310 10962 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 16229 10962 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 16148 10962 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 16067 10962 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15986 10962 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15905 10962 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15824 10962 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15743 10962 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15662 10962 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15581 10962 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15500 10962 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15419 10962 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15338 10962 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15257 10962 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15176 10962 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15095 10962 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 15014 10962 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14933 10962 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14852 10962 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14771 10962 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14690 10962 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14609 10962 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14527 10962 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14445 10962 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14363 10962 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14281 10962 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14199 10962 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14117 10962 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 14035 10962 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 13953 10962 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 13871 10962 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 13789 10962 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 13707 10962 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10922 13625 10962 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 4432 10938 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 4346 10938 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 4260 10938 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 4174 10938 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 4088 10938 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 4002 10938 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 3916 10938 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 3830 10938 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 3744 10938 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 3658 10938 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10898 3572 10938 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10873 17065 10913 17105 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10873 16972 10913 17012 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10873 16879 10913 16919 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10873 16786 10913 16826 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10873 16694 10913 16734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10873 16602 10913 16642 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 16472 10882 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 16391 10882 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 16310 10882 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 16229 10882 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 16148 10882 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 16067 10882 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15986 10882 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15905 10882 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15824 10882 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15743 10882 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15662 10882 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15581 10882 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15500 10882 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15419 10882 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15338 10882 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15257 10882 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15176 10882 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15095 10882 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 15014 10882 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14933 10882 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14852 10882 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14771 10882 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14690 10882 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14609 10882 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14527 10882 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14445 10882 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14363 10882 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14281 10882 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14199 10882 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14117 10882 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 14035 10882 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 13953 10882 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 13871 10882 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 13789 10882 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 13707 10882 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10842 13625 10882 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 4432 10857 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 4346 10857 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 4260 10857 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 4174 10857 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 4088 10857 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 4002 10857 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 3916 10857 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 3830 10857 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 3744 10857 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 3658 10857 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10817 3572 10857 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10777 17065 10817 17105 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10777 16972 10817 17012 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10777 16879 10817 16919 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10777 16786 10817 16826 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10777 16694 10817 16734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10777 16602 10817 16642 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 16472 10802 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 16391 10802 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 16310 10802 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 16229 10802 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 16148 10802 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 16067 10802 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15986 10802 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15905 10802 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15824 10802 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15743 10802 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15662 10802 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15581 10802 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15500 10802 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15419 10802 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15338 10802 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15257 10802 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15176 10802 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15095 10802 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 15014 10802 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14933 10802 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14852 10802 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14771 10802 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14690 10802 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14609 10802 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14527 10802 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14445 10802 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14363 10802 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14281 10802 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14199 10802 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14117 10802 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 14035 10802 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 13953 10802 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 13871 10802 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 13789 10802 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 13707 10802 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10762 13625 10802 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 4432 10776 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 4346 10776 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 4260 10776 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 4174 10776 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 4088 10776 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 4002 10776 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 3916 10776 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 3830 10776 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 3744 10776 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 3658 10776 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10736 3572 10776 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 16472 10722 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 16391 10722 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 16310 10722 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 16229 10722 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 16148 10722 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 16067 10722 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15986 10722 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15905 10722 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15824 10722 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15743 10722 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15662 10722 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15581 10722 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15500 10722 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15419 10722 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15338 10722 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15257 10722 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15176 10722 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15095 10722 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 15014 10722 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14933 10722 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14852 10722 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14771 10722 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14690 10722 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14609 10722 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14527 10722 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14445 10722 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14363 10722 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14281 10722 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14199 10722 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14117 10722 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 14035 10722 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 13953 10722 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 13871 10722 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 13789 10722 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 13707 10722 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10682 13625 10722 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10668 16804 10708 16844 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10668 16694 10708 16734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10668 16584 10708 16624 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 4432 10695 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 4346 10695 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 4260 10695 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 4174 10695 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 4088 10695 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 4002 10695 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 3916 10695 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 3830 10695 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 3744 10695 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 3658 10695 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10655 3572 10695 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 16472 10642 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 16391 10642 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 16310 10642 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 16229 10642 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 16148 10642 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 16067 10642 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15986 10642 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15905 10642 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15824 10642 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15743 10642 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15662 10642 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15581 10642 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15500 10642 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15419 10642 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15338 10642 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15257 10642 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15176 10642 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15095 10642 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 15014 10642 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14933 10642 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14852 10642 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14771 10642 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14690 10642 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14609 10642 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14527 10642 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14445 10642 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14363 10642 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14281 10642 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14199 10642 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14117 10642 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 14035 10642 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 13953 10642 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 13871 10642 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 13789 10642 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 13707 10642 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10602 13625 10642 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 4432 10614 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 4346 10614 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 4260 10614 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 4174 10614 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 4088 10614 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 4002 10614 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 3916 10614 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 3830 10614 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 3744 10614 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 3658 10614 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10574 3572 10614 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 16472 10562 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 16391 10562 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 16310 10562 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 16229 10562 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 16148 10562 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 16067 10562 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15986 10562 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15905 10562 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15824 10562 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15743 10562 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15662 10562 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15581 10562 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15500 10562 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15419 10562 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15338 10562 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15257 10562 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15176 10562 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15095 10562 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 15014 10562 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14933 10562 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14852 10562 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14771 10562 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14690 10562 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14609 10562 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14527 10562 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14445 10562 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14363 10562 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14281 10562 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14199 10562 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14117 10562 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 14035 10562 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 13953 10562 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 13871 10562 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 13789 10562 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 13707 10562 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10522 13625 10562 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 16804 10550 16844 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 16694 10550 16734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10510 16584 10550 16624 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 4432 10533 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 4346 10533 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 4260 10533 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 4174 10533 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 4088 10533 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 4002 10533 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 3916 10533 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 3830 10533 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 3744 10533 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 3658 10533 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10493 3572 10533 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 16472 10482 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 16391 10482 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 16310 10482 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 16229 10482 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 16148 10482 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 16067 10482 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15986 10482 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15905 10482 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15824 10482 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15743 10482 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15662 10482 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15581 10482 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15500 10482 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15419 10482 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15338 10482 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15257 10482 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15176 10482 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15095 10482 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 15014 10482 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14933 10482 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14852 10482 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14771 10482 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14690 10482 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14609 10482 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14527 10482 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14445 10482 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14363 10482 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14281 10482 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14199 10482 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14117 10482 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 14035 10482 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 13953 10482 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 13871 10482 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 13789 10482 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 13707 10482 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10442 13625 10482 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 4432 10452 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 4346 10452 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 4260 10452 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 4174 10452 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 4088 10452 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 4002 10452 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 3916 10452 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 3830 10452 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 3744 10452 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 3658 10452 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10412 3572 10452 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 16472 10402 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 16391 10402 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 16310 10402 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 16229 10402 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 16148 10402 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 16067 10402 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15986 10402 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15905 10402 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15824 10402 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15743 10402 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15662 10402 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15581 10402 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15500 10402 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15419 10402 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15338 10402 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15257 10402 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15176 10402 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15095 10402 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 15014 10402 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14933 10402 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14852 10402 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14771 10402 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14690 10402 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14609 10402 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14527 10402 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14445 10402 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14363 10402 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14281 10402 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14199 10402 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14117 10402 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 14035 10402 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 13953 10402 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 13871 10402 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 13789 10402 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 13707 10402 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10362 13625 10402 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 4432 10371 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 4346 10371 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 4260 10371 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 4174 10371 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 4088 10371 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 4002 10371 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 3916 10371 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 3830 10371 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 3744 10371 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 3658 10371 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10331 3572 10371 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 16472 10322 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 16391 10322 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 16310 10322 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 16229 10322 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 16148 10322 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 16067 10322 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15986 10322 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15905 10322 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15824 10322 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15743 10322 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15662 10322 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15581 10322 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15500 10322 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15419 10322 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15338 10322 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15257 10322 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15176 10322 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15095 10322 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 15014 10322 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14933 10322 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14852 10322 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14771 10322 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14690 10322 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14609 10322 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14527 10322 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14445 10322 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14363 10322 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14281 10322 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14199 10322 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14117 10322 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 14035 10322 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 13953 10322 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 13871 10322 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 13789 10322 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 13707 10322 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10282 13625 10322 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 4432 10290 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 4346 10290 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 4260 10290 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 4174 10290 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 4088 10290 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 4002 10290 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 3916 10290 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 3830 10290 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 3744 10290 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 3658 10290 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10250 3572 10290 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 16472 10242 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 16391 10242 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 16310 10242 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 16229 10242 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 16148 10242 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 16067 10242 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15986 10242 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15905 10242 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15824 10242 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15743 10242 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15662 10242 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15581 10242 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15500 10242 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15419 10242 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15338 10242 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15257 10242 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15176 10242 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15095 10242 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 15014 10242 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14933 10242 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14852 10242 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14771 10242 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14690 10242 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14609 10242 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14527 10242 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14445 10242 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14363 10242 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14281 10242 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14199 10242 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14117 10242 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 14035 10242 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 13953 10242 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 13871 10242 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 13789 10242 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 13707 10242 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10202 13625 10242 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 4432 10209 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 4346 10209 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 4260 10209 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 4174 10209 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 4088 10209 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 4002 10209 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 3916 10209 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 3830 10209 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 3744 10209 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 3658 10209 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 10169 3572 10209 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 4432 4882 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 4346 4882 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 4260 4882 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 4174 4882 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 4088 4882 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 4002 4882 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 3916 4882 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 3830 4882 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 3744 4882 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 3658 4882 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4842 3572 4882 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 16472 4849 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 16391 4849 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 16310 4849 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 16229 4849 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 16148 4849 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 16067 4849 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 15986 4849 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 15905 4849 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 15824 4849 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 15743 4849 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 15662 4849 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 15581 4849 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 15500 4849 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 15419 4849 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 15338 4849 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 15257 4849 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 15176 4849 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 15095 4849 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 15014 4849 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 14933 4849 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 14852 4849 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 14771 4849 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 14690 4849 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 14609 4849 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 14527 4849 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 14445 4849 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 14363 4849 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 14281 4849 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 14199 4849 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 14117 4849 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 14035 4849 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 13953 4849 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 13871 4849 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 13789 4849 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 13707 4849 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4809 13625 4849 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 4432 4800 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 4346 4800 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 4260 4800 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 4174 4800 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 4088 4800 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 4002 4800 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 3916 4800 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 3830 4800 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 3744 4800 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 3658 4800 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4760 3572 4800 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 16472 4769 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 16391 4769 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 16310 4769 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 16229 4769 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 16148 4769 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 16067 4769 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 15986 4769 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 15905 4769 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 15824 4769 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 15743 4769 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 15662 4769 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 15581 4769 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 15500 4769 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 15419 4769 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 15338 4769 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 15257 4769 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 15176 4769 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 15095 4769 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 15014 4769 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 14933 4769 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 14852 4769 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 14771 4769 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 14690 4769 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 14609 4769 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 14527 4769 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 14445 4769 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 14363 4769 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 14281 4769 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 14199 4769 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 14117 4769 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 14035 4769 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 13953 4769 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 13871 4769 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 13789 4769 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 13707 4769 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4729 13625 4769 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 4432 4718 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 4346 4718 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 4260 4718 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 4174 4718 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 4088 4718 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 4002 4718 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 3916 4718 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 3830 4718 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 3744 4718 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 3658 4718 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4678 3572 4718 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 16472 4689 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 16391 4689 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 16310 4689 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 16229 4689 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 16148 4689 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 16067 4689 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 15986 4689 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 15905 4689 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 15824 4689 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 15743 4689 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 15662 4689 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 15581 4689 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 15500 4689 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 15419 4689 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 15338 4689 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 15257 4689 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 15176 4689 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 15095 4689 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 15014 4689 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 14933 4689 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 14852 4689 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 14771 4689 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 14690 4689 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 14609 4689 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 14527 4689 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 14445 4689 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 14363 4689 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 14281 4689 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 14199 4689 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 14117 4689 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 14035 4689 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 13953 4689 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 13871 4689 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 13789 4689 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 13707 4689 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4649 13625 4689 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 4432 4636 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 4346 4636 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 4260 4636 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 4174 4636 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 4088 4636 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 4002 4636 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 3916 4636 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 3830 4636 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 3744 4636 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 3658 4636 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4596 3572 4636 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 16472 4609 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 16391 4609 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 16310 4609 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 16229 4609 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 16148 4609 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 16067 4609 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 15986 4609 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 15905 4609 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 15824 4609 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 15743 4609 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 15662 4609 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 15581 4609 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 15500 4609 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 15419 4609 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 15338 4609 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 15257 4609 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 15176 4609 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 15095 4609 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 15014 4609 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 14933 4609 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 14852 4609 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 14771 4609 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 14690 4609 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 14609 4609 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 14527 4609 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 14445 4609 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 14363 4609 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 14281 4609 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 14199 4609 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 14117 4609 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 14035 4609 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 13953 4609 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 13871 4609 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 13789 4609 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 13707 4609 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4569 13625 4609 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 4432 4554 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 4346 4554 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 4260 4554 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 4174 4554 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 4088 4554 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 4002 4554 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 3916 4554 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 3830 4554 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 3744 4554 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 3658 4554 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4514 3572 4554 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4501 16804 4541 16844 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4501 16694 4541 16734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4501 16584 4541 16624 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 16472 4529 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 16391 4529 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 16310 4529 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 16229 4529 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 16148 4529 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 16067 4529 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 15986 4529 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 15905 4529 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 15824 4529 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 15743 4529 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 15662 4529 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 15581 4529 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 15500 4529 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 15419 4529 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 15338 4529 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 15257 4529 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 15176 4529 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 15095 4529 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 15014 4529 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 14933 4529 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 14852 4529 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 14771 4529 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 14690 4529 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 14609 4529 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 14527 4529 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 14445 4529 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 14363 4529 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 14281 4529 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 14199 4529 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 14117 4529 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 14035 4529 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 13953 4529 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 13871 4529 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 13789 4529 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 13707 4529 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4489 13625 4529 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 4432 4472 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 4346 4472 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 4260 4472 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 4174 4472 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 4088 4472 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 4002 4472 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 3916 4472 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 3830 4472 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 3744 4472 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 3658 4472 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4432 3572 4472 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 16472 4449 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 16391 4449 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 16310 4449 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 16229 4449 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 16148 4449 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 16067 4449 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 15986 4449 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 15905 4449 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 15824 4449 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 15743 4449 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 15662 4449 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 15581 4449 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 15500 4449 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 15419 4449 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 15338 4449 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 15257 4449 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 15176 4449 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 15095 4449 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 15014 4449 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 14933 4449 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 14852 4449 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 14771 4449 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 14690 4449 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 14609 4449 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 14527 4449 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 14445 4449 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 14363 4449 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 14281 4449 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 14199 4449 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 14117 4449 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 14035 4449 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 13953 4449 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 13871 4449 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 13789 4449 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 13707 4449 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4409 13625 4449 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 4432 4390 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 4346 4390 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 4260 4390 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 4174 4390 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 4088 4390 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 4002 4390 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 3916 4390 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 3830 4390 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 3744 4390 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 3658 4390 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4350 3572 4390 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4343 16804 4383 16844 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4343 16694 4383 16734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4343 16584 4383 16624 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 16472 4369 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 16391 4369 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 16310 4369 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 16229 4369 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 16148 4369 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 16067 4369 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 15986 4369 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 15905 4369 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 15824 4369 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 15743 4369 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 15662 4369 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 15581 4369 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 15500 4369 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 15419 4369 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 15338 4369 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 15257 4369 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 15176 4369 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 15095 4369 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 15014 4369 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 14933 4369 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 14852 4369 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 14771 4369 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 14690 4369 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 14609 4369 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 14527 4369 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 14445 4369 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 14363 4369 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 14281 4369 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 14199 4369 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 14117 4369 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 14035 4369 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 13953 4369 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 13871 4369 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 13789 4369 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 13707 4369 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4329 13625 4369 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 4432 4309 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 4346 4309 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 4260 4309 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 4174 4309 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 4088 4309 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 4002 4309 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 3916 4309 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 3830 4309 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 3744 4309 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 3658 4309 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4269 3572 4309 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 16472 4289 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 16391 4289 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 16310 4289 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 16229 4289 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 16148 4289 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 16067 4289 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 15986 4289 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 15905 4289 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 15824 4289 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 15743 4289 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 15662 4289 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 15581 4289 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 15500 4289 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 15419 4289 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 15338 4289 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 15257 4289 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 15176 4289 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 15095 4289 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 15014 4289 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 14933 4289 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 14852 4289 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 14771 4289 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 14690 4289 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 14609 4289 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 14527 4289 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 14445 4289 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 14363 4289 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 14281 4289 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 14199 4289 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 14117 4289 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 14035 4289 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 13953 4289 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 13871 4289 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 13789 4289 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 13707 4289 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4249 13625 4289 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4234 17065 4274 17105 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4234 16972 4274 17012 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4234 16879 4274 16919 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4234 16786 4274 16826 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4234 16694 4274 16734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4234 16602 4274 16642 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 4432 4228 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 4346 4228 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 4260 4228 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 4174 4228 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 4088 4228 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 4002 4228 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 3916 4228 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 3830 4228 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 3744 4228 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 3658 4228 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4188 3572 4228 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 16472 4209 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 16391 4209 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 16310 4209 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 16229 4209 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 16148 4209 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 16067 4209 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 15986 4209 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 15905 4209 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 15824 4209 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 15743 4209 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 15662 4209 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 15581 4209 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 15500 4209 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 15419 4209 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 15338 4209 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 15257 4209 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 15176 4209 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 15095 4209 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 15014 4209 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 14933 4209 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 14852 4209 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 14771 4209 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 14690 4209 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 14609 4209 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 14527 4209 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 14445 4209 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 14363 4209 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 14281 4209 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 14199 4209 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 14117 4209 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 14035 4209 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 13953 4209 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 13871 4209 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 13789 4209 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 13707 4209 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4169 13625 4209 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4138 17065 4178 17105 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4138 16972 4178 17012 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4138 16879 4178 16919 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4138 16786 4178 16826 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4138 16694 4178 16734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4138 16602 4178 16642 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 4432 4147 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 4346 4147 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 4260 4147 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 4174 4147 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 4088 4147 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 4002 4147 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 3916 4147 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 3830 4147 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 3744 4147 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 3658 4147 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4107 3572 4147 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 16472 4129 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 16391 4129 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 16310 4129 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 16229 4129 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 16148 4129 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 16067 4129 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 15986 4129 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 15905 4129 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 15824 4129 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 15743 4129 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 15662 4129 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 15581 4129 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 15500 4129 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 15419 4129 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 15338 4129 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 15257 4129 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 15176 4129 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 15095 4129 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 15014 4129 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 14933 4129 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 14852 4129 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 14771 4129 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 14690 4129 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 14609 4129 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 14527 4129 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 14445 4129 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 14363 4129 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 14281 4129 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 14199 4129 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 14117 4129 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 14035 4129 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 13953 4129 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 13871 4129 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 13789 4129 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 13707 4129 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4089 13625 4129 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4042 17065 4082 17105 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4042 16972 4082 17012 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4042 16879 4082 16919 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4042 16786 4082 16826 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4042 16694 4082 16734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4042 16602 4082 16642 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 4432 4066 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 4346 4066 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 4260 4066 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 4174 4066 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 4088 4066 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 4002 4066 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 3916 4066 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 3830 4066 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 3744 4066 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 3658 4066 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4026 3572 4066 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 16472 4049 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 16391 4049 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 16310 4049 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 16229 4049 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 16148 4049 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 16067 4049 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 15986 4049 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 15905 4049 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 15824 4049 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 15743 4049 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 15662 4049 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 15581 4049 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 15500 4049 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 15419 4049 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 15338 4049 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 15257 4049 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 15176 4049 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 15095 4049 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 15014 4049 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 14933 4049 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 14852 4049 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 14771 4049 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 14690 4049 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 14609 4049 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 14527 4049 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 14445 4049 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 14363 4049 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 14281 4049 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 14199 4049 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 14117 4049 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 14035 4049 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 13953 4049 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 13871 4049 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 13789 4049 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 13707 4049 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 4009 13625 4049 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3960 17350 4000 17390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3960 17262 4000 17302 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3960 17175 4000 17215 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3946 17065 3986 17105 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3946 16972 3986 17012 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3946 16879 3986 16919 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3946 16786 3986 16826 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3946 16694 3986 16734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3946 16602 3986 16642 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 4432 3985 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 4346 3985 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 4260 3985 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 4174 3985 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 4088 3985 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 4002 3985 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 3916 3985 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 3830 3985 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 3744 3985 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 3658 3985 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3945 3572 3985 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 16472 3969 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 16391 3969 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 16310 3969 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 16229 3969 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 16148 3969 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 16067 3969 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 15986 3969 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 15905 3969 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 15824 3969 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 15743 3969 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 15662 3969 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 15581 3969 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 15500 3969 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 15419 3969 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 15338 3969 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 15257 3969 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 15176 3969 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 15095 3969 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 15014 3969 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 14933 3969 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 14852 3969 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 14771 3969 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 14690 3969 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 14609 3969 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 14527 3969 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 14445 3969 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 14363 3969 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 14281 3969 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 14199 3969 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 14117 3969 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 14035 3969 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 13953 3969 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 13871 3969 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 13789 3969 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 13707 3969 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3929 13625 3969 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 4432 3904 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 4346 3904 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 4260 3904 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 4174 3904 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 4088 3904 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 4002 3904 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 3916 3904 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 3830 3904 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 3744 3904 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 3658 3904 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3864 3572 3904 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3850 17065 3890 17105 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3850 16972 3890 17012 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3850 16879 3890 16919 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3850 16786 3890 16826 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3850 16694 3890 16734 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3850 16602 3890 16642 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 16472 3889 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 16391 3889 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 16310 3889 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 16229 3889 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 16148 3889 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 16067 3889 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 15986 3889 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 15905 3889 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 15824 3889 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 15743 3889 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 15662 3889 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 15581 3889 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 15500 3889 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 15419 3889 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 15338 3889 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 15257 3889 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 15176 3889 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 15095 3889 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 15014 3889 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 14933 3889 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 14852 3889 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 14771 3889 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 14690 3889 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 14609 3889 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 14527 3889 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 14445 3889 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 14363 3889 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 14281 3889 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 14199 3889 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 14117 3889 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 14035 3889 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 13953 3889 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 13871 3889 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 13789 3889 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 13707 3889 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3849 13625 3889 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3812 17350 3852 17390 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3812 17262 3852 17302 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3812 17175 3852 17215 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 4432 3823 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 4346 3823 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 4260 3823 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 4174 3823 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 4088 3823 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 4002 3823 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 3916 3823 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 3830 3823 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 3744 3823 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 3658 3823 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3783 3572 3823 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 16472 3809 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 16391 3809 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 16310 3809 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 16229 3809 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 16148 3809 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 16067 3809 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 15986 3809 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 15905 3809 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 15824 3809 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 15743 3809 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 15662 3809 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 15581 3809 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 15500 3809 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 15419 3809 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 15338 3809 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 15257 3809 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 15176 3809 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 15095 3809 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 15014 3809 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 14933 3809 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 14852 3809 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 14771 3809 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 14690 3809 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 14609 3809 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 14527 3809 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 14445 3809 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 14363 3809 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 14281 3809 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 14199 3809 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 14117 3809 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 14035 3809 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 13953 3809 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 13871 3809 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 13789 3809 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 13707 3809 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3769 13625 3809 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3713 17575 3753 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3713 17494 3753 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3713 17413 3753 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3713 17332 3753 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3713 17251 3753 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3713 17171 3753 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3713 17091 3753 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3713 17011 3753 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3713 16931 3753 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3713 16851 3753 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3713 16771 3753 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3713 16691 3753 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3713 16611 3753 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 4432 3742 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 4346 3742 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 4260 3742 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 4174 3742 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 4088 3742 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 4002 3742 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 3916 3742 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 3830 3742 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 3744 3742 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 3658 3742 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3702 3572 3742 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 16472 3729 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 16391 3729 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 16310 3729 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 16229 3729 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 16148 3729 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 16067 3729 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 15986 3729 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 15905 3729 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 15824 3729 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 15743 3729 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 15662 3729 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 15581 3729 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 15500 3729 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 15419 3729 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 15338 3729 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 15257 3729 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 15176 3729 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 15095 3729 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 15014 3729 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 14933 3729 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 14852 3729 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 14771 3729 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 14690 3729 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 14609 3729 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 14527 3729 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 14445 3729 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 14363 3729 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 14281 3729 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 14199 3729 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 14117 3729 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 14035 3729 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 13953 3729 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 13871 3729 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 13789 3729 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 13707 3729 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3689 13625 3729 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3631 17575 3671 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3631 17494 3671 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3631 17413 3671 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3631 17332 3671 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3631 17251 3671 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3631 17171 3671 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3631 17091 3671 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3631 17011 3671 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3631 16931 3671 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3631 16851 3671 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3631 16771 3671 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3631 16691 3671 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3631 16611 3671 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 4432 3661 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 4346 3661 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 4260 3661 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 4174 3661 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 4088 3661 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 4002 3661 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 3916 3661 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 3830 3661 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 3744 3661 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 3658 3661 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3621 3572 3661 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 16472 3649 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 16391 3649 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 16310 3649 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 16229 3649 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 16148 3649 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 16067 3649 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 15986 3649 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 15905 3649 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 15824 3649 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 15743 3649 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 15662 3649 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 15581 3649 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 15500 3649 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 15419 3649 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 15338 3649 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 15257 3649 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 15176 3649 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 15095 3649 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 15014 3649 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 14933 3649 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 14852 3649 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 14771 3649 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 14690 3649 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 14609 3649 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 14527 3649 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 14445 3649 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 14363 3649 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 14281 3649 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 14199 3649 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 14117 3649 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 14035 3649 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 13953 3649 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 13871 3649 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 13789 3649 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 13707 3649 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3609 13625 3649 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3549 17575 3589 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3549 17494 3589 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3549 17413 3589 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3549 17332 3589 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3549 17251 3589 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3549 17171 3589 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3549 17091 3589 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3549 17011 3589 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3549 16931 3589 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3549 16851 3589 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3549 16771 3589 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3549 16691 3589 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3549 16611 3589 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 4432 3580 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 4346 3580 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 4260 3580 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 4174 3580 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 4088 3580 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 4002 3580 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 3916 3580 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 3830 3580 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 3744 3580 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 3658 3580 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3540 3572 3580 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 16472 3569 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 16391 3569 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 16310 3569 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 16229 3569 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 16148 3569 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 16067 3569 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 15986 3569 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 15905 3569 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 15824 3569 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 15743 3569 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 15662 3569 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 15581 3569 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 15500 3569 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 15419 3569 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 15338 3569 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 15257 3569 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 15176 3569 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 15095 3569 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 15014 3569 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 14933 3569 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 14852 3569 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 14771 3569 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 14690 3569 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 14609 3569 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 14527 3569 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 14445 3569 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 14363 3569 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 14281 3569 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 14199 3569 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 14117 3569 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 14035 3569 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 13953 3569 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 13871 3569 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 13789 3569 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 13707 3569 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3529 13625 3569 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3467 17575 3507 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3467 17494 3507 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3467 17413 3507 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3467 17332 3507 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3467 17251 3507 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3467 17171 3507 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3467 17091 3507 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3467 17011 3507 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3467 16931 3507 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3467 16851 3507 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3467 16771 3507 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3467 16691 3507 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3467 16611 3507 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 4432 3499 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 4346 3499 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 4260 3499 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 4174 3499 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 4088 3499 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 4002 3499 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 3916 3499 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 3830 3499 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 3744 3499 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 3658 3499 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3459 3572 3499 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3452 17853 3492 17893 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3452 17769 3492 17809 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3452 17686 3492 17726 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 16472 3489 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 16391 3489 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 16310 3489 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 16229 3489 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 16148 3489 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 16067 3489 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 15986 3489 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 15905 3489 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 15824 3489 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 15743 3489 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 15662 3489 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 15581 3489 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 15500 3489 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 15419 3489 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 15338 3489 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 15257 3489 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 15176 3489 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 15095 3489 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 15014 3489 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 14933 3489 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 14852 3489 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 14771 3489 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 14690 3489 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 14609 3489 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 14527 3489 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 14445 3489 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 14363 3489 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 14281 3489 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 14199 3489 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 14117 3489 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 14035 3489 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 13953 3489 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 13871 3489 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 13789 3489 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 13707 3489 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3449 13625 3489 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3385 17575 3425 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3385 17494 3425 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3385 17413 3425 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3385 17332 3425 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3385 17251 3425 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3385 17171 3425 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3385 17091 3425 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3385 17011 3425 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3385 16931 3425 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3385 16851 3425 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3385 16771 3425 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3385 16691 3425 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3385 16611 3425 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 4432 3418 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 4346 3418 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 4260 3418 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 4174 3418 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 4088 3418 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 4002 3418 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 3916 3418 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 3830 3418 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 3744 3418 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 3658 3418 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3378 3572 3418 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 16472 3409 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 16391 3409 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 16310 3409 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 16229 3409 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 16148 3409 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 16067 3409 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 15986 3409 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 15905 3409 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 15824 3409 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 15743 3409 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 15662 3409 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 15581 3409 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 15500 3409 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 15419 3409 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 15338 3409 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 15257 3409 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 15176 3409 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 15095 3409 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 15014 3409 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 14933 3409 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 14852 3409 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 14771 3409 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 14690 3409 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 14609 3409 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 14527 3409 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 14445 3409 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 14363 3409 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 14281 3409 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 14199 3409 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 14117 3409 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 14035 3409 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 13953 3409 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 13871 3409 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 13789 3409 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 13707 3409 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3369 13625 3409 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3303 17575 3343 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3303 17494 3343 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3303 17413 3343 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3303 17332 3343 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3303 17251 3343 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3303 17171 3343 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3303 17091 3343 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3303 17011 3343 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3303 16931 3343 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3303 16851 3343 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3303 16771 3343 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3303 16691 3343 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3303 16611 3343 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 4432 3337 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 4346 3337 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 4260 3337 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 4174 3337 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 4088 3337 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 4002 3337 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 3916 3337 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 3830 3337 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 3744 3337 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 3658 3337 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3297 3572 3337 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3296 17853 3336 17893 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3296 17769 3336 17809 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3296 17686 3336 17726 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 16472 3329 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 16391 3329 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 16310 3329 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 16229 3329 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 16148 3329 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 16067 3329 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 15986 3329 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 15905 3329 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 15824 3329 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 15743 3329 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 15662 3329 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 15581 3329 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 15500 3329 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 15419 3329 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 15338 3329 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 15257 3329 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 15176 3329 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 15095 3329 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 15014 3329 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 14933 3329 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 14852 3329 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 14771 3329 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 14690 3329 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 14609 3329 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 14527 3329 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 14445 3329 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 14363 3329 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 14281 3329 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 14199 3329 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 14117 3329 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 14035 3329 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 13953 3329 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 13871 3329 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 13789 3329 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 13707 3329 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3289 13625 3329 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3221 17575 3261 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3221 17494 3261 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3221 17413 3261 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3221 17332 3261 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3221 17251 3261 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3221 17171 3261 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3221 17091 3261 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3221 17011 3261 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3221 16931 3261 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3221 16851 3261 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3221 16771 3261 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3221 16691 3261 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3221 16611 3261 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 4432 3256 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 4346 3256 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 4260 3256 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 4174 3256 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 4088 3256 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 4002 3256 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 3916 3256 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 3830 3256 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 3744 3256 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 3658 3256 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3216 3572 3256 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 16472 3249 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 16391 3249 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 16310 3249 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 16229 3249 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 16148 3249 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 16067 3249 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 15986 3249 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 15905 3249 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 15824 3249 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 15743 3249 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 15662 3249 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 15581 3249 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 15500 3249 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 15419 3249 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 15338 3249 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 15257 3249 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 15176 3249 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 15095 3249 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 15014 3249 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 14933 3249 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 14852 3249 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 14771 3249 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 14690 3249 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 14609 3249 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 14527 3249 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 14445 3249 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 14363 3249 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 14281 3249 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 14199 3249 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 14117 3249 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 14035 3249 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 13953 3249 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 13871 3249 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 13789 3249 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 13707 3249 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3209 13625 3249 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3196 18111 3236 18151 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3196 18025 3236 18065 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3196 17939 3236 17979 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3196 17853 3236 17893 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3196 17767 3236 17807 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3196 17682 3236 17722 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3139 17575 3179 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3139 17494 3179 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3139 17413 3179 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3139 17332 3179 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3139 17251 3179 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3139 17171 3179 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3139 17091 3179 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3139 17011 3179 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3139 16931 3179 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3139 16851 3179 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3139 16771 3179 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3139 16691 3179 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3139 16611 3179 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 4432 3175 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 4346 3175 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 4260 3175 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 4174 3175 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 4088 3175 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 4002 3175 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 3916 3175 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 3830 3175 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 3744 3175 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 3658 3175 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3135 3572 3175 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 16472 3169 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 16391 3169 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 16310 3169 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 16229 3169 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 16148 3169 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 16067 3169 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 15986 3169 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 15905 3169 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 15824 3169 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 15743 3169 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 15662 3169 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 15581 3169 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 15500 3169 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 15419 3169 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 15338 3169 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 15257 3169 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 15176 3169 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 15095 3169 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 15014 3169 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 14933 3169 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 14852 3169 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 14771 3169 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 14690 3169 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 14609 3169 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 14527 3169 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 14445 3169 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 14363 3169 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 14281 3169 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 14199 3169 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 14117 3169 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 14035 3169 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 13953 3169 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 13871 3169 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 13789 3169 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 13707 3169 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3129 13625 3169 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3114 18111 3154 18151 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3114 18025 3154 18065 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3114 17939 3154 17979 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3114 17853 3154 17893 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3114 17767 3154 17807 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3114 17682 3154 17722 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3057 17575 3097 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3057 17494 3097 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3057 17413 3097 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3057 17332 3097 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3057 17251 3097 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3057 17171 3097 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3057 17091 3097 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3057 17011 3097 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3057 16931 3097 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3057 16851 3097 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3057 16771 3097 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3057 16691 3097 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3057 16611 3097 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 4432 3094 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 4346 3094 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 4260 3094 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 4174 3094 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 4088 3094 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 4002 3094 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 3916 3094 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 3830 3094 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 3744 3094 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 3658 3094 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3054 3572 3094 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 16472 3089 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 16391 3089 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 16310 3089 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 16229 3089 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 16148 3089 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 16067 3089 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 15986 3089 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 15905 3089 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 15824 3089 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 15743 3089 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 15662 3089 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 15581 3089 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 15500 3089 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 15419 3089 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 15338 3089 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 15257 3089 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 15176 3089 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 15095 3089 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 15014 3089 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 14933 3089 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 14852 3089 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 14771 3089 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 14690 3089 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 14609 3089 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 14527 3089 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 14445 3089 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 14363 3089 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 14281 3089 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 14199 3089 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 14117 3089 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 14035 3089 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 13953 3089 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 13871 3089 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 13789 3089 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 13707 3089 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3049 13625 3089 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3032 18111 3072 18151 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3032 18025 3072 18065 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3032 17939 3072 17979 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3032 17853 3072 17893 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3032 17767 3072 17807 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3032 17682 3072 17722 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3020 18289 3060 18329 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 3020 18203 3060 18243 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2975 17575 3015 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2975 17494 3015 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2975 17413 3015 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2975 17332 3015 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2975 17251 3015 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2975 17171 3015 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2975 17091 3015 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2975 17011 3015 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2975 16931 3015 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2975 16851 3015 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2975 16771 3015 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2975 16691 3015 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2975 16611 3015 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 4432 3013 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 4346 3013 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 4260 3013 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 4174 3013 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 4088 3013 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 4002 3013 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 3916 3013 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 3830 3013 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 3744 3013 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 3658 3013 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2973 3572 3013 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 16472 3009 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 16391 3009 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 16310 3009 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 16229 3009 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 16148 3009 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 16067 3009 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 15986 3009 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 15905 3009 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 15824 3009 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 15743 3009 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 15662 3009 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 15581 3009 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 15500 3009 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 15419 3009 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 15338 3009 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 15257 3009 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 15176 3009 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 15095 3009 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 15014 3009 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 14933 3009 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 14852 3009 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 14771 3009 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 14690 3009 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 14609 3009 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 14527 3009 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 14445 3009 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 14363 3009 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 14281 3009 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 14199 3009 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 14117 3009 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 14035 3009 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 13953 3009 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 13871 3009 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 13789 3009 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 13707 3009 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2969 13625 3009 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2950 18111 2990 18151 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2950 18025 2990 18065 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2950 17939 2990 17979 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2950 17853 2990 17893 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2950 17767 2990 17807 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2950 17682 2990 17722 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2893 17575 2933 17615 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2893 17494 2933 17534 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2893 17413 2933 17453 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2893 17332 2933 17372 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2893 17251 2933 17291 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2893 17171 2933 17211 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2893 17091 2933 17131 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2893 17011 2933 17051 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2893 16931 2933 16971 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2893 16851 2933 16891 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2893 16771 2933 16811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2893 16691 2933 16731 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2893 16611 2933 16651 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 4432 2932 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 4346 2932 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 4260 2932 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 4174 2932 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 4088 2932 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 4002 2932 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 3916 2932 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 3830 2932 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 3744 2932 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 3658 2932 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2892 3572 2932 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 16472 2929 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 16391 2929 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 16310 2929 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 16229 2929 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 16148 2929 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 16067 2929 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 15986 2929 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 15905 2929 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 15824 2929 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 15743 2929 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 15662 2929 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 15581 2929 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 15500 2929 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 15419 2929 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 15338 2929 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 15257 2929 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 15176 2929 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 15095 2929 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 15014 2929 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 14933 2929 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 14852 2929 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 14771 2929 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 14690 2929 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 14609 2929 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 14527 2929 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 14445 2929 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 14363 2929 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 14281 2929 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 14199 2929 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 14117 2929 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 14035 2929 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 13953 2929 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 13871 2929 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 13789 2929 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 13707 2929 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2889 13625 2929 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2868 18111 2908 18151 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2868 18025 2908 18065 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2868 17939 2908 17979 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2868 17853 2908 17893 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2868 17767 2908 17807 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2868 17682 2908 17722 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2864 18289 2904 18329 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2864 18203 2904 18243 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 4432 2851 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 4346 2851 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 4260 2851 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 4174 2851 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 4088 2851 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 4002 2851 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 3916 2851 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 3830 2851 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 3744 2851 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 3658 2851 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2811 3572 2851 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 16472 2849 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 16391 2849 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 16310 2849 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 16229 2849 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 16148 2849 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 16067 2849 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 15986 2849 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 15905 2849 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 15824 2849 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 15743 2849 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 15662 2849 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 15581 2849 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 15500 2849 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 15419 2849 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 15338 2849 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 15257 2849 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 15176 2849 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 15095 2849 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 15014 2849 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 14933 2849 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 14852 2849 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 14771 2849 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 14690 2849 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 14609 2849 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 14527 2849 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 14445 2849 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 14363 2849 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 14281 2849 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 14199 2849 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 14117 2849 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 14035 2849 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 13953 2849 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 13871 2849 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 13789 2849 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 13707 2849 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2809 13625 2849 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2768 18539 2808 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2768 18457 2808 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2768 18375 2808 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2768 18293 2808 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2768 18211 2808 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2768 18129 2808 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2768 18047 2808 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2768 17965 2808 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2768 17883 2808 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2768 17801 2808 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2768 17719 2808 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2768 17637 2808 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2768 17555 2808 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2768 17473 2808 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2768 17391 2808 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2768 17309 2808 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2768 17227 2808 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2768 17145 2808 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2768 17063 2808 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2768 16981 2808 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2768 16899 2808 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2768 16817 2808 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2768 16735 2808 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2768 16653 2808 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2768 16571 2808 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 4432 2770 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 4346 2770 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 4260 2770 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 4174 2770 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 4088 2770 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 4002 2770 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 3916 2770 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 3830 2770 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 3744 2770 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 3658 2770 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2730 3572 2770 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 16472 2769 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 16391 2769 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 16310 2769 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 16229 2769 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 16148 2769 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 16067 2769 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 15986 2769 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 15905 2769 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 15824 2769 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 15743 2769 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 15662 2769 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 15581 2769 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 15500 2769 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 15419 2769 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 15338 2769 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 15257 2769 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 15176 2769 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 15095 2769 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 15014 2769 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 14933 2769 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 14852 2769 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 14771 2769 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 14690 2769 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 14609 2769 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 14527 2769 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 14445 2769 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 14363 2769 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 14281 2769 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 14199 2769 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 14117 2769 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 14035 2769 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 13953 2769 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 13871 2769 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 13789 2769 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 13707 2769 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2729 13625 2769 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2687 18539 2727 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2687 18457 2727 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2687 18375 2727 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2687 18293 2727 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2687 18211 2727 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2687 18129 2727 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2687 18047 2727 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2687 17965 2727 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2687 17883 2727 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2687 17801 2727 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2687 17719 2727 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2687 17637 2727 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2687 17555 2727 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2687 17473 2727 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2687 17391 2727 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2687 17309 2727 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2687 17227 2727 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2687 17145 2727 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2687 17063 2727 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2687 16981 2727 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2687 16899 2727 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2687 16817 2727 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2687 16735 2727 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2687 16653 2727 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2687 16571 2727 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 16472 2689 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 16391 2689 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 16310 2689 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 16229 2689 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 16148 2689 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 16067 2689 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 15986 2689 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 15905 2689 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 15824 2689 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 15743 2689 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 15662 2689 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 15581 2689 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 15500 2689 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 15419 2689 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 15338 2689 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 15257 2689 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 15176 2689 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 15095 2689 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 15014 2689 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 14933 2689 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 14852 2689 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 14771 2689 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 14690 2689 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 14609 2689 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 14527 2689 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 14445 2689 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 14363 2689 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 14281 2689 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 14199 2689 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 14117 2689 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 14035 2689 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 13953 2689 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 13871 2689 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 13789 2689 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 13707 2689 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 13625 2689 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 4432 2689 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 4346 2689 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 4260 2689 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 4174 2689 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 4088 2689 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 4002 2689 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 3916 2689 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 3830 2689 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 3744 2689 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 3658 2689 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2649 3572 2689 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2606 18539 2646 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2606 18457 2646 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2606 18375 2646 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2606 18293 2646 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2606 18211 2646 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2606 18129 2646 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2606 18047 2646 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2606 17965 2646 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2606 17883 2646 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2606 17801 2646 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2606 17719 2646 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2606 17637 2646 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2606 17555 2646 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2606 17473 2646 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2606 17391 2646 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2606 17309 2646 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2606 17227 2646 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2606 17145 2646 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2606 17063 2646 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2606 16981 2646 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2606 16899 2646 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2606 16817 2646 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2606 16735 2646 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2606 16653 2646 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2606 16571 2646 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 16472 2609 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 16391 2609 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 16310 2609 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 16229 2609 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 16148 2609 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 16067 2609 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 15986 2609 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 15905 2609 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 15824 2609 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 15743 2609 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 15662 2609 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 15581 2609 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 15500 2609 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 15419 2609 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 15338 2609 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 15257 2609 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 15176 2609 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 15095 2609 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 15014 2609 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 14933 2609 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 14852 2609 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 14771 2609 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 14690 2609 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 14609 2609 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 14527 2609 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 14445 2609 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 14363 2609 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 14281 2609 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 14199 2609 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 14117 2609 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 14035 2609 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 13953 2609 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 13871 2609 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 13789 2609 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 13707 2609 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2569 13625 2609 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 4432 2608 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 4346 2608 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 4260 2608 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 4174 2608 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 4088 2608 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 4002 2608 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 3916 2608 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 3830 2608 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 3744 2608 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 3658 2608 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2568 3572 2608 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2525 18539 2565 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2525 18457 2565 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2525 18375 2565 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2525 18293 2565 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2525 18211 2565 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2525 18129 2565 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2525 18047 2565 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2525 17965 2565 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2525 17883 2565 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2525 17801 2565 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2525 17719 2565 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2525 17637 2565 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2525 17555 2565 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2525 17473 2565 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2525 17391 2565 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2525 17309 2565 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2525 17227 2565 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2525 17145 2565 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2525 17063 2565 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2525 16981 2565 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2525 16899 2565 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2525 16817 2565 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2525 16735 2565 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2525 16653 2565 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2525 16571 2565 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 16472 2529 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 16391 2529 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 16310 2529 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 16229 2529 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 16148 2529 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 16067 2529 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 15986 2529 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 15905 2529 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 15824 2529 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 15743 2529 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 15662 2529 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 15581 2529 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 15500 2529 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 15419 2529 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 15338 2529 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 15257 2529 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 15176 2529 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 15095 2529 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 15014 2529 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 14933 2529 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 14852 2529 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 14771 2529 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 14690 2529 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 14609 2529 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 14527 2529 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 14445 2529 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 14363 2529 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 14281 2529 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 14199 2529 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 14117 2529 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 14035 2529 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 13953 2529 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 13871 2529 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 13789 2529 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 13707 2529 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2489 13625 2529 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 4432 2527 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 4346 2527 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 4260 2527 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 4174 2527 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 4088 2527 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 4002 2527 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 3916 2527 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 3830 2527 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 3744 2527 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 3658 2527 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2487 3572 2527 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2443 18539 2483 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2443 18457 2483 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2443 18375 2483 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2443 18293 2483 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2443 18211 2483 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2443 18129 2483 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2443 18047 2483 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2443 17965 2483 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2443 17883 2483 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2443 17801 2483 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2443 17719 2483 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2443 17637 2483 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2443 17555 2483 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2443 17473 2483 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2443 17391 2483 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2443 17309 2483 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2443 17227 2483 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2443 17145 2483 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2443 17063 2483 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2443 16981 2483 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2443 16899 2483 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2443 16817 2483 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2443 16735 2483 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2443 16653 2483 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2443 16571 2483 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 16472 2449 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 16391 2449 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 16310 2449 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 16229 2449 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 16148 2449 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 16067 2449 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 15986 2449 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 15905 2449 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 15824 2449 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 15743 2449 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 15662 2449 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 15581 2449 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 15500 2449 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 15419 2449 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 15338 2449 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 15257 2449 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 15176 2449 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 15095 2449 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 15014 2449 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 14933 2449 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 14852 2449 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 14771 2449 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 14690 2449 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 14609 2449 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 14527 2449 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 14445 2449 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 14363 2449 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 14281 2449 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 14199 2449 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 14117 2449 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 14035 2449 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 13953 2449 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 13871 2449 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 13789 2449 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 13707 2449 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2409 13625 2449 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 4432 2446 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 4346 2446 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 4260 2446 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 4174 2446 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 4088 2446 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 4002 2446 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 3916 2446 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 3830 2446 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 3744 2446 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 3658 2446 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2406 3572 2446 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2361 18539 2401 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2361 18457 2401 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2361 18375 2401 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2361 18293 2401 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2361 18211 2401 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2361 18129 2401 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2361 18047 2401 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2361 17965 2401 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2361 17883 2401 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2361 17801 2401 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2361 17719 2401 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2361 17637 2401 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2361 17555 2401 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2361 17473 2401 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2361 17391 2401 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2361 17309 2401 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2361 17227 2401 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2361 17145 2401 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2361 17063 2401 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2361 16981 2401 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2361 16899 2401 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2361 16817 2401 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2361 16735 2401 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2361 16653 2401 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2361 16571 2401 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 16472 2369 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 16391 2369 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 16310 2369 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 16229 2369 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 16148 2369 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 16067 2369 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 15986 2369 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 15905 2369 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 15824 2369 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 15743 2369 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 15662 2369 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 15581 2369 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 15500 2369 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 15419 2369 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 15338 2369 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 15257 2369 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 15176 2369 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 15095 2369 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 15014 2369 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 14933 2369 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 14852 2369 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 14771 2369 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 14690 2369 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 14609 2369 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 14527 2369 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 14445 2369 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 14363 2369 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 14281 2369 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 14199 2369 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 14117 2369 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 14035 2369 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 13953 2369 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 13871 2369 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 13789 2369 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 13707 2369 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2329 13625 2369 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 4432 2365 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 4346 2365 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 4260 2365 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 4174 2365 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 4088 2365 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 4002 2365 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 3916 2365 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 3830 2365 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 3744 2365 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 3658 2365 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2325 3572 2365 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2279 18539 2319 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2279 18457 2319 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2279 18375 2319 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2279 18293 2319 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2279 18211 2319 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2279 18129 2319 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2279 18047 2319 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2279 17965 2319 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2279 17883 2319 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2279 17801 2319 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2279 17719 2319 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2279 17637 2319 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2279 17555 2319 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2279 17473 2319 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2279 17391 2319 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2279 17309 2319 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2279 17227 2319 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2279 17145 2319 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2279 17063 2319 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2279 16981 2319 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2279 16899 2319 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2279 16817 2319 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2279 16735 2319 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2279 16653 2319 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2279 16571 2319 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 16472 2289 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 16391 2289 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 16310 2289 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 16229 2289 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 16148 2289 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 16067 2289 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 15986 2289 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 15905 2289 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 15824 2289 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 15743 2289 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 15662 2289 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 15581 2289 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 15500 2289 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 15419 2289 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 15338 2289 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 15257 2289 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 15176 2289 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 15095 2289 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 15014 2289 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 14933 2289 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 14852 2289 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 14771 2289 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 14690 2289 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 14609 2289 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 14527 2289 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 14445 2289 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 14363 2289 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 14281 2289 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 14199 2289 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 14117 2289 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 14035 2289 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 13953 2289 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 13871 2289 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 13789 2289 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 13707 2289 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2249 13625 2289 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 4432 2284 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 4346 2284 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 4260 2284 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 4174 2284 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 4088 2284 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 4002 2284 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 3916 2284 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 3830 2284 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 3744 2284 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 3658 2284 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2244 3572 2284 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2197 18539 2237 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2197 18457 2237 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2197 18375 2237 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2197 18293 2237 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2197 18211 2237 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2197 18129 2237 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2197 18047 2237 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2197 17965 2237 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2197 17883 2237 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2197 17801 2237 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2197 17719 2237 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2197 17637 2237 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2197 17555 2237 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2197 17473 2237 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2197 17391 2237 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2197 17309 2237 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2197 17227 2237 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2197 17145 2237 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2197 17063 2237 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2197 16981 2237 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2197 16899 2237 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2197 16817 2237 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2197 16735 2237 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2197 16653 2237 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2197 16571 2237 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 16472 2209 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 16391 2209 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 16310 2209 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 16229 2209 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 16148 2209 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 16067 2209 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 15986 2209 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 15905 2209 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 15824 2209 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 15743 2209 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 15662 2209 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 15581 2209 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 15500 2209 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 15419 2209 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 15338 2209 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 15257 2209 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 15176 2209 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 15095 2209 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 15014 2209 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 14933 2209 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 14852 2209 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 14771 2209 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 14690 2209 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 14609 2209 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 14527 2209 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 14445 2209 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 14363 2209 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 14281 2209 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 14199 2209 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 14117 2209 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 14035 2209 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 13953 2209 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 13871 2209 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 13789 2209 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 13707 2209 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2169 13625 2209 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 4432 2203 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 4346 2203 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 4260 2203 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 4174 2203 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 4088 2203 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 4002 2203 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 3916 2203 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 3830 2203 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 3744 2203 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 3658 2203 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2163 3572 2203 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2115 18539 2155 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2115 18457 2155 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2115 18375 2155 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2115 18293 2155 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2115 18211 2155 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2115 18129 2155 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2115 18047 2155 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2115 17965 2155 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2115 17883 2155 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2115 17801 2155 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2115 17719 2155 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2115 17637 2155 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2115 17555 2155 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2115 17473 2155 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2115 17391 2155 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2115 17309 2155 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2115 17227 2155 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2115 17145 2155 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2115 17063 2155 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2115 16981 2155 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2115 16899 2155 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2115 16817 2155 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2115 16735 2155 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2115 16653 2155 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2115 16571 2155 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 16472 2129 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 16391 2129 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 16310 2129 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 16229 2129 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 16148 2129 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 16067 2129 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 15986 2129 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 15905 2129 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 15824 2129 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 15743 2129 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 15662 2129 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 15581 2129 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 15500 2129 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 15419 2129 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 15338 2129 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 15257 2129 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 15176 2129 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 15095 2129 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 15014 2129 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 14933 2129 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 14852 2129 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 14771 2129 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 14690 2129 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 14609 2129 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 14527 2129 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 14445 2129 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 14363 2129 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 14281 2129 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 14199 2129 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 14117 2129 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 14035 2129 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 13953 2129 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 13871 2129 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 13789 2129 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 13707 2129 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2089 13625 2129 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 4432 2122 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 4346 2122 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 4260 2122 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 4174 2122 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 4088 2122 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 4002 2122 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 3916 2122 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 3830 2122 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 3744 2122 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 3658 2122 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2082 3572 2122 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2033 18539 2073 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2033 18457 2073 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2033 18375 2073 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2033 18293 2073 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2033 18211 2073 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2033 18129 2073 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2033 18047 2073 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2033 17965 2073 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2033 17883 2073 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2033 17801 2073 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2033 17719 2073 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2033 17637 2073 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2033 17555 2073 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2033 17473 2073 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2033 17391 2073 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2033 17309 2073 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2033 17227 2073 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2033 17145 2073 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2033 17063 2073 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2033 16981 2073 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2033 16899 2073 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2033 16817 2073 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2033 16735 2073 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2033 16653 2073 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2033 16571 2073 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 16472 2049 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 16391 2049 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 16310 2049 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 16229 2049 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 16148 2049 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 16067 2049 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 15986 2049 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 15905 2049 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 15824 2049 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 15743 2049 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 15662 2049 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 15581 2049 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 15500 2049 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 15419 2049 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 15338 2049 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 15257 2049 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 15176 2049 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 15095 2049 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 15014 2049 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 14933 2049 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 14852 2049 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 14771 2049 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 14690 2049 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 14609 2049 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 14527 2049 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 14445 2049 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 14363 2049 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 14281 2049 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 14199 2049 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 14117 2049 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 14035 2049 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 13953 2049 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 13871 2049 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 13789 2049 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 13707 2049 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2009 13625 2049 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 4432 2041 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 4346 2041 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 4260 2041 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 4174 2041 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 4088 2041 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 4002 2041 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 3916 2041 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 3830 2041 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 3744 2041 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 3658 2041 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 2001 3572 2041 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1951 18539 1991 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1951 18457 1991 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1951 18375 1991 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1951 18293 1991 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1951 18211 1991 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1951 18129 1991 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1951 18047 1991 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1951 17965 1991 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1951 17883 1991 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1951 17801 1991 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1951 17719 1991 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1951 17637 1991 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1951 17555 1991 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1951 17473 1991 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1951 17391 1991 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1951 17309 1991 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1951 17227 1991 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1951 17145 1991 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1951 17063 1991 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1951 16981 1991 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1951 16899 1991 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1951 16817 1991 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1951 16735 1991 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1951 16653 1991 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1951 16571 1991 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 16472 1969 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 16391 1969 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 16310 1969 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 16229 1969 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 16148 1969 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 16067 1969 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 15986 1969 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 15905 1969 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 15824 1969 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 15743 1969 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 15662 1969 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 15581 1969 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 15500 1969 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 15419 1969 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 15338 1969 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 15257 1969 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 15176 1969 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 15095 1969 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 15014 1969 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 14933 1969 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 14852 1969 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 14771 1969 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 14690 1969 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 14609 1969 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 14527 1969 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 14445 1969 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 14363 1969 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 14281 1969 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 14199 1969 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 14117 1969 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 14035 1969 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 13953 1969 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 13871 1969 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 13789 1969 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 13707 1969 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1929 13625 1969 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 4432 1960 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 4346 1960 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 4260 1960 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 4174 1960 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 4088 1960 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 4002 1960 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 3916 1960 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 3830 1960 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 3744 1960 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 3658 1960 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1920 3572 1960 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1869 18539 1909 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1869 18457 1909 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1869 18375 1909 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1869 18293 1909 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1869 18211 1909 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1869 18129 1909 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1869 18047 1909 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1869 17965 1909 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1869 17883 1909 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1869 17801 1909 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1869 17719 1909 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1869 17637 1909 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1869 17555 1909 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1869 17473 1909 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1869 17391 1909 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1869 17309 1909 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1869 17227 1909 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1869 17145 1909 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1869 17063 1909 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1869 16981 1909 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1869 16899 1909 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1869 16817 1909 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1869 16735 1909 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1869 16653 1909 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1869 16571 1909 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 16472 1889 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 16391 1889 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 16310 1889 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 16229 1889 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 16148 1889 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 16067 1889 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 15986 1889 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 15905 1889 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 15824 1889 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 15743 1889 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 15662 1889 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 15581 1889 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 15500 1889 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 15419 1889 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 15338 1889 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 15257 1889 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 15176 1889 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 15095 1889 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 15014 1889 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 14933 1889 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 14852 1889 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 14771 1889 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 14690 1889 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 14609 1889 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 14527 1889 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 14445 1889 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 14363 1889 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 14281 1889 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 14199 1889 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 14117 1889 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 14035 1889 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 13953 1889 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 13871 1889 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 13789 1889 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 13707 1889 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1849 13625 1889 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 4432 1879 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 4346 1879 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 4260 1879 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 4174 1879 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 4088 1879 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 4002 1879 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 3916 1879 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 3830 1879 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 3744 1879 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 3658 1879 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1839 3572 1879 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1787 18539 1827 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1787 18457 1827 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1787 18375 1827 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1787 18293 1827 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1787 18211 1827 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1787 18129 1827 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1787 18047 1827 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1787 17965 1827 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1787 17883 1827 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1787 17801 1827 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1787 17719 1827 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1787 17637 1827 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1787 17555 1827 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1787 17473 1827 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1787 17391 1827 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1787 17309 1827 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1787 17227 1827 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1787 17145 1827 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1787 17063 1827 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1787 16981 1827 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1787 16899 1827 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1787 16817 1827 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1787 16735 1827 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1787 16653 1827 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1787 16571 1827 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 16472 1809 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 16391 1809 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 16310 1809 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 16229 1809 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 16148 1809 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 16067 1809 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 15986 1809 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 15905 1809 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 15824 1809 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 15743 1809 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 15662 1809 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 15581 1809 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 15500 1809 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 15419 1809 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 15338 1809 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 15257 1809 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 15176 1809 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 15095 1809 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 15014 1809 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 14933 1809 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 14852 1809 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 14771 1809 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 14690 1809 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 14609 1809 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 14527 1809 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 14445 1809 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 14363 1809 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 14281 1809 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 14199 1809 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 14117 1809 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 14035 1809 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 13953 1809 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 13871 1809 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 13789 1809 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 13707 1809 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1769 13625 1809 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 4432 1798 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 4346 1798 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 4260 1798 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 4174 1798 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 4088 1798 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 4002 1798 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 3916 1798 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 3830 1798 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 3744 1798 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 3658 1798 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1758 3572 1798 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1705 18539 1745 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1705 18457 1745 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1705 18375 1745 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1705 18293 1745 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1705 18211 1745 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1705 18129 1745 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1705 18047 1745 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1705 17965 1745 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1705 17883 1745 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1705 17801 1745 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1705 17719 1745 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1705 17637 1745 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1705 17555 1745 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1705 17473 1745 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1705 17391 1745 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1705 17309 1745 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1705 17227 1745 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1705 17145 1745 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1705 17063 1745 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1705 16981 1745 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1705 16899 1745 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1705 16817 1745 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1705 16735 1745 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1705 16653 1745 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1705 16571 1745 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 16472 1729 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 16391 1729 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 16310 1729 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 16229 1729 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 16148 1729 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 16067 1729 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 15986 1729 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 15905 1729 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 15824 1729 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 15743 1729 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 15662 1729 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 15581 1729 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 15500 1729 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 15419 1729 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 15338 1729 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 15257 1729 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 15176 1729 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 15095 1729 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 15014 1729 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 14933 1729 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 14852 1729 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 14771 1729 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 14690 1729 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 14609 1729 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 14527 1729 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 14445 1729 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 14363 1729 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 14281 1729 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 14199 1729 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 14117 1729 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 14035 1729 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 13953 1729 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 13871 1729 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 13789 1729 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 13707 1729 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1689 13625 1729 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 4432 1717 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 4346 1717 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 4260 1717 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 4174 1717 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 4088 1717 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 4002 1717 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 3916 1717 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 3830 1717 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 3744 1717 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 3658 1717 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1677 3572 1717 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1623 18539 1663 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1623 18457 1663 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1623 18375 1663 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1623 18293 1663 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1623 18211 1663 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1623 18129 1663 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1623 18047 1663 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1623 17965 1663 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1623 17883 1663 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1623 17801 1663 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1623 17719 1663 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1623 17637 1663 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1623 17555 1663 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1623 17473 1663 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1623 17391 1663 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1623 17309 1663 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1623 17227 1663 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1623 17145 1663 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1623 17063 1663 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1623 16981 1663 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1623 16899 1663 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1623 16817 1663 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1623 16735 1663 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1623 16653 1663 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1623 16571 1663 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 16472 1649 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 16391 1649 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 16310 1649 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 16229 1649 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 16148 1649 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 16067 1649 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 15986 1649 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 15905 1649 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 15824 1649 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 15743 1649 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 15662 1649 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 15581 1649 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 15500 1649 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 15419 1649 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 15338 1649 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 15257 1649 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 15176 1649 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 15095 1649 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 15014 1649 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 14933 1649 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 14852 1649 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 14771 1649 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 14690 1649 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 14609 1649 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 14527 1649 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 14445 1649 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 14363 1649 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 14281 1649 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 14199 1649 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 14117 1649 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 14035 1649 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 13953 1649 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 13871 1649 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 13789 1649 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 13707 1649 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1609 13625 1649 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 4432 1636 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 4346 1636 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 4260 1636 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 4174 1636 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 4088 1636 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 4002 1636 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 3916 1636 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 3830 1636 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 3744 1636 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 3658 1636 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1596 3572 1636 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1541 18539 1581 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1541 18457 1581 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1541 18375 1581 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1541 18293 1581 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1541 18211 1581 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1541 18129 1581 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1541 18047 1581 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1541 17965 1581 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1541 17883 1581 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1541 17801 1581 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1541 17719 1581 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1541 17637 1581 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1541 17555 1581 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1541 17473 1581 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1541 17391 1581 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1541 17309 1581 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1541 17227 1581 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1541 17145 1581 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1541 17063 1581 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1541 16981 1581 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1541 16899 1581 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1541 16817 1581 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1541 16735 1581 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1541 16653 1581 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1541 16571 1581 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 16472 1569 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 16391 1569 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 16310 1569 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 16229 1569 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 16148 1569 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 16067 1569 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 15986 1569 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 15905 1569 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 15824 1569 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 15743 1569 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 15662 1569 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 15581 1569 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 15500 1569 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 15419 1569 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 15338 1569 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 15257 1569 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 15176 1569 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 15095 1569 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 15014 1569 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 14933 1569 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 14852 1569 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 14771 1569 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 14690 1569 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 14609 1569 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 14527 1569 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 14445 1569 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 14363 1569 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 14281 1569 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 14199 1569 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 14117 1569 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 14035 1569 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 13953 1569 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 13871 1569 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 13789 1569 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 13707 1569 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1529 13625 1569 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 4432 1555 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 4346 1555 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 4260 1555 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 4174 1555 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 4088 1555 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 4002 1555 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 3916 1555 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 3830 1555 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 3744 1555 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 3658 1555 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1515 3572 1555 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1459 18539 1499 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1459 18457 1499 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1459 18375 1499 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1459 18293 1499 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1459 18211 1499 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1459 18129 1499 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1459 18047 1499 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1459 17965 1499 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1459 17883 1499 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1459 17801 1499 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1459 17719 1499 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1459 17637 1499 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1459 17555 1499 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1459 17473 1499 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1459 17391 1499 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1459 17309 1499 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1459 17227 1499 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1459 17145 1499 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1459 17063 1499 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1459 16981 1499 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1459 16899 1499 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1459 16817 1499 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1459 16735 1499 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1459 16653 1499 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1459 16571 1499 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 16472 1489 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 16391 1489 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 16310 1489 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 16229 1489 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 16148 1489 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 16067 1489 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 15986 1489 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 15905 1489 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 15824 1489 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 15743 1489 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 15662 1489 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 15581 1489 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 15500 1489 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 15419 1489 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 15338 1489 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 15257 1489 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 15176 1489 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 15095 1489 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 15014 1489 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 14933 1489 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 14852 1489 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 14771 1489 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 14690 1489 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 14609 1489 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 14527 1489 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 14445 1489 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 14363 1489 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 14281 1489 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 14199 1489 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 14117 1489 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 14035 1489 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 13953 1489 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 13871 1489 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 13789 1489 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 13707 1489 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1449 13625 1489 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 4432 1474 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 4346 1474 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 4260 1474 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 4174 1474 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 4088 1474 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 4002 1474 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 3916 1474 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 3830 1474 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 3744 1474 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 3658 1474 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1434 3572 1474 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1377 18539 1417 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1377 18457 1417 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1377 18375 1417 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1377 18293 1417 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1377 18211 1417 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1377 18129 1417 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1377 18047 1417 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1377 17965 1417 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1377 17883 1417 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1377 17801 1417 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1377 17719 1417 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1377 17637 1417 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1377 17555 1417 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1377 17473 1417 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1377 17391 1417 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1377 17309 1417 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1377 17227 1417 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1377 17145 1417 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1377 17063 1417 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1377 16981 1417 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1377 16899 1417 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1377 16817 1417 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1377 16735 1417 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1377 16653 1417 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1377 16571 1417 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 16472 1409 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 16391 1409 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 16310 1409 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 16229 1409 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 16148 1409 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 16067 1409 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 15986 1409 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 15905 1409 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 15824 1409 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 15743 1409 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 15662 1409 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 15581 1409 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 15500 1409 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 15419 1409 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 15338 1409 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 15257 1409 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 15176 1409 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 15095 1409 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 15014 1409 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 14933 1409 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 14852 1409 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 14771 1409 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 14690 1409 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 14609 1409 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 14527 1409 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 14445 1409 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 14363 1409 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 14281 1409 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 14199 1409 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 14117 1409 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 14035 1409 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 13953 1409 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 13871 1409 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 13789 1409 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 13707 1409 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1369 13625 1409 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 4432 1393 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 4346 1393 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 4260 1393 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 4174 1393 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 4088 1393 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 4002 1393 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 3916 1393 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 3830 1393 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 3744 1393 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 3658 1393 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1353 3572 1393 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1295 18539 1335 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1295 18457 1335 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1295 18375 1335 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1295 18293 1335 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1295 18211 1335 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1295 18129 1335 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1295 18047 1335 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1295 17965 1335 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1295 17883 1335 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1295 17801 1335 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1295 17719 1335 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1295 17637 1335 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1295 17555 1335 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1295 17473 1335 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1295 17391 1335 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1295 17309 1335 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1295 17227 1335 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1295 17145 1335 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1295 17063 1335 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1295 16981 1335 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1295 16899 1335 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1295 16817 1335 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1295 16735 1335 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1295 16653 1335 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1295 16571 1335 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 16472 1329 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 16391 1329 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 16310 1329 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 16229 1329 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 16148 1329 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 16067 1329 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 15986 1329 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 15905 1329 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 15824 1329 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 15743 1329 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 15662 1329 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 15581 1329 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 15500 1329 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 15419 1329 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 15338 1329 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 15257 1329 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 15176 1329 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 15095 1329 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 15014 1329 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 14933 1329 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 14852 1329 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 14771 1329 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 14690 1329 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 14609 1329 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 14527 1329 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 14445 1329 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 14363 1329 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 14281 1329 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 14199 1329 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 14117 1329 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 14035 1329 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 13953 1329 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 13871 1329 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 13789 1329 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 13707 1329 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1289 13625 1329 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 4432 1312 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 4346 1312 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 4260 1312 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 4174 1312 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 4088 1312 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 4002 1312 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 3916 1312 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 3830 1312 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 3744 1312 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 3658 1312 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1272 3572 1312 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1213 18539 1253 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1213 18457 1253 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1213 18375 1253 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1213 18293 1253 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1213 18211 1253 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1213 18129 1253 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1213 18047 1253 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1213 17965 1253 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1213 17883 1253 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1213 17801 1253 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1213 17719 1253 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1213 17637 1253 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1213 17555 1253 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1213 17473 1253 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1213 17391 1253 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1213 17309 1253 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1213 17227 1253 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1213 17145 1253 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1213 17063 1253 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1213 16981 1253 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1213 16899 1253 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1213 16817 1253 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1213 16735 1253 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1213 16653 1253 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1213 16571 1253 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 16472 1249 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 16391 1249 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 16310 1249 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 16229 1249 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 16148 1249 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 16067 1249 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 15986 1249 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 15905 1249 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 15824 1249 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 15743 1249 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 15662 1249 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 15581 1249 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 15500 1249 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 15419 1249 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 15338 1249 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 15257 1249 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 15176 1249 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 15095 1249 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 15014 1249 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 14933 1249 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 14852 1249 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 14771 1249 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 14690 1249 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 14609 1249 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 14527 1249 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 14445 1249 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 14363 1249 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 14281 1249 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 14199 1249 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 14117 1249 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 14035 1249 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 13953 1249 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 13871 1249 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 13789 1249 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 13707 1249 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1209 13625 1249 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 4432 1231 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 4346 1231 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 4260 1231 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 4174 1231 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 4088 1231 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 4002 1231 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 3916 1231 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 3830 1231 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 3744 1231 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 3658 1231 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1191 3572 1231 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1131 18539 1171 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1131 18457 1171 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1131 18375 1171 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1131 18293 1171 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1131 18211 1171 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1131 18129 1171 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1131 18047 1171 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1131 17965 1171 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1131 17883 1171 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1131 17801 1171 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1131 17719 1171 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1131 17637 1171 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1131 17555 1171 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1131 17473 1171 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1131 17391 1171 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1131 17309 1171 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1131 17227 1171 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1131 17145 1171 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1131 17063 1171 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1131 16981 1171 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1131 16899 1171 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1131 16817 1171 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1131 16735 1171 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1131 16653 1171 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1131 16571 1171 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 16472 1169 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 16391 1169 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 16310 1169 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 16229 1169 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 16148 1169 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 16067 1169 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 15986 1169 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 15905 1169 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 15824 1169 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 15743 1169 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 15662 1169 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 15581 1169 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 15500 1169 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 15419 1169 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 15338 1169 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 15257 1169 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 15176 1169 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 15095 1169 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 15014 1169 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 14933 1169 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 14852 1169 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 14771 1169 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 14690 1169 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 14609 1169 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 14527 1169 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 14445 1169 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 14363 1169 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 14281 1169 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 14199 1169 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 14117 1169 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 14035 1169 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 13953 1169 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 13871 1169 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 13789 1169 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 13707 1169 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1129 13625 1169 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 4432 1150 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 4346 1150 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 4260 1150 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 4174 1150 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 4088 1150 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 4002 1150 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 3916 1150 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 3830 1150 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 3744 1150 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 3658 1150 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1110 3572 1150 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 18539 1089 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 18457 1089 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 18375 1089 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 18293 1089 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 18211 1089 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 18129 1089 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 18047 1089 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 17965 1089 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 17883 1089 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 17801 1089 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 17719 1089 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 17637 1089 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 17555 1089 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 17473 1089 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 17391 1089 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 17309 1089 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 17227 1089 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 17145 1089 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 17063 1089 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 16981 1089 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 16899 1089 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 16817 1089 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 16735 1089 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 16653 1089 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 16571 1089 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 16472 1089 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 16391 1089 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 16310 1089 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 16229 1089 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 16148 1089 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 16067 1089 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 15986 1089 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 15905 1089 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 15824 1089 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 15743 1089 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 15662 1089 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 15581 1089 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 15500 1089 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 15419 1089 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 15338 1089 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 15257 1089 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 15176 1089 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 15095 1089 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 15014 1089 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 14933 1089 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 14852 1089 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 14771 1089 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 14690 1089 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 14609 1089 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 14527 1089 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 14445 1089 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 14363 1089 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 14281 1089 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 14199 1089 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 14117 1089 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 14035 1089 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 13953 1089 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 13871 1089 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 13789 1089 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 13707 1089 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1049 13625 1089 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 4432 1069 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 4346 1069 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 4260 1069 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 4174 1069 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 4088 1069 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 4002 1069 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 3916 1069 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 3830 1069 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 3744 1069 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 3658 1069 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 1029 3572 1069 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 16472 1009 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 16391 1009 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 16310 1009 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 16229 1009 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 16148 1009 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 16067 1009 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 15986 1009 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 15905 1009 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 15824 1009 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 15743 1009 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 15662 1009 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 15581 1009 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 15500 1009 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 15419 1009 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 15338 1009 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 15257 1009 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 15176 1009 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 15095 1009 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 15014 1009 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 14933 1009 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 14852 1009 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 14771 1009 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 14690 1009 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 14609 1009 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 14527 1009 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 14445 1009 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 14363 1009 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 14281 1009 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 14199 1009 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 14117 1009 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 14035 1009 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 13953 1009 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 13871 1009 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 13789 1009 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 13707 1009 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 969 13625 1009 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 967 18539 1007 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 967 18457 1007 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 967 18375 1007 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 967 18293 1007 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 967 18211 1007 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 967 18129 1007 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 967 18047 1007 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 967 17965 1007 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 967 17883 1007 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 967 17801 1007 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 967 17719 1007 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 967 17637 1007 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 967 17555 1007 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 967 17473 1007 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 967 17391 1007 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 967 17309 1007 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 967 17227 1007 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 967 17145 1007 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 967 17063 1007 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 967 16981 1007 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 967 16899 1007 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 967 16817 1007 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 967 16735 1007 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 967 16653 1007 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 967 16571 1007 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 4432 988 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 4346 988 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 4260 988 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 4174 988 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 4088 988 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 4002 988 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 3916 988 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 3830 988 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 3744 988 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 3658 988 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 948 3572 988 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 16472 929 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 16391 929 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 16310 929 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 16229 929 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 16148 929 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 16067 929 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 15986 929 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 15905 929 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 15824 929 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 15743 929 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 15662 929 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 15581 929 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 15500 929 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 15419 929 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 15338 929 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 15257 929 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 15176 929 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 15095 929 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 15014 929 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 14933 929 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 14852 929 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 14771 929 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 14690 929 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 14609 929 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 14527 929 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 14445 929 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 14363 929 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 14281 929 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 14199 929 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 14117 929 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 14035 929 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 13953 929 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 13871 929 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 13789 929 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 13707 929 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 889 13625 929 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 885 18539 925 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 885 18457 925 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 885 18375 925 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 885 18293 925 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 885 18211 925 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 885 18129 925 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 885 18047 925 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 885 17965 925 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 885 17883 925 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 885 17801 925 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 885 17719 925 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 885 17637 925 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 885 17555 925 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 885 17473 925 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 885 17391 925 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 885 17309 925 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 885 17227 925 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 885 17145 925 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 885 17063 925 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 885 16981 925 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 885 16899 925 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 885 16817 925 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 885 16735 925 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 885 16653 925 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 885 16571 925 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 4432 907 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 4346 907 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 4260 907 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 4174 907 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 4088 907 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 4002 907 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 3916 907 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 3830 907 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 3744 907 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 3658 907 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 867 3572 907 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 16472 849 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 16391 849 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 16310 849 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 16229 849 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 16148 849 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 16067 849 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 15986 849 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 15905 849 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 15824 849 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 15743 849 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 15662 849 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 15581 849 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 15500 849 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 15419 849 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 15338 849 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 15257 849 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 15176 849 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 15095 849 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 15014 849 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 14933 849 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 14852 849 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 14771 849 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 14690 849 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 14609 849 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 14527 849 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 14445 849 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 14363 849 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 14281 849 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 14199 849 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 14117 849 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 14035 849 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 13953 849 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 13871 849 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 13789 849 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 13707 849 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 809 13625 849 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 803 18539 843 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 803 18457 843 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 803 18375 843 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 803 18293 843 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 803 18211 843 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 803 18129 843 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 803 18047 843 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 803 17965 843 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 803 17883 843 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 803 17801 843 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 803 17719 843 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 803 17637 843 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 803 17555 843 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 803 17473 843 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 803 17391 843 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 803 17309 843 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 803 17227 843 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 803 17145 843 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 803 17063 843 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 803 16981 843 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 803 16899 843 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 803 16817 843 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 803 16735 843 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 803 16653 843 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 803 16571 843 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 4432 826 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 4346 826 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 4260 826 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 4174 826 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 4088 826 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 4002 826 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 3916 826 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 3830 826 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 3744 826 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 3658 826 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 786 3572 826 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 16472 769 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 16391 769 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 16310 769 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 16229 769 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 16148 769 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 16067 769 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 15986 769 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 15905 769 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 15824 769 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 15743 769 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 15662 769 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 15581 769 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 15500 769 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 15419 769 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 15338 769 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 15257 769 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 15176 769 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 15095 769 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 15014 769 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 14933 769 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 14852 769 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 14771 769 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 14690 769 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 14609 769 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 14527 769 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 14445 769 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 14363 769 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 14281 769 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 14199 769 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 14117 769 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 14035 769 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 13953 769 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 13871 769 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 13789 769 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 13707 769 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 729 13625 769 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 721 18539 761 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 721 18457 761 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 721 18375 761 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 721 18293 761 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 721 18211 761 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 721 18129 761 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 721 18047 761 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 721 17965 761 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 721 17883 761 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 721 17801 761 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 721 17719 761 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 721 17637 761 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 721 17555 761 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 721 17473 761 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 721 17391 761 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 721 17309 761 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 721 17227 761 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 721 17145 761 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 721 17063 761 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 721 16981 761 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 721 16899 761 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 721 16817 761 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 721 16735 761 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 721 16653 761 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 721 16571 761 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 4432 745 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 4346 745 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 4260 745 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 4174 745 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 4088 745 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 4002 745 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 3916 745 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 3830 745 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 3744 745 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 3658 745 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 705 3572 745 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 16472 689 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 16391 689 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 16310 689 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 16229 689 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 16148 689 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 16067 689 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 15986 689 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 15905 689 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 15824 689 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 15743 689 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 15662 689 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 15581 689 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 15500 689 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 15419 689 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 15338 689 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 15257 689 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 15176 689 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 15095 689 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 15014 689 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 14933 689 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 14852 689 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 14771 689 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 14690 689 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 14609 689 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 14527 689 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 14445 689 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 14363 689 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 14281 689 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 14199 689 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 14117 689 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 14035 689 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 13953 689 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 13871 689 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 13789 689 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 13707 689 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 649 13625 689 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 639 18539 679 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 639 18457 679 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 639 18375 679 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 639 18293 679 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 639 18211 679 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 639 18129 679 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 639 18047 679 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 639 17965 679 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 639 17883 679 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 639 17801 679 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 639 17719 679 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 639 17637 679 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 639 17555 679 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 639 17473 679 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 639 17391 679 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 639 17309 679 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 639 17227 679 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 639 17145 679 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 639 17063 679 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 639 16981 679 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 639 16899 679 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 639 16817 679 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 639 16735 679 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 639 16653 679 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 639 16571 679 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 4432 664 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 4346 664 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 4260 664 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 4174 664 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 4088 664 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 4002 664 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 3916 664 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 3830 664 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 3744 664 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 3658 664 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 624 3572 664 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 16472 609 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 16391 609 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 16310 609 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 16229 609 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 16148 609 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 16067 609 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 15986 609 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 15905 609 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 15824 609 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 15743 609 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 15662 609 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 15581 609 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 15500 609 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 15419 609 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 15338 609 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 15257 609 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 15176 609 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 15095 609 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 15014 609 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 14933 609 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 14852 609 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 14771 609 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 14690 609 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 14609 609 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 14527 609 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 14445 609 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 14363 609 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 14281 609 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 14199 609 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 14117 609 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 14035 609 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 13953 609 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 13871 609 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 13789 609 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 13707 609 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 569 13625 609 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 18539 597 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 18457 597 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 18375 597 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 18293 597 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 18211 597 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 18129 597 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 18047 597 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 17965 597 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 17883 597 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 17801 597 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 17719 597 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 17637 597 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 17555 597 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 17473 597 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 17391 597 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 17309 597 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 17227 597 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 17145 597 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 17063 597 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 16981 597 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 16899 597 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 16817 597 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 16735 597 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 16653 597 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 557 16571 597 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 4432 583 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 4346 583 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 4260 583 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 4174 583 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 4088 583 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 4002 583 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 3916 583 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 3830 583 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 3744 583 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 3658 583 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 543 3572 583 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 16472 529 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 16391 529 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 16310 529 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 16229 529 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 16148 529 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 16067 529 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 15986 529 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 15905 529 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 15824 529 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 15743 529 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 15662 529 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 15581 529 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 15500 529 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 15419 529 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 15338 529 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 15257 529 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 15176 529 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 15095 529 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 15014 529 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 14933 529 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 14852 529 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 14771 529 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 14690 529 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 14609 529 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 14527 529 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 14445 529 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 14363 529 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 14281 529 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 14199 529 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 14117 529 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 14035 529 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 13953 529 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 13871 529 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 13789 529 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 13707 529 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 489 13625 529 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 475 18539 515 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 475 18457 515 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 475 18375 515 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 475 18293 515 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 475 18211 515 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 475 18129 515 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 475 18047 515 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 475 17965 515 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 475 17883 515 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 475 17801 515 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 475 17719 515 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 475 17637 515 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 475 17555 515 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 475 17473 515 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 475 17391 515 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 475 17309 515 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 475 17227 515 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 475 17145 515 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 475 17063 515 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 475 16981 515 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 475 16899 515 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 475 16817 515 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 475 16735 515 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 475 16653 515 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 475 16571 515 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 4432 502 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 4346 502 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 4260 502 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 4174 502 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 4088 502 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 4002 502 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 3916 502 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 3830 502 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 3744 502 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 3658 502 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 462 3572 502 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 16472 449 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 16391 449 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 16310 449 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 16229 449 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 16148 449 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 16067 449 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 15986 449 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 15905 449 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 15824 449 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 15743 449 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 15662 449 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 15581 449 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 15500 449 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 15419 449 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 15338 449 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 15257 449 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 15176 449 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 15095 449 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 15014 449 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 14933 449 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 14852 449 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 14771 449 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 14690 449 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 14609 449 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 14527 449 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 14445 449 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 14363 449 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 14281 449 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 14199 449 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 14117 449 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 14035 449 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 13953 449 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 13871 449 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 13789 449 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 13707 449 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 409 13625 449 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 393 18539 433 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 393 18457 433 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 393 18375 433 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 393 18293 433 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 393 18211 433 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 393 18129 433 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 393 18047 433 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 393 17965 433 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 393 17883 433 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 393 17801 433 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 393 17719 433 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 393 17637 433 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 393 17555 433 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 393 17473 433 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 393 17391 433 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 393 17309 433 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 393 17227 433 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 393 17145 433 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 393 17063 433 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 393 16981 433 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 393 16899 433 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 393 16817 433 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 393 16735 433 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 393 16653 433 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 393 16571 433 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 4432 421 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 4346 421 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 4260 421 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 4174 421 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 4088 421 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 4002 421 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 3916 421 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 3830 421 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 3744 421 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 3658 421 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 381 3572 421 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 16472 369 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 16391 369 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 16310 369 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 16229 369 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 16148 369 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 16067 369 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 15986 369 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 15905 369 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 15824 369 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 15743 369 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 15662 369 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 15581 369 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 15500 369 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 15419 369 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 15338 369 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 15257 369 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 15176 369 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 15095 369 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 15014 369 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 14933 369 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 14852 369 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 14771 369 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 14690 369 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 14609 369 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 14527 369 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 14445 369 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 14363 369 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 14281 369 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 14199 369 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 14117 369 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 14035 369 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 13953 369 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 13871 369 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 13789 369 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 13707 369 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 329 13625 369 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 311 18539 351 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 311 18457 351 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 311 18375 351 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 311 18293 351 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 311 18211 351 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 311 18129 351 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 311 18047 351 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 311 17965 351 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 311 17883 351 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 311 17801 351 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 311 17719 351 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 311 17637 351 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 311 17555 351 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 311 17473 351 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 311 17391 351 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 311 17309 351 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 311 17227 351 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 311 17145 351 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 311 17063 351 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 311 16981 351 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 311 16899 351 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 311 16817 351 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 311 16735 351 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 311 16653 351 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 311 16571 351 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 4432 340 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 4346 340 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 4260 340 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 4174 340 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 4088 340 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 4002 340 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 3916 340 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 3830 340 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 3744 340 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 3658 340 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 300 3572 340 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 16472 289 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 16391 289 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 16310 289 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 16229 289 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 16148 289 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 16067 289 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 15986 289 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 15905 289 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 15824 289 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 15743 289 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 15662 289 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 15581 289 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 15500 289 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 15419 289 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 15338 289 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 15257 289 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 15176 289 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 15095 289 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 15014 289 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 14933 289 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 14852 289 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 14771 289 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 14690 289 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 14609 289 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 14527 289 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 14445 289 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 14363 289 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 14281 289 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 14199 289 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 14117 289 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 14035 289 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 13953 289 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 13871 289 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 13789 289 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 13707 289 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 249 13625 289 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 229 18539 269 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 229 18457 269 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 229 18375 269 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 229 18293 269 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 229 18211 269 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 229 18129 269 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 229 18047 269 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 229 17965 269 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 229 17883 269 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 229 17801 269 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 229 17719 269 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 229 17637 269 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 229 17555 269 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 229 17473 269 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 229 17391 269 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 229 17309 269 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 229 17227 269 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 229 17145 269 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 229 17063 269 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 229 16981 269 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 229 16899 269 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 229 16817 269 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 229 16735 269 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 229 16653 269 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 229 16571 269 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 4432 259 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 4346 259 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 4260 259 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 4174 259 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 4088 259 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 4002 259 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 3916 259 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 3830 259 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 3744 259 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 3658 259 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 219 3572 259 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 16472 209 16512 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 16391 209 16431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 16310 209 16350 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 16229 209 16269 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 16148 209 16188 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 16067 209 16107 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 15986 209 16026 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 15905 209 15945 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 15824 209 15864 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 15743 209 15783 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 15662 209 15702 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 15581 209 15621 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 15500 209 15540 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 15419 209 15459 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 15338 209 15378 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 15257 209 15297 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 15176 209 15216 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 15095 209 15135 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 15014 209 15054 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 14933 209 14973 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 14852 209 14892 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 14771 209 14811 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 14690 209 14730 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 14609 209 14649 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 14527 209 14567 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 14445 209 14485 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 14363 209 14403 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 14281 209 14321 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 14199 209 14239 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 14117 209 14157 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 14035 209 14075 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 13953 209 13993 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 13871 209 13911 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 13789 209 13829 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 13707 209 13747 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 169 13625 209 13665 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 147 18539 187 18579 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 147 18457 187 18497 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 147 18375 187 18415 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 147 18293 187 18333 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 147 18211 187 18251 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 147 18129 187 18169 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 147 18047 187 18087 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 147 17965 187 18005 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 147 17883 187 17923 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 147 17801 187 17841 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 147 17719 187 17759 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 147 17637 187 17677 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 147 17555 187 17595 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 147 17473 187 17513 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 147 17391 187 17431 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 147 17309 187 17349 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 147 17227 187 17267 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 147 17145 187 17185 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 147 17063 187 17103 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 147 16981 187 17021 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 147 16899 187 16939 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 147 16817 187 16857 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 147 16735 187 16775 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 147 16653 187 16693 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 147 16571 187 16611 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 4432 178 4472 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 4346 178 4386 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 4260 178 4300 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 4174 178 4214 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 4088 178 4128 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 4002 178 4042 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 3916 178 3956 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 3830 178 3870 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 3744 178 3784 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 3658 178 3698 6 VDDIO
port 7 nsew power bidirectional
rlabel metal3 s 138 3572 178 3612 6 VDDIO
port 7 nsew power bidirectional
rlabel metal5 s 0 5997 254 6647 6 VSWITCH
port 8 nsew power bidirectional
rlabel metal5 s 14746 5997 15000 6647 6 VSWITCH
port 8 nsew power bidirectional
rlabel metal4 s 0 5977 254 6667 6 VSWITCH
port 8 nsew power bidirectional
rlabel metal4 s 14746 5977 15000 6667 6 VSWITCH
port 8 nsew power bidirectional
rlabel metal4 s 14746 5977 15000 6667 6 VSWITCH
port 8 nsew power bidirectional
rlabel metal5 s 0 5997 254 6647 6 VSWITCH
port 8 nsew power bidirectional
rlabel metal5 s 14746 5997 15000 6647 6 VSWITCH
port 8 nsew power bidirectional
rlabel metal4 s 14746 5977 15000 6667 6 VSWITCH
port 8 nsew power bidirectional
rlabel metal5 s 0 5997 254 6647 6 VSWITCH
port 8 nsew power bidirectional
rlabel metal5 s 14746 5997 15000 6647 6 VSWITCH
port 8 nsew power bidirectional
rlabel metal5 s 0 11267 254 12117 6 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal5 s 14746 11267 15000 12117 6 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal4 s 0 11247 254 12137 6 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal4 s 14746 11247 15000 12137 6 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal4 s 14746 11247 15000 12137 6 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal5 s 0 11267 254 12117 6 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal5 s 14746 11267 15000 12117 6 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal4 s 14746 11247 15000 12137 6 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal5 s 0 11267 254 12117 6 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal5 s 14746 11267 15000 12117 6 VSSIO_Q
port 9 nsew ground bidirectional
rlabel metal5 s 0 4787 254 5677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal5 s 0 34757 254 39600 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal5 s 14746 4787 15000 5677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal5 s 14746 34757 15000 39600 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 0 4767 254 5697 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 0 34757 254 39600 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14746 4767 15000 5697 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14746 34757 15000 39600 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 0 4767 254 5697 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14746 34757 15000 39600 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14746 4767 15000 5697 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal5 s 0 34757 254 39600 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal5 s 0 4787 254 5677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal5 s 14746 34757 15000 39600 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal5 s 14746 4787 15000 5677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 0 4767 254 5697 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14746 34757 15000 39600 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 14746 4767 15000 5697 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal5 s 0 34757 254 39600 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal5 s 0 4787 254 5677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal5 s 14746 34757 15000 39600 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal5 s 14746 4787 15000 5677 6 VSSIO
port 10 nsew ground bidirectional
rlabel metal4 s 0 10225 15000 10821 6 AMUXBUS_A
port 11 nsew signal bidirectional
rlabel metal4 s 0 10225 254 10821 6 AMUXBUS_A
port 11 nsew signal bidirectional
rlabel metal4 s 14746 10225 15000 10821 6 AMUXBUS_A
port 11 nsew signal bidirectional
rlabel metal4 s 14746 10225 15000 10821 6 AMUXBUS_A
port 11 nsew signal bidirectional
rlabel metal4 s 0 9273 15000 9869 6 AMUXBUS_B
port 12 nsew signal bidirectional
rlabel metal4 s 0 9273 254 9869 6 AMUXBUS_B
port 12 nsew signal bidirectional
rlabel metal4 s 14746 9273 15000 9869 6 AMUXBUS_B
port 12 nsew signal bidirectional
rlabel metal4 s 14746 9273 15000 9869 6 AMUXBUS_B
port 12 nsew signal bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 15000 39600
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 17269118
string GDS_START 16685534
<< end >>
