* NGSPICE file created from Bandgap1v8.ext - technology: sky130A


* Top level circuit Bandgap1v8

X0 G1011 G1011 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u M=44
X1 G1011 D6 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u M=10
X2 D5 G1011 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u M=4
X3 GND GND VBJTS sky130_fd_pr__pnp_05v0 area=0p M=-nan
X4 D9 G4 D5 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=500000u M=6
X5 G3 Vref GND sky130_fd_pr__res_xhigh_po w=1.41e+06u l=1.8e+06u
X6 VDD G1011 Vref VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u M=4
X7 GND GND G4 sky130_fd_pr__pnp_05v0 area=0p
X8 GND D9 D9 GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u M=4
X9 D5 G3 D6 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+07u l=500000u M=6
X10 D6 D9 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=500000u M=4
X11 a_523_n9665# a_n7_n8873# GND sky130_fd_pr__res_xhigh_po w=1.41e+06u l=1.8e+06u
X12 a_2643_n9665# a_3173_n8873# GND sky130_fd_pr__res_xhigh_po w=1.41e+06u l=1.8e+06u
X13 D1011 G1011 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=1e+06u M=2
X14 G4 D1011 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+07u l=1e+06u M=2
X15 VDD G1011 D2 VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u M=4
X16 G3 a_n7_n8873# GND sky130_fd_pr__res_xhigh_po w=1.41e+06u l=1.8e+06u
X17 G4 a_3173_n8873# GND sky130_fd_pr__res_xhigh_po w=1.41e+06u l=1.8e+06u
X18 D1011 G1011 GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=2e+07u
X19 a_2643_n9665# a_2113_n8873# GND sky130_fd_pr__res_xhigh_po w=1.41e+06u l=1.8e+06u
X20 VBJTS a_1053_n8873# GND sky130_fd_pr__res_xhigh_po w=1.41e+06u l=1.8e+06u
X21 D2 a_2113_n8873# GND sky130_fd_pr__res_xhigh_po w=1.41e+06u l=1.8e+06u
X22 a_523_n9665# a_1053_n8873# GND sky130_fd_pr__res_xhigh_po w=1.41e+06u l=1.8e+06u
.end

