magic
tech sky130A
magscale 1 2
timestamp 1624884114
<< metal3 >>
rect 10078 11648 14858 12536
rect 99 5168 4879 6096
rect 10078 5168 14858 6096
<< obsm3 >>
rect 99 12616 14858 40000
rect 99 11648 9998 12616
<< metal4 >>
rect 0 39984 254 40000
rect 0 35186 2695 39984
rect 2726 39434 12265 39986
rect 14746 39984 15000 40000
rect 2719 39246 2851 39394
rect 12136 39246 12268 39394
rect 0 35157 254 35186
rect 12301 35186 15000 39984
rect 14746 35157 15000 35186
rect 0 14007 254 19000
rect 14746 14007 15000 19000
rect 0 12817 254 13707
rect 14746 12817 15000 13707
rect 0 11647 4874 12537
rect 10083 11647 15000 12537
rect 0 11281 15000 11347
rect 0 10625 15000 11221
rect 0 10329 254 10565
rect 14746 10329 15000 10565
rect 0 9673 15000 10269
rect 0 9547 15000 9613
rect 0 8317 254 9247
rect 14746 8317 15000 9247
rect 0 7347 254 8037
rect 14746 7347 15000 8037
rect 0 6377 254 7067
rect 14746 6377 15000 7067
rect 0 5167 4874 6097
rect 10083 5167 15000 6097
rect 0 3957 254 4887
rect 14746 3957 15000 4887
rect 0 2987 193 3677
rect 14807 2987 15000 3677
rect 0 1777 254 2707
rect 14746 1777 15000 2707
rect 0 407 254 1497
rect 14746 407 15000 1497
<< obsm4 >>
rect 2931 39166 12056 39354
rect 2775 35106 12221 39166
rect 334 35077 14666 35106
rect 193 19080 14807 35077
rect 334 13927 14666 19080
rect 193 13787 14807 13927
rect 334 12737 14666 13787
rect 193 12617 14807 12737
rect 4954 11567 10003 12617
rect 193 11427 14807 11567
rect 334 10349 14666 10545
rect 193 9327 14807 9467
rect 334 8237 14666 9327
rect 193 8117 14807 8237
rect 334 7267 14666 8117
rect 193 7147 14807 7267
rect 334 6297 14666 7147
rect 193 6177 14807 6297
rect 4954 5087 10003 6177
rect 193 4967 14807 5087
rect 334 3877 14666 4967
rect 193 3757 14807 3877
rect 273 2907 14727 3757
rect 193 2787 14807 2907
rect 334 1697 14666 2787
rect 193 1577 14807 1697
rect 334 407 14666 1577
<< metal5 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 0 14007 254 18997
rect 0 12837 254 13687
rect 0 11667 254 12517
rect 0 9547 254 11347
rect 0 8337 254 9227
rect 0 7368 254 8017
rect 14746 14007 15000 18997
rect 14746 12837 15000 13687
rect 14746 11667 15000 12517
rect 14746 9547 15000 11347
rect 14746 8337 15000 9227
rect 14746 7368 15000 8017
rect 0 6397 254 7047
rect 0 5187 254 6077
rect 0 3977 254 4867
rect 14746 6397 15000 7047
rect 14746 5187 15000 6077
rect 14746 3977 15000 4867
rect 0 3007 193 3657
rect 14807 3007 15000 3657
rect 0 1797 254 2687
rect 0 427 254 1477
rect 14746 1797 15000 2687
rect 14746 427 15000 1477
<< obsm5 >>
rect 574 34837 14426 40000
rect 0 19317 15000 34837
rect 574 7368 14426 19317
rect 0 7367 15000 7368
rect 574 3657 14426 7367
rect 513 3007 14487 3657
rect 574 427 14426 3007
<< labels >>
rlabel metal5 s 0 9547 254 11347 6 VSSA
port 1 nsew ground bidirectional
rlabel metal5 s 0 7368 254 8017 6 VSSA
port 1 nsew ground bidirectional
rlabel metal5 s 14746 9547 15000 11347 6 VSSA
port 1 nsew ground bidirectional
rlabel metal5 s 14746 7368 15000 8017 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 0 11281 15000 11347 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 0 9547 15000 9613 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 0 10329 254 10565 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 0 7347 254 8037 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 14746 11281 15000 11347 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 14746 9547 15000 9613 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 14746 10329 15000 10565 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 14746 7347 15000 8037 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 0 9547 254 9613 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 0 10329 254 10565 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 0 11281 254 11347 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 14746 7347 15000 8037 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 14746 9547 15000 9613 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 14746 10329 15000 10565 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 14746 11281 15000 11347 6 VSSA
port 1 nsew ground bidirectional
rlabel metal5 s 0 7368 254 8017 6 VSSA
port 1 nsew ground bidirectional
rlabel metal5 s 0 9547 254 11347 6 VSSA
port 1 nsew ground bidirectional
rlabel metal5 s 14746 7368 15000 8017 6 VSSA
port 1 nsew ground bidirectional
rlabel metal5 s 14746 9547 15000 11347 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 0 9547 254 9613 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 0 10329 254 10565 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 0 11281 254 11347 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 14746 7347 15000 8037 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 14746 9547 15000 9613 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 14746 10329 15000 10565 6 VSSA
port 1 nsew ground bidirectional
rlabel metal4 s 14746 11281 15000 11347 6 VSSA
port 1 nsew ground bidirectional
rlabel metal5 s 0 7368 254 8017 6 VSSA
port 1 nsew ground bidirectional
rlabel metal5 s 0 9547 254 11347 6 VSSA
port 1 nsew ground bidirectional
rlabel metal5 s 14746 7368 15000 8017 6 VSSA
port 1 nsew ground bidirectional
rlabel metal5 s 14746 9547 15000 11347 6 VSSA
port 1 nsew ground bidirectional
rlabel metal5 s 0 14007 254 18997 6 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 0 3977 254 4867 6 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 14746 14007 15000 18997 6 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 14746 3977 15000 4867 6 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 0 3957 254 4887 6 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 0 14007 254 19000 6 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 14746 3957 15000 4887 6 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 14746 14007 15000 19000 6 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 0 14007 254 19000 6 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 14746 3957 15000 4887 6 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 14746 14007 15000 19000 6 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 0 3977 254 4867 6 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 0 14007 254 18997 6 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 14746 3977 15000 4867 6 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 14746 14007 15000 18997 6 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 0 14007 254 19000 6 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 14746 3957 15000 4887 6 VDDIO
port 2 nsew power bidirectional
rlabel metal4 s 14746 14007 15000 19000 6 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 0 3977 254 4867 6 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 0 14007 254 18997 6 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 14746 3977 15000 4867 6 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 14746 14007 15000 18997 6 VDDIO
port 2 nsew power bidirectional
rlabel metal5 s 0 12837 254 13687 6 VDDIO_Q
port 3 nsew power bidirectional
rlabel metal5 s 14746 12837 15000 13687 6 VDDIO_Q
port 3 nsew power bidirectional
rlabel metal4 s 0 12817 254 13707 6 VDDIO_Q
port 3 nsew power bidirectional
rlabel metal4 s 14746 12817 15000 13707 6 VDDIO_Q
port 3 nsew power bidirectional
rlabel metal4 s 14746 12817 15000 13707 6 VDDIO_Q
port 3 nsew power bidirectional
rlabel metal5 s 0 12837 254 13687 6 VDDIO_Q
port 3 nsew power bidirectional
rlabel metal5 s 14746 12837 15000 13687 6 VDDIO_Q
port 3 nsew power bidirectional
rlabel metal4 s 14746 12817 15000 13707 6 VDDIO_Q
port 3 nsew power bidirectional
rlabel metal5 s 0 12837 254 13687 6 VDDIO_Q
port 3 nsew power bidirectional
rlabel metal5 s 14746 12837 15000 13687 6 VDDIO_Q
port 3 nsew power bidirectional
rlabel metal5 s 0 8337 254 9227 6 VSSD
port 4 nsew ground bidirectional
rlabel metal5 s 14746 8337 15000 9227 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 0 8317 254 9247 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 14746 8317 15000 9247 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 14746 8317 15000 9247 6 VSSD
port 4 nsew ground bidirectional
rlabel metal5 s 0 8337 254 9227 6 VSSD
port 4 nsew ground bidirectional
rlabel metal5 s 14746 8337 15000 9227 6 VSSD
port 4 nsew ground bidirectional
rlabel metal4 s 14746 8317 15000 9247 6 VSSD
port 4 nsew ground bidirectional
rlabel metal5 s 0 8337 254 9227 6 VSSD
port 4 nsew ground bidirectional
rlabel metal5 s 14746 8337 15000 9227 6 VSSD
port 4 nsew ground bidirectional
rlabel metal5 s 0 5187 254 6077 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 14746 5187 15000 6077 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 14746 35157 15000 40000 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 0 35157 254 40000 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 0 5167 254 6097 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14746 5167 15000 6097 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14746 35157 15000 40000 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 0 35157 254 40000 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 126 38320 128 38322 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 99 5168 4879 6096 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10078 5168 14858 6096 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 0 39984 254 40000 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 0 35186 2695 39984 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 0 35157 254 35186 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 0 5167 4874 6097 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2719 39246 2851 39394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2726 39434 12265 39986 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 10083 5167 15000 6097 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12136 39246 12268 39394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14746 39984 15000 40000 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14746 35157 15000 35186 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12301 35186 15000 39984 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 0 35157 254 40000 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 0 5187 254 6077 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 14746 35157 15000 40000 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 14746 5187 15000 6077 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 6042 14840 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5956 14840 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5870 14840 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5784 14840 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5698 14840 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5612 14840 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5526 14840 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5440 14840 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5354 14840 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5268 14840 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5182 14840 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14786 39919 14850 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14786 39838 14850 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14786 39757 14850 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14786 39676 14850 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14786 39595 14850 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14786 39514 14850 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14786 39433 14850 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14786 39352 14850 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14786 39271 14850 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14786 39190 14850 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14786 39109 14850 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14786 39028 14850 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12306 35187 14850 39011 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 38879 14838 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 38799 14838 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 38719 14838 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 38639 14838 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 38559 14838 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 38479 14838 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 38399 14838 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 38319 14838 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 38239 14838 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 38159 14838 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 38079 14838 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 37999 14838 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 37919 14838 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 37839 14838 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 37759 14838 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 37679 14838 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 37599 14838 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 37519 14838 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 37439 14838 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 37359 14838 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 37279 14838 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 37199 14838 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 37119 14838 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 37039 14838 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 36959 14838 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 36879 14838 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 36799 14838 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 36719 14838 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 36639 14838 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 36559 14838 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 36479 14838 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 36399 14838 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 36319 14838 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 36239 14838 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 36159 14838 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 36079 14838 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 35999 14838 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 35919 14838 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 35839 14838 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 35759 14838 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 35679 14838 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 35599 14838 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 35519 14838 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 35439 14838 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 35359 14838 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 35279 14838 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 35199 14838 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 6042 14759 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5956 14759 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5870 14759 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5784 14759 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5698 14759 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5612 14759 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5526 14759 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5440 14759 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5354 14759 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5268 14759 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5182 14759 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14706 39919 14770 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14706 39838 14770 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14706 39757 14770 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14706 39676 14770 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14706 39595 14770 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14706 39514 14770 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14706 39433 14770 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14706 39352 14770 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14706 39271 14770 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14706 39190 14770 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14706 39109 14770 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14706 39028 14770 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 38959 14758 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 38879 14758 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 38799 14758 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 38719 14758 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 38639 14758 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 38559 14758 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 38479 14758 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 38399 14758 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 38319 14758 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 38239 14758 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 38159 14758 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 38079 14758 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 37999 14758 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 37919 14758 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 37839 14758 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 37759 14758 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 37679 14758 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 37599 14758 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 37519 14758 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 37439 14758 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 37359 14758 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 37279 14758 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 37199 14758 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 37119 14758 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 37039 14758 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 36959 14758 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 36879 14758 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 36799 14758 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 36719 14758 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 36639 14758 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 36559 14758 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 36479 14758 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 36399 14758 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 36319 14758 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 36239 14758 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 36159 14758 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 36079 14758 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 35999 14758 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 35919 14758 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 35839 14758 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 35759 14758 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 35679 14758 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 35599 14758 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 35519 14758 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 35439 14758 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 35359 14758 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 35279 14758 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 35199 14758 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14626 39919 14690 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14626 39838 14690 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14626 39757 14690 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14626 39676 14690 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14626 39595 14690 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14626 39514 14690 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14626 39433 14690 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14626 39352 14690 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14626 39271 14690 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14626 39190 14690 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14626 39109 14690 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14626 39028 14690 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 38959 14678 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 38879 14678 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 38799 14678 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 38719 14678 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 38639 14678 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 38559 14678 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 38479 14678 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 38399 14678 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 38319 14678 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 38239 14678 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 38159 14678 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 38079 14678 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 37999 14678 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 37919 14678 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 37839 14678 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 37759 14678 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 37679 14678 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 37599 14678 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 37519 14678 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 37439 14678 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 37359 14678 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 37279 14678 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 37199 14678 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 37119 14678 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 37039 14678 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 36959 14678 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 36879 14678 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 36799 14678 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 36719 14678 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 36639 14678 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 36559 14678 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 36479 14678 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 36399 14678 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 36319 14678 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 36239 14678 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 36159 14678 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 36079 14678 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 35999 14678 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 35919 14678 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 35839 14678 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 35759 14678 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 35679 14678 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 35599 14678 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 35519 14678 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 35439 14678 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 35359 14678 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 35279 14678 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 35199 14678 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 6042 14678 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 5956 14678 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 5870 14678 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 5784 14678 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 5698 14678 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 5612 14678 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 5526 14678 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 5440 14678 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 5354 14678 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 5268 14678 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 5182 14678 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14546 39919 14610 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14546 39838 14610 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14546 39757 14610 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14546 39676 14610 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14546 39595 14610 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14546 39514 14610 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14546 39433 14610 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14546 39352 14610 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14546 39271 14610 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14546 39190 14610 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14546 39109 14610 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14546 39028 14610 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 38959 14598 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 38879 14598 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 38799 14598 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 38719 14598 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 38639 14598 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 38559 14598 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 38479 14598 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 38399 14598 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 38319 14598 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 38239 14598 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 38159 14598 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 38079 14598 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 37999 14598 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 37919 14598 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 37839 14598 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 37759 14598 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 37679 14598 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 37599 14598 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 37519 14598 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 37439 14598 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 37359 14598 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 37279 14598 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 37199 14598 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 37119 14598 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 37039 14598 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 36959 14598 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 36879 14598 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 36799 14598 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 36719 14598 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 36639 14598 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 36559 14598 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 36479 14598 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 36399 14598 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 36319 14598 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 36239 14598 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 36159 14598 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 36079 14598 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 35999 14598 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 35919 14598 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 35839 14598 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 35759 14598 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 35679 14598 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 35599 14598 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 35519 14598 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 35439 14598 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 35359 14598 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 35279 14598 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 35199 14598 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 6042 14597 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5956 14597 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5870 14597 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5784 14597 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5698 14597 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5612 14597 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5526 14597 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5440 14597 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5354 14597 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5268 14597 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5182 14597 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14466 39919 14530 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14466 39838 14530 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14466 39757 14530 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14466 39676 14530 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14466 39595 14530 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14466 39514 14530 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14466 39433 14530 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14466 39352 14530 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14466 39271 14530 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14466 39190 14530 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14466 39109 14530 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14466 39028 14530 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 38959 14518 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 38879 14518 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 38799 14518 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 38719 14518 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 38639 14518 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 38559 14518 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 38479 14518 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 38399 14518 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 38319 14518 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 38239 14518 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 38159 14518 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 38079 14518 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 37999 14518 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 37919 14518 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 37839 14518 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 37759 14518 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 37679 14518 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 37599 14518 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 37519 14518 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 37439 14518 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 37359 14518 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 37279 14518 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 37199 14518 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 37119 14518 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 37039 14518 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 36959 14518 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 36879 14518 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 36799 14518 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 36719 14518 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 36639 14518 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 36559 14518 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 36479 14518 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 36399 14518 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 36319 14518 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 36239 14518 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 36159 14518 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 36079 14518 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 35999 14518 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 35919 14518 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 35839 14518 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 35759 14518 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 35679 14518 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 35599 14518 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 35519 14518 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 35439 14518 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 35359 14518 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 35279 14518 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 35199 14518 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14476 6042 14516 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14476 5956 14516 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14476 5870 14516 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14476 5784 14516 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14476 5698 14516 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14476 5612 14516 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14476 5526 14516 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14476 5440 14516 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14476 5354 14516 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14476 5268 14516 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14476 5182 14516 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14386 39919 14450 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14386 39838 14450 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14386 39757 14450 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14386 39676 14450 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14386 39595 14450 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14386 39514 14450 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14386 39433 14450 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14386 39352 14450 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14386 39271 14450 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14386 39190 14450 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14386 39109 14450 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14386 39028 14450 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 38959 14438 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 38879 14438 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 38799 14438 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 38719 14438 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 38639 14438 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 38559 14438 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 38479 14438 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 38399 14438 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 38319 14438 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 38239 14438 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 38159 14438 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 38079 14438 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 37999 14438 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 37919 14438 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 37839 14438 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 37759 14438 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 37679 14438 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 37599 14438 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 37519 14438 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 37439 14438 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 37359 14438 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 37279 14438 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 37199 14438 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 37119 14438 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 37039 14438 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 36959 14438 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 36879 14438 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 36799 14438 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 36719 14438 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 36639 14438 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 36559 14438 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 36479 14438 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 36399 14438 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 36319 14438 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 36239 14438 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 36159 14438 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 36079 14438 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 35999 14438 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 35919 14438 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 35839 14438 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 35759 14438 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 35679 14438 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 35599 14438 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 35519 14438 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 35439 14438 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 35359 14438 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 35279 14438 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 35199 14438 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14395 6042 14435 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14395 5956 14435 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14395 5870 14435 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14395 5784 14435 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14395 5698 14435 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14395 5612 14435 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14395 5526 14435 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14395 5440 14435 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14395 5354 14435 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14395 5268 14435 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14395 5182 14435 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14306 39919 14370 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14306 39838 14370 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14306 39757 14370 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14306 39676 14370 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14306 39595 14370 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14306 39514 14370 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14306 39433 14370 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14306 39352 14370 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14306 39271 14370 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14306 39190 14370 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14306 39109 14370 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14306 39028 14370 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 38959 14358 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 38879 14358 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 38799 14358 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 38719 14358 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 38639 14358 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 38559 14358 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 38479 14358 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 38399 14358 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 38319 14358 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 38239 14358 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 38159 14358 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 38079 14358 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 37999 14358 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 37919 14358 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 37839 14358 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 37759 14358 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 37679 14358 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 37599 14358 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 37519 14358 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 37439 14358 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 37359 14358 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 37279 14358 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 37199 14358 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 37119 14358 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 37039 14358 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 36959 14358 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 36879 14358 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 36799 14358 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 36719 14358 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 36639 14358 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 36559 14358 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 36479 14358 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 36399 14358 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 36319 14358 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 36239 14358 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 36159 14358 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 36079 14358 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 35999 14358 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 35919 14358 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 35839 14358 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 35759 14358 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 35679 14358 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 35599 14358 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 35519 14358 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 35439 14358 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 35359 14358 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 35279 14358 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 35199 14358 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14314 6042 14354 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14314 5956 14354 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14314 5870 14354 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14314 5784 14354 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14314 5698 14354 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14314 5612 14354 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14314 5526 14354 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14314 5440 14354 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14314 5354 14354 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14314 5268 14354 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14314 5182 14354 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14226 39919 14290 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14226 39838 14290 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14226 39757 14290 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14226 39676 14290 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14226 39595 14290 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14226 39514 14290 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14226 39433 14290 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14226 39352 14290 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14226 39271 14290 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14226 39190 14290 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14226 39109 14290 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14226 39028 14290 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 38959 14278 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 38879 14278 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 38799 14278 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 38719 14278 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 38639 14278 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 38559 14278 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 38479 14278 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 38399 14278 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 38319 14278 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 38239 14278 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 38159 14278 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 38079 14278 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 37999 14278 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 37919 14278 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 37839 14278 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 37759 14278 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 37679 14278 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 37599 14278 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 37519 14278 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 37439 14278 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 37359 14278 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 37279 14278 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 37199 14278 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 37119 14278 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 37039 14278 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 36959 14278 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 36879 14278 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 36799 14278 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 36719 14278 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 36639 14278 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 36559 14278 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 36479 14278 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 36399 14278 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 36319 14278 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 36239 14278 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 36159 14278 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 36079 14278 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 35999 14278 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 35919 14278 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 35839 14278 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 35759 14278 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 35679 14278 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 35599 14278 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 35519 14278 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 35439 14278 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 35359 14278 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 35279 14278 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 35199 14278 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 6042 14273 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5956 14273 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5870 14273 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5784 14273 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5698 14273 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5612 14273 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5526 14273 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5440 14273 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5354 14273 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5268 14273 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5182 14273 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14146 39919 14210 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14146 39838 14210 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14146 39757 14210 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14146 39676 14210 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14146 39595 14210 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14146 39514 14210 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14146 39433 14210 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14146 39352 14210 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14146 39271 14210 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14146 39190 14210 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14146 39109 14210 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14146 39028 14210 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 38959 14198 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 38879 14198 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 38799 14198 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 38719 14198 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 38639 14198 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 38559 14198 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 38479 14198 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 38399 14198 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 38319 14198 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 38239 14198 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 38159 14198 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 38079 14198 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 37999 14198 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 37919 14198 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 37839 14198 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 37759 14198 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 37679 14198 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 37599 14198 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 37519 14198 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 37439 14198 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 37359 14198 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 37279 14198 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 37199 14198 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 37119 14198 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 37039 14198 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 36959 14198 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 36879 14198 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 36799 14198 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 36719 14198 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 36639 14198 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 36559 14198 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 36479 14198 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 36399 14198 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 36319 14198 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 36239 14198 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 36159 14198 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 36079 14198 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 35999 14198 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 35919 14198 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 35839 14198 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 35759 14198 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 35679 14198 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 35599 14198 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 35519 14198 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 35439 14198 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 35359 14198 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 35279 14198 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 35199 14198 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14152 6042 14192 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14152 5956 14192 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14152 5870 14192 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14152 5784 14192 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14152 5698 14192 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14152 5612 14192 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14152 5526 14192 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14152 5440 14192 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14152 5354 14192 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14152 5268 14192 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14152 5182 14192 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14066 39919 14130 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14066 39838 14130 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14066 39757 14130 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14066 39676 14130 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14066 39595 14130 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14066 39514 14130 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14066 39433 14130 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14066 39352 14130 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14066 39271 14130 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14066 39190 14130 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14066 39109 14130 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14066 39028 14130 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 38959 14118 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 38879 14118 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 38799 14118 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 38719 14118 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 38639 14118 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 38559 14118 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 38479 14118 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 38399 14118 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 38319 14118 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 38239 14118 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 38159 14118 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 38079 14118 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 37999 14118 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 37919 14118 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 37839 14118 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 37759 14118 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 37679 14118 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 37599 14118 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 37519 14118 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 37439 14118 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 37359 14118 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 37279 14118 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 37199 14118 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 37119 14118 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 37039 14118 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 36959 14118 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 36879 14118 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 36799 14118 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 36719 14118 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 36639 14118 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 36559 14118 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 36479 14118 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 36399 14118 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 36319 14118 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 36239 14118 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 36159 14118 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 36079 14118 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 35999 14118 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 35919 14118 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 35839 14118 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 35759 14118 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 35679 14118 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 35599 14118 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 35519 14118 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 35439 14118 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 35359 14118 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 35279 14118 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 35199 14118 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14071 6042 14111 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14071 5956 14111 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14071 5870 14111 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14071 5784 14111 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14071 5698 14111 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14071 5612 14111 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14071 5526 14111 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14071 5440 14111 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14071 5354 14111 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14071 5268 14111 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14071 5182 14111 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13986 39919 14050 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13986 39838 14050 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13986 39757 14050 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13986 39676 14050 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13986 39595 14050 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13986 39514 14050 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13986 39433 14050 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13986 39352 14050 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13986 39271 14050 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13986 39190 14050 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13986 39109 14050 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13986 39028 14050 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 38959 14038 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 38879 14038 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 38799 14038 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 38719 14038 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 38639 14038 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 38559 14038 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 38479 14038 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 38399 14038 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 38319 14038 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 38239 14038 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 38159 14038 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 38079 14038 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 37999 14038 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 37919 14038 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 37839 14038 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 37759 14038 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 37679 14038 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 37599 14038 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 37519 14038 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 37439 14038 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 37359 14038 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 37279 14038 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 37199 14038 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 37119 14038 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 37039 14038 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 36959 14038 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 36879 14038 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 36799 14038 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 36719 14038 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 36639 14038 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 36559 14038 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 36479 14038 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 36399 14038 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 36319 14038 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 36239 14038 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 36159 14038 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 36079 14038 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 35999 14038 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 35919 14038 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 35839 14038 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 35759 14038 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 35679 14038 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 35599 14038 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 35519 14038 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 35439 14038 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 35359 14038 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 35279 14038 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 35199 14038 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13990 6042 14030 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13990 5956 14030 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13990 5870 14030 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13990 5784 14030 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13990 5698 14030 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13990 5612 14030 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13990 5526 14030 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13990 5440 14030 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13990 5354 14030 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13990 5268 14030 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13990 5182 14030 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13906 39919 13970 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13906 39838 13970 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13906 39757 13970 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13906 39676 13970 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13906 39595 13970 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13906 39514 13970 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13906 39433 13970 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13906 39352 13970 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13906 39271 13970 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13906 39190 13970 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13906 39109 13970 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13906 39028 13970 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 38959 13958 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 38879 13958 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 38799 13958 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 38719 13958 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 38639 13958 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 38559 13958 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 38479 13958 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 38399 13958 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 38319 13958 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 38239 13958 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 38159 13958 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 38079 13958 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 37999 13958 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 37919 13958 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 37839 13958 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 37759 13958 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 37679 13958 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 37599 13958 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 37519 13958 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 37439 13958 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 37359 13958 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 37279 13958 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 37199 13958 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 37119 13958 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 37039 13958 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 36959 13958 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 36879 13958 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 36799 13958 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 36719 13958 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 36639 13958 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 36559 13958 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 36479 13958 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 36399 13958 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 36319 13958 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 36239 13958 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 36159 13958 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 36079 13958 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 35999 13958 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 35919 13958 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 35839 13958 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 35759 13958 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 35679 13958 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 35599 13958 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 35519 13958 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 35439 13958 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 35359 13958 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 35279 13958 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 35199 13958 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 6042 13949 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5956 13949 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5870 13949 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5784 13949 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5698 13949 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5612 13949 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5526 13949 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5440 13949 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5354 13949 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5268 13949 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5182 13949 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13826 39919 13890 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13826 39838 13890 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13826 39757 13890 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13826 39676 13890 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13826 39595 13890 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13826 39514 13890 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13826 39433 13890 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13826 39352 13890 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13826 39271 13890 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13826 39190 13890 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13826 39109 13890 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13826 39028 13890 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 38959 13878 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 38879 13878 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 38799 13878 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 38719 13878 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 38639 13878 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 38559 13878 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 38479 13878 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 38399 13878 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 38319 13878 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 38239 13878 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 38159 13878 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 38079 13878 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 37999 13878 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 37919 13878 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 37839 13878 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 37759 13878 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 37679 13878 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 37599 13878 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 37519 13878 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 37439 13878 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 37359 13878 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 37279 13878 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 37199 13878 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 37119 13878 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 37039 13878 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 36959 13878 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 36879 13878 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 36799 13878 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 36719 13878 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 36639 13878 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 36559 13878 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 36479 13878 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 36399 13878 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 36319 13878 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 36239 13878 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 36159 13878 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 36079 13878 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 35999 13878 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 35919 13878 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 35839 13878 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 35759 13878 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 35679 13878 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 35599 13878 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 35519 13878 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 35439 13878 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 35359 13878 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 35279 13878 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 35199 13878 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13828 6042 13868 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13828 5956 13868 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13828 5870 13868 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13828 5784 13868 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13828 5698 13868 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13828 5612 13868 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13828 5526 13868 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13828 5440 13868 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13828 5354 13868 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13828 5268 13868 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13828 5182 13868 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13746 39919 13810 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13746 39838 13810 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13746 39757 13810 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13746 39676 13810 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13746 39595 13810 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13746 39514 13810 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13746 39433 13810 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13746 39352 13810 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13746 39271 13810 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13746 39190 13810 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13746 39109 13810 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13746 39028 13810 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 38959 13798 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 38879 13798 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 38799 13798 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 38719 13798 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 38639 13798 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 38559 13798 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 38479 13798 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 38399 13798 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 38319 13798 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 38239 13798 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 38159 13798 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 38079 13798 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 37999 13798 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 37919 13798 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 37839 13798 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 37759 13798 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 37679 13798 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 37599 13798 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 37519 13798 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 37439 13798 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 37359 13798 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 37279 13798 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 37199 13798 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 37119 13798 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 37039 13798 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 36959 13798 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 36879 13798 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 36799 13798 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 36719 13798 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 36639 13798 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 36559 13798 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 36479 13798 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 36399 13798 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 36319 13798 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 36239 13798 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 36159 13798 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 36079 13798 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 35999 13798 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 35919 13798 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 35839 13798 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 35759 13798 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 35679 13798 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 35599 13798 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 35519 13798 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 35439 13798 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 35359 13798 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 35279 13798 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 35199 13798 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13747 6042 13787 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13747 5956 13787 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13747 5870 13787 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13747 5784 13787 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13747 5698 13787 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13747 5612 13787 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13747 5526 13787 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13747 5440 13787 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13747 5354 13787 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13747 5268 13787 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13747 5182 13787 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 39919 13730 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 39838 13730 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 39757 13730 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 39676 13730 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 39595 13730 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 39514 13730 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 39433 13730 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 39352 13730 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 39271 13730 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 39190 13730 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 39109 13730 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 39028 13730 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 38959 13718 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 38879 13718 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 38799 13718 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 38719 13718 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 38639 13718 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 38559 13718 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 38479 13718 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 38399 13718 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 38319 13718 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 38239 13718 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 38159 13718 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 38079 13718 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 37999 13718 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 37919 13718 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 37839 13718 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 37759 13718 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 37679 13718 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 37599 13718 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 37519 13718 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 37439 13718 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 37359 13718 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 37279 13718 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 37199 13718 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 37119 13718 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 37039 13718 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 36959 13718 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 36879 13718 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 36799 13718 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 36719 13718 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 36639 13718 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 36559 13718 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 36479 13718 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 36399 13718 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 36319 13718 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 36239 13718 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 36159 13718 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 36079 13718 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 35999 13718 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 35919 13718 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 35839 13718 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 35759 13718 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 35679 13718 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 35599 13718 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 35519 13718 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 35439 13718 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 35359 13718 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 35279 13718 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 35199 13718 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 6042 13706 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 5956 13706 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 5870 13706 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 5784 13706 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 5698 13706 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 5612 13706 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 5526 13706 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 5440 13706 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 5354 13706 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 5268 13706 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 5182 13706 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13586 39919 13650 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13586 39838 13650 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13586 39757 13650 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13586 39676 13650 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13586 39595 13650 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13586 39514 13650 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13586 39433 13650 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13586 39352 13650 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13586 39271 13650 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13586 39190 13650 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13586 39109 13650 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13586 39028 13650 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 38959 13638 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 38879 13638 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 38799 13638 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 38719 13638 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 38639 13638 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 38559 13638 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 38479 13638 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 38399 13638 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 38319 13638 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 38239 13638 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 38159 13638 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 38079 13638 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 37999 13638 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 37919 13638 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 37839 13638 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 37759 13638 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 37679 13638 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 37599 13638 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 37519 13638 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 37439 13638 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 37359 13638 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 37279 13638 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 37199 13638 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 37119 13638 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 37039 13638 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 36959 13638 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 36879 13638 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 36799 13638 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 36719 13638 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 36639 13638 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 36559 13638 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 36479 13638 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 36399 13638 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 36319 13638 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 36239 13638 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 36159 13638 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 36079 13638 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 35999 13638 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 35919 13638 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 35839 13638 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 35759 13638 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 35679 13638 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 35599 13638 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 35519 13638 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 35439 13638 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 35359 13638 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 35279 13638 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 35199 13638 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 6042 13625 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5956 13625 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5870 13625 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5784 13625 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5698 13625 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5612 13625 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5526 13625 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5440 13625 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5354 13625 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5268 13625 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5182 13625 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13506 39919 13570 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13506 39838 13570 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13506 39757 13570 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13506 39676 13570 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13506 39595 13570 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13506 39514 13570 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13506 39433 13570 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13506 39352 13570 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13506 39271 13570 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13506 39190 13570 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13506 39109 13570 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13506 39028 13570 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 38959 13558 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 38879 13558 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 38799 13558 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 38719 13558 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 38639 13558 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 38559 13558 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 38479 13558 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 38399 13558 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 38319 13558 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 38239 13558 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 38159 13558 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 38079 13558 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 37999 13558 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 37919 13558 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 37839 13558 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 37759 13558 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 37679 13558 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 37599 13558 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 37519 13558 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 37439 13558 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 37359 13558 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 37279 13558 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 37199 13558 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 37119 13558 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 37039 13558 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 36959 13558 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 36879 13558 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 36799 13558 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 36719 13558 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 36639 13558 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 36559 13558 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 36479 13558 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 36399 13558 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 36319 13558 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 36239 13558 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 36159 13558 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 36079 13558 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 35999 13558 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 35919 13558 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 35839 13558 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 35759 13558 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 35679 13558 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 35599 13558 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 35519 13558 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 35439 13558 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 35359 13558 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 35279 13558 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 35199 13558 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13504 6042 13544 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13504 5956 13544 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13504 5870 13544 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13504 5784 13544 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13504 5698 13544 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13504 5612 13544 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13504 5526 13544 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13504 5440 13544 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13504 5354 13544 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13504 5268 13544 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13504 5182 13544 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13426 39919 13490 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13426 39838 13490 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13426 39757 13490 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13426 39676 13490 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13426 39595 13490 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13426 39514 13490 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13426 39433 13490 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13426 39352 13490 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13426 39271 13490 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13426 39190 13490 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13426 39109 13490 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13426 39028 13490 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 38959 13478 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 38879 13478 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 38799 13478 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 38719 13478 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 38639 13478 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 38559 13478 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 38479 13478 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 38399 13478 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 38319 13478 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 38239 13478 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 38159 13478 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 38079 13478 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 37999 13478 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 37919 13478 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 37839 13478 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 37759 13478 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 37679 13478 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 37599 13478 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 37519 13478 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 37439 13478 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 37359 13478 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 37279 13478 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 37199 13478 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 37119 13478 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 37039 13478 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 36959 13478 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 36879 13478 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 36799 13478 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 36719 13478 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 36639 13478 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 36559 13478 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 36479 13478 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 36399 13478 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 36319 13478 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 36239 13478 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 36159 13478 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 36079 13478 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 35999 13478 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 35919 13478 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 35839 13478 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 35759 13478 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 35679 13478 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 35599 13478 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 35519 13478 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 35439 13478 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 35359 13478 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 35279 13478 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 35199 13478 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13423 6042 13463 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13423 5956 13463 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13423 5870 13463 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13423 5784 13463 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13423 5698 13463 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13423 5612 13463 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13423 5526 13463 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13423 5440 13463 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13423 5354 13463 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13423 5268 13463 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13423 5182 13463 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13346 39919 13410 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13346 39838 13410 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13346 39757 13410 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13346 39676 13410 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13346 39595 13410 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13346 39514 13410 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13346 39433 13410 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13346 39352 13410 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13346 39271 13410 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13346 39190 13410 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13346 39109 13410 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13346 39028 13410 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 38959 13398 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 38879 13398 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 38799 13398 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 38719 13398 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 38639 13398 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 38559 13398 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 38479 13398 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 38399 13398 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 38319 13398 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 38239 13398 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 38159 13398 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 38079 13398 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 37999 13398 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 37919 13398 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 37839 13398 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 37759 13398 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 37679 13398 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 37599 13398 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 37519 13398 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 37439 13398 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 37359 13398 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 37279 13398 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 37199 13398 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 37119 13398 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 37039 13398 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 36959 13398 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 36879 13398 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 36799 13398 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 36719 13398 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 36639 13398 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 36559 13398 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 36479 13398 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 36399 13398 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 36319 13398 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 36239 13398 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 36159 13398 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 36079 13398 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 35999 13398 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 35919 13398 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 35839 13398 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 35759 13398 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 35679 13398 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 35599 13398 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 35519 13398 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 35439 13398 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 35359 13398 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 35279 13398 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 35199 13398 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13342 6042 13382 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13342 5956 13382 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13342 5870 13382 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13342 5784 13382 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13342 5698 13382 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13342 5612 13382 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13342 5526 13382 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13342 5440 13382 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13342 5354 13382 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13342 5268 13382 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13342 5182 13382 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13266 39919 13330 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13266 39838 13330 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13266 39757 13330 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13266 39676 13330 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13266 39595 13330 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13266 39514 13330 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13266 39433 13330 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13266 39352 13330 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13266 39271 13330 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13266 39190 13330 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13266 39109 13330 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13266 39028 13330 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 38959 13318 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 38879 13318 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 38799 13318 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 38719 13318 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 38639 13318 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 38559 13318 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 38479 13318 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 38399 13318 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 38319 13318 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 38239 13318 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 38159 13318 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 38079 13318 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 37999 13318 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 37919 13318 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 37839 13318 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 37759 13318 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 37679 13318 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 37599 13318 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 37519 13318 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 37439 13318 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 37359 13318 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 37279 13318 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 37199 13318 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 37119 13318 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 37039 13318 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 36959 13318 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 36879 13318 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 36799 13318 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 36719 13318 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 36639 13318 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 36559 13318 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 36479 13318 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 36399 13318 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 36319 13318 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 36239 13318 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 36159 13318 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 36079 13318 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 35999 13318 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 35919 13318 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 35839 13318 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 35759 13318 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 35679 13318 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 35599 13318 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 35519 13318 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 35439 13318 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 35359 13318 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 35279 13318 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 35199 13318 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 6042 13301 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5956 13301 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5870 13301 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5784 13301 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5698 13301 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5612 13301 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5526 13301 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5440 13301 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5354 13301 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5268 13301 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5182 13301 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13186 39919 13250 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13186 39838 13250 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13186 39757 13250 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13186 39676 13250 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13186 39595 13250 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13186 39514 13250 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13186 39433 13250 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13186 39352 13250 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13186 39271 13250 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13186 39190 13250 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13186 39109 13250 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13186 39028 13250 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 38959 13238 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 38879 13238 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 38799 13238 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 38719 13238 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 38639 13238 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 38559 13238 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 38479 13238 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 38399 13238 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 38319 13238 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 38239 13238 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 38159 13238 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 38079 13238 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 37999 13238 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 37919 13238 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 37839 13238 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 37759 13238 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 37679 13238 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 37599 13238 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 37519 13238 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 37439 13238 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 37359 13238 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 37279 13238 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 37199 13238 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 37119 13238 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 37039 13238 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 36959 13238 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 36879 13238 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 36799 13238 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 36719 13238 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 36639 13238 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 36559 13238 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 36479 13238 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 36399 13238 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 36319 13238 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 36239 13238 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 36159 13238 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 36079 13238 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 35999 13238 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 35919 13238 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 35839 13238 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 35759 13238 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 35679 13238 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 35599 13238 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 35519 13238 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 35439 13238 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 35359 13238 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 35279 13238 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 35199 13238 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13180 6042 13220 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13180 5956 13220 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13180 5870 13220 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13180 5784 13220 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13180 5698 13220 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13180 5612 13220 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13180 5526 13220 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13180 5440 13220 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13180 5354 13220 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13180 5268 13220 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13180 5182 13220 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13106 39919 13170 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13106 39838 13170 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13106 39757 13170 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13106 39676 13170 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13106 39595 13170 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13106 39514 13170 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13106 39433 13170 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13106 39352 13170 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13106 39271 13170 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13106 39190 13170 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13106 39109 13170 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13106 39028 13170 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 38959 13158 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 38879 13158 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 38799 13158 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 38719 13158 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 38639 13158 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 38559 13158 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 38479 13158 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 38399 13158 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 38319 13158 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 38239 13158 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 38159 13158 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 38079 13158 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 37999 13158 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 37919 13158 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 37839 13158 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 37759 13158 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 37679 13158 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 37599 13158 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 37519 13158 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 37439 13158 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 37359 13158 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 37279 13158 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 37199 13158 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 37119 13158 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 37039 13158 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 36959 13158 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 36879 13158 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 36799 13158 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 36719 13158 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 36639 13158 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 36559 13158 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 36479 13158 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 36399 13158 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 36319 13158 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 36239 13158 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 36159 13158 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 36079 13158 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 35999 13158 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 35919 13158 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 35839 13158 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 35759 13158 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 35679 13158 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 35599 13158 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 35519 13158 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 35439 13158 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 35359 13158 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 35279 13158 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 35199 13158 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13099 6042 13139 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13099 5956 13139 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13099 5870 13139 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13099 5784 13139 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13099 5698 13139 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13099 5612 13139 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13099 5526 13139 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13099 5440 13139 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13099 5354 13139 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13099 5268 13139 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13099 5182 13139 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13026 39919 13090 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13026 39838 13090 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13026 39757 13090 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13026 39676 13090 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13026 39595 13090 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13026 39514 13090 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13026 39433 13090 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13026 39352 13090 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13026 39271 13090 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13026 39190 13090 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13026 39109 13090 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13026 39028 13090 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 38959 13078 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 38879 13078 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 38799 13078 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 38719 13078 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 38639 13078 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 38559 13078 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 38479 13078 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 38399 13078 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 38319 13078 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 38239 13078 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 38159 13078 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 38079 13078 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 37999 13078 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 37919 13078 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 37839 13078 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 37759 13078 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 37679 13078 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 37599 13078 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 37519 13078 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 37439 13078 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 37359 13078 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 37279 13078 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 37199 13078 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 37119 13078 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 37039 13078 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 36959 13078 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 36879 13078 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 36799 13078 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 36719 13078 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 36639 13078 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 36559 13078 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 36479 13078 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 36399 13078 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 36319 13078 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 36239 13078 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 36159 13078 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 36079 13078 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 35999 13078 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 35919 13078 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 35839 13078 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 35759 13078 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 35679 13078 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 35599 13078 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 35519 13078 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 35439 13078 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 35359 13078 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 35279 13078 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 35199 13078 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13018 6042 13058 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13018 5956 13058 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13018 5870 13058 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13018 5784 13058 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13018 5698 13058 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13018 5612 13058 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13018 5526 13058 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13018 5440 13058 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13018 5354 13058 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13018 5268 13058 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13018 5182 13058 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12946 39919 13010 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12946 39838 13010 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12946 39757 13010 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12946 39676 13010 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12946 39595 13010 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12946 39514 13010 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12946 39433 13010 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12946 39352 13010 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12946 39271 13010 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12946 39190 13010 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12946 39109 13010 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12946 39028 13010 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 38959 12998 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 38879 12998 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 38799 12998 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 38719 12998 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 38639 12998 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 38559 12998 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 38479 12998 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 38399 12998 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 38319 12998 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 38239 12998 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 38159 12998 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 38079 12998 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 37999 12998 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 37919 12998 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 37839 12998 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 37759 12998 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 37679 12998 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 37599 12998 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 37519 12998 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 37439 12998 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 37359 12998 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 37279 12998 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 37199 12998 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 37119 12998 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 37039 12998 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 36959 12998 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 36879 12998 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 36799 12998 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 36719 12998 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 36639 12998 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 36559 12998 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 36479 12998 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 36399 12998 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 36319 12998 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 36239 12998 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 36159 12998 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 36079 12998 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 35999 12998 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 35919 12998 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 35839 12998 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 35759 12998 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 35679 12998 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 35599 12998 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 35519 12998 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 35439 12998 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 35359 12998 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 35279 12998 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 35199 12998 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 6042 12977 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5956 12977 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5870 12977 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5784 12977 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5698 12977 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5612 12977 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5526 12977 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5440 12977 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5354 12977 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5268 12977 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5182 12977 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12866 39919 12930 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12866 39838 12930 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12866 39757 12930 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12866 39676 12930 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12866 39595 12930 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12866 39514 12930 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12866 39433 12930 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12866 39352 12930 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12866 39271 12930 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12866 39190 12930 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12866 39109 12930 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12866 39028 12930 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 38959 12918 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 38879 12918 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 38799 12918 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 38719 12918 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 38639 12918 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 38559 12918 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 38479 12918 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 38399 12918 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 38319 12918 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 38239 12918 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 38159 12918 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 38079 12918 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 37999 12918 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 37919 12918 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 37839 12918 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 37759 12918 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 37679 12918 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 37599 12918 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 37519 12918 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 37439 12918 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 37359 12918 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 37279 12918 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 37199 12918 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 37119 12918 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 37039 12918 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 36959 12918 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 36879 12918 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 36799 12918 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 36719 12918 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 36639 12918 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 36559 12918 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 36479 12918 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 36399 12918 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 36319 12918 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 36239 12918 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 36159 12918 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 36079 12918 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 35999 12918 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 35919 12918 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 35839 12918 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 35759 12918 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 35679 12918 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 35599 12918 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 35519 12918 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 35439 12918 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 35359 12918 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 35279 12918 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 35199 12918 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12856 6042 12896 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12856 5956 12896 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12856 5870 12896 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12856 5784 12896 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12856 5698 12896 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12856 5612 12896 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12856 5526 12896 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12856 5440 12896 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12856 5354 12896 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12856 5268 12896 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12856 5182 12896 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12786 39919 12850 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12786 39838 12850 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12786 39757 12850 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12786 39676 12850 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12786 39595 12850 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12786 39514 12850 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12786 39433 12850 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12786 39352 12850 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12786 39271 12850 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12786 39190 12850 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12786 39109 12850 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12786 39028 12850 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 38959 12838 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 38879 12838 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 38799 12838 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 38719 12838 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 38639 12838 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 38559 12838 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 38479 12838 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 38399 12838 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 38319 12838 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 38239 12838 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 38159 12838 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 38079 12838 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 37999 12838 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 37919 12838 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 37839 12838 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 37759 12838 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 37679 12838 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 37599 12838 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 37519 12838 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 37439 12838 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 37359 12838 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 37279 12838 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 37199 12838 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 37119 12838 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 37039 12838 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 36959 12838 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 36879 12838 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 36799 12838 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 36719 12838 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 36639 12838 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 36559 12838 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 36479 12838 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 36399 12838 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 36319 12838 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 36239 12838 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 36159 12838 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 36079 12838 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 35999 12838 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 35919 12838 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 35839 12838 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 35759 12838 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 35679 12838 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 35599 12838 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 35519 12838 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 35439 12838 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 35359 12838 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 35279 12838 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 35199 12838 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12775 6042 12815 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12775 5956 12815 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12775 5870 12815 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12775 5784 12815 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12775 5698 12815 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12775 5612 12815 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12775 5526 12815 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12775 5440 12815 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12775 5354 12815 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12775 5268 12815 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12775 5182 12815 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12706 39919 12770 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12706 39838 12770 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12706 39757 12770 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12706 39676 12770 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12706 39595 12770 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12706 39514 12770 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12706 39433 12770 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12706 39352 12770 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12706 39271 12770 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12706 39190 12770 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12706 39109 12770 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12706 39028 12770 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 38959 12758 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 38879 12758 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 38799 12758 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 38719 12758 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 38639 12758 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 38559 12758 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 38479 12758 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 38399 12758 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 38319 12758 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 38239 12758 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 38159 12758 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 38079 12758 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 37999 12758 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 37919 12758 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 37839 12758 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 37759 12758 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 37679 12758 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 37599 12758 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 37519 12758 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 37439 12758 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 37359 12758 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 37279 12758 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 37199 12758 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 37119 12758 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 37039 12758 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 36959 12758 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 36879 12758 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 36799 12758 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 36719 12758 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 36639 12758 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 36559 12758 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 36479 12758 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 36399 12758 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 36319 12758 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 36239 12758 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 36159 12758 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 36079 12758 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 35999 12758 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 35919 12758 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 35839 12758 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 35759 12758 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 35679 12758 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 35599 12758 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 35519 12758 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 35439 12758 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 35359 12758 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 35279 12758 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 35199 12758 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12694 6042 12734 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12694 5956 12734 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12694 5870 12734 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12694 5784 12734 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12694 5698 12734 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12694 5612 12734 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12694 5526 12734 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12694 5440 12734 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12694 5354 12734 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12694 5268 12734 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12694 5182 12734 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12626 39919 12690 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12626 39838 12690 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12626 39757 12690 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12626 39676 12690 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12626 39595 12690 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12626 39514 12690 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12626 39433 12690 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12626 39352 12690 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12626 39271 12690 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12626 39190 12690 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12626 39109 12690 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12626 39028 12690 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 38959 12678 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 38879 12678 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 38799 12678 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 38719 12678 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 38639 12678 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 38559 12678 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 38479 12678 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 38399 12678 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 38319 12678 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 38239 12678 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 38159 12678 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 38079 12678 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 37999 12678 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 37919 12678 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 37839 12678 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 37759 12678 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 37679 12678 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 37599 12678 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 37519 12678 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 37439 12678 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 37359 12678 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 37279 12678 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 37199 12678 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 37119 12678 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 37039 12678 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 36959 12678 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 36879 12678 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 36799 12678 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 36719 12678 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 36639 12678 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 36559 12678 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 36479 12678 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 36399 12678 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 36319 12678 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 36239 12678 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 36159 12678 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 36079 12678 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 35999 12678 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 35919 12678 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 35839 12678 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 35759 12678 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 35679 12678 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 35599 12678 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 35519 12678 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 35439 12678 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 35359 12678 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 35279 12678 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 35199 12678 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 6042 12653 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5956 12653 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5870 12653 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5784 12653 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5698 12653 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5612 12653 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5526 12653 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5440 12653 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5354 12653 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5268 12653 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5182 12653 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12546 39919 12610 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12546 39838 12610 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12546 39757 12610 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12546 39676 12610 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12546 39595 12610 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12546 39514 12610 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12546 39433 12610 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12546 39352 12610 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12546 39271 12610 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12546 39190 12610 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12546 39109 12610 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12546 39028 12610 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 38959 12598 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 38879 12598 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 38799 12598 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 38719 12598 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 38639 12598 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 38559 12598 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 38479 12598 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 38399 12598 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 38319 12598 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 38239 12598 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 38159 12598 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 38079 12598 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 37999 12598 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 37919 12598 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 37839 12598 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 37759 12598 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 37679 12598 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 37599 12598 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 37519 12598 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 37439 12598 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 37359 12598 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 37279 12598 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 37199 12598 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 37119 12598 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 37039 12598 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 36959 12598 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 36879 12598 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 36799 12598 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 36719 12598 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 36639 12598 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 36559 12598 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 36479 12598 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 36399 12598 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 36319 12598 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 36239 12598 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 36159 12598 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 36079 12598 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 35999 12598 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 35919 12598 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 35839 12598 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 35759 12598 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 35679 12598 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 35599 12598 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 35519 12598 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 35439 12598 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 35359 12598 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 35279 12598 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 35199 12598 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12532 6042 12572 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12532 5956 12572 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12532 5870 12572 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12532 5784 12572 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12532 5698 12572 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12532 5612 12572 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12532 5526 12572 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12532 5440 12572 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12532 5354 12572 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12532 5268 12572 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12532 5182 12572 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12466 39919 12530 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12466 39838 12530 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12466 39757 12530 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12466 39676 12530 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12466 39595 12530 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12466 39514 12530 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12466 39433 12530 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12466 39352 12530 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12466 39271 12530 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12466 39190 12530 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12466 39109 12530 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12466 39028 12530 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 38959 12518 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 38879 12518 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 38799 12518 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 38719 12518 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 38639 12518 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 38559 12518 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 38479 12518 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 38399 12518 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 38319 12518 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 38239 12518 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 38159 12518 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 38079 12518 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 37999 12518 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 37919 12518 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 37839 12518 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 37759 12518 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 37679 12518 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 37599 12518 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 37519 12518 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 37439 12518 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 37359 12518 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 37279 12518 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 37199 12518 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 37119 12518 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 37039 12518 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 36959 12518 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 36879 12518 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 36799 12518 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 36719 12518 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 36639 12518 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 36559 12518 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 36479 12518 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 36399 12518 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 36319 12518 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 36239 12518 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 36159 12518 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 36079 12518 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 35999 12518 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 35919 12518 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 35839 12518 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 35759 12518 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 35679 12518 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 35599 12518 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 35519 12518 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 35439 12518 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 35359 12518 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 35279 12518 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 35199 12518 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12451 6042 12491 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12451 5956 12491 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12451 5870 12491 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12451 5784 12491 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12451 5698 12491 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12451 5612 12491 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12451 5526 12491 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12451 5440 12491 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12451 5354 12491 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12451 5268 12491 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12451 5182 12491 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12386 39919 12450 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12386 39838 12450 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12386 39757 12450 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12386 39676 12450 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12386 39595 12450 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12386 39514 12450 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12386 39433 12450 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12386 39352 12450 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12386 39271 12450 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12386 39190 12450 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12386 39109 12450 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12386 39028 12450 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 38959 12438 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 38879 12438 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 38799 12438 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 38719 12438 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 38639 12438 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 38559 12438 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 38479 12438 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 38399 12438 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 38319 12438 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 38239 12438 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 38159 12438 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 38079 12438 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 37999 12438 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 37919 12438 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 37839 12438 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 37759 12438 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 37679 12438 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 37599 12438 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 37519 12438 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 37439 12438 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 37359 12438 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 37279 12438 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 37199 12438 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 37119 12438 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 37039 12438 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 36959 12438 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 36879 12438 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 36799 12438 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 36719 12438 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 36639 12438 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 36559 12438 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 36479 12438 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 36399 12438 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 36319 12438 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 36239 12438 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 36159 12438 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 36079 12438 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 35999 12438 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 35919 12438 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 35839 12438 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 35759 12438 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 35679 12438 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 35599 12438 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 35519 12438 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 35439 12438 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 35359 12438 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 35279 12438 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 35199 12438 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12370 6042 12410 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12370 5956 12410 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12370 5870 12410 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12370 5784 12410 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12370 5698 12410 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12370 5612 12410 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12370 5526 12410 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12370 5440 12410 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12370 5354 12410 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12370 5268 12410 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12370 5182 12410 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12306 39919 12370 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12306 39838 12370 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12306 39757 12370 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12306 39676 12370 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12306 39595 12370 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12306 39514 12370 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12306 39433 12370 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12306 39352 12370 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12306 39271 12370 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12306 39190 12370 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12306 39109 12370 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12306 39028 12370 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 38959 12358 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 38879 12358 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 38799 12358 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 38719 12358 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 38639 12358 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 38559 12358 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 38479 12358 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 38399 12358 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 38319 12358 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 38239 12358 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 38159 12358 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 38079 12358 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 37999 12358 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 37919 12358 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 37839 12358 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 37759 12358 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 37679 12358 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 37599 12358 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 37519 12358 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 37439 12358 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 37359 12358 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 37279 12358 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 37199 12358 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 37119 12358 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 37039 12358 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 36959 12358 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 36879 12358 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 36799 12358 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 36719 12358 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 36639 12358 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 36559 12358 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 36479 12358 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 36399 12358 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 36319 12358 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 36239 12358 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 36159 12358 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 36079 12358 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 35999 12358 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 35919 12358 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 35839 12358 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 35759 12358 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 35679 12358 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 35599 12358 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 35519 12358 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 35439 12358 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 35359 12358 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 35279 12358 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 35199 12358 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 6042 12329 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5956 12329 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5870 12329 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5784 12329 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5698 12329 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5612 12329 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5526 12329 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5440 12329 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5354 12329 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5268 12329 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5182 12329 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7417 39438 12264 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12212 39850 12252 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12212 39770 12252 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12212 39690 12252 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12212 39610 12252 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12212 39530 12252 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12212 39450 12252 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12208 6042 12248 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12208 5956 12248 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12208 5870 12248 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12208 5784 12248 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12208 5698 12248 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12208 5612 12248 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12208 5526 12248 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12208 5440 12248 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12208 5354 12248 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12208 5268 12248 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12208 5182 12248 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12170 39329 12234 39393 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12170 39247 12234 39311 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12132 39930 12172 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12132 39850 12172 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12132 39770 12172 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12132 39690 12172 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12132 39610 12172 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12132 39530 12172 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12132 39450 12172 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12127 6042 12167 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12127 5956 12167 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12127 5870 12167 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12127 5784 12167 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12127 5698 12167 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12127 5612 12167 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12127 5526 12167 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12127 5440 12167 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12127 5354 12167 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12127 5268 12167 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12127 5182 12167 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12052 39930 12092 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12052 39850 12092 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12052 39770 12092 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12052 39690 12092 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12052 39610 12092 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12052 39530 12092 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12052 39450 12092 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12046 6042 12086 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12046 5956 12086 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12046 5870 12086 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12046 5784 12086 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12046 5698 12086 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12046 5612 12086 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12046 5526 12086 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12046 5440 12086 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12046 5354 12086 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12046 5268 12086 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12046 5182 12086 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11972 39930 12012 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11972 39850 12012 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11972 39770 12012 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11972 39690 12012 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11972 39610 12012 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11972 39530 12012 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11972 39450 12012 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 6042 12005 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5956 12005 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5870 12005 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5784 12005 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5698 12005 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5612 12005 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5526 12005 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5440 12005 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5354 12005 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5268 12005 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5182 12005 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11892 39930 11932 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11892 39850 11932 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11892 39770 11932 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11892 39690 11932 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11892 39610 11932 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11892 39530 11932 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11892 39450 11932 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11884 6042 11924 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11884 5956 11924 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11884 5870 11924 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11884 5784 11924 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11884 5698 11924 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11884 5612 11924 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11884 5526 11924 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11884 5440 11924 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11884 5354 11924 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11884 5268 11924 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11884 5182 11924 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11812 39930 11852 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11812 39850 11852 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11812 39770 11852 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11812 39690 11852 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11812 39610 11852 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11812 39530 11852 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11812 39450 11852 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11803 6042 11843 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11803 5956 11843 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11803 5870 11843 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11803 5784 11843 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11803 5698 11843 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11803 5612 11843 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11803 5526 11843 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11803 5440 11843 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11803 5354 11843 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11803 5268 11843 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11803 5182 11843 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11732 39930 11772 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11732 39850 11772 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11732 39770 11772 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11732 39690 11772 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11732 39610 11772 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11732 39530 11772 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11732 39450 11772 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11722 6042 11762 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11722 5956 11762 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11722 5870 11762 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11722 5784 11762 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11722 5698 11762 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11722 5612 11762 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11722 5526 11762 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11722 5440 11762 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11722 5354 11762 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11722 5268 11762 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11722 5182 11762 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11652 39930 11692 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11652 39850 11692 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11652 39770 11692 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11652 39690 11692 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11652 39610 11692 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11652 39530 11692 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11652 39450 11692 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 6042 11681 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5956 11681 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5870 11681 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5784 11681 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5698 11681 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5612 11681 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5526 11681 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5440 11681 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5354 11681 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5268 11681 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5182 11681 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11572 39930 11612 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11572 39850 11612 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11572 39770 11612 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11572 39690 11612 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11572 39610 11612 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11572 39530 11612 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11572 39450 11612 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11560 6042 11600 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11560 5956 11600 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11560 5870 11600 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11560 5784 11600 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11560 5698 11600 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11560 5612 11600 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11560 5526 11600 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11560 5440 11600 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11560 5354 11600 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11560 5268 11600 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11560 5182 11600 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11492 39930 11532 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11492 39850 11532 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11492 39770 11532 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11492 39690 11532 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11492 39610 11532 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11492 39530 11532 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11492 39450 11532 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11479 6042 11519 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11479 5956 11519 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11479 5870 11519 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11479 5784 11519 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11479 5698 11519 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11479 5612 11519 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11479 5526 11519 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11479 5440 11519 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11479 5354 11519 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11479 5268 11519 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11479 5182 11519 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11412 39930 11452 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11412 39850 11452 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11412 39770 11452 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11412 39690 11452 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11412 39610 11452 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11412 39530 11452 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11412 39450 11452 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11398 6042 11438 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11398 5956 11438 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11398 5870 11438 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11398 5784 11438 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11398 5698 11438 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11398 5612 11438 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11398 5526 11438 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11398 5440 11438 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11398 5354 11438 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11398 5268 11438 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11398 5182 11438 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11332 39930 11372 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11332 39850 11372 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11332 39770 11372 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11332 39690 11372 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11332 39610 11372 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11332 39530 11372 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11332 39450 11372 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 6042 11357 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5956 11357 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5870 11357 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5784 11357 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5698 11357 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5612 11357 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5526 11357 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5440 11357 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5354 11357 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5268 11357 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5182 11357 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11252 39930 11292 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11252 39850 11292 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11252 39770 11292 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11252 39690 11292 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11252 39610 11292 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11252 39530 11292 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11252 39450 11292 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11236 6042 11276 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11236 5956 11276 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11236 5870 11276 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11236 5784 11276 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11236 5698 11276 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11236 5612 11276 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11236 5526 11276 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11236 5440 11276 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11236 5354 11276 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11236 5268 11276 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11236 5182 11276 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11172 39930 11212 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11172 39850 11212 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11172 39770 11212 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11172 39690 11212 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11172 39610 11212 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11172 39530 11212 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11172 39450 11212 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11155 6042 11195 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11155 5956 11195 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11155 5870 11195 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11155 5784 11195 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11155 5698 11195 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11155 5612 11195 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11155 5526 11195 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11155 5440 11195 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11155 5354 11195 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11155 5268 11195 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11155 5182 11195 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11092 39930 11132 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11092 39850 11132 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11092 39770 11132 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11092 39690 11132 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11092 39610 11132 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11092 39530 11132 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11092 39450 11132 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11074 6042 11114 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11074 5956 11114 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11074 5870 11114 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11074 5784 11114 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11074 5698 11114 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11074 5612 11114 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11074 5526 11114 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11074 5440 11114 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11074 5354 11114 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11074 5268 11114 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11074 5182 11114 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11012 39930 11052 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11012 39850 11052 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11012 39770 11052 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11012 39690 11052 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11012 39610 11052 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11012 39530 11052 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11012 39450 11052 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 6042 11033 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5956 11033 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5870 11033 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5784 11033 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5698 11033 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5612 11033 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5526 11033 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5440 11033 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5354 11033 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5268 11033 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5182 11033 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10932 39930 10972 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10932 39850 10972 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10932 39770 10972 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10932 39690 10972 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10932 39610 10972 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10932 39530 10972 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10932 39450 10972 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10912 6042 10952 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10912 5956 10952 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10912 5870 10952 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10912 5784 10952 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10912 5698 10952 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10912 5612 10952 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10912 5526 10952 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10912 5440 10952 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10912 5354 10952 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10912 5268 10952 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10912 5182 10952 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10852 39930 10892 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10852 39850 10892 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10852 39770 10892 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10852 39690 10892 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10852 39610 10892 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10852 39530 10892 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10852 39450 10892 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10831 6042 10871 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10831 5956 10871 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10831 5870 10871 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10831 5784 10871 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10831 5698 10871 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10831 5612 10871 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10831 5526 10871 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10831 5440 10871 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10831 5354 10871 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10831 5268 10871 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10831 5182 10871 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10772 39930 10812 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10772 39850 10812 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10772 39770 10812 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10772 39690 10812 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10772 39610 10812 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10772 39530 10812 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10772 39450 10812 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10750 6042 10790 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10750 5956 10790 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10750 5870 10790 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10750 5784 10790 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10750 5698 10790 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10750 5612 10790 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10750 5526 10790 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10750 5440 10790 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10750 5354 10790 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10750 5268 10790 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10750 5182 10790 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10692 39930 10732 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10692 39850 10732 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10692 39770 10732 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10692 39690 10732 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10692 39610 10732 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10692 39530 10732 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10692 39450 10732 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 6042 10709 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5956 10709 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5870 10709 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5784 10709 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5698 10709 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5612 10709 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5526 10709 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5440 10709 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5354 10709 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5268 10709 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5182 10709 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10612 39930 10652 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10612 39850 10652 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10612 39770 10652 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10612 39690 10652 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10612 39610 10652 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10612 39530 10652 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10612 39450 10652 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10588 6042 10628 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10588 5956 10628 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10588 5870 10628 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10588 5784 10628 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10588 5698 10628 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10588 5612 10628 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10588 5526 10628 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10588 5440 10628 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10588 5354 10628 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10588 5268 10628 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10588 5182 10628 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10532 39930 10572 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10532 39850 10572 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10532 39770 10572 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10532 39690 10572 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10532 39610 10572 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10532 39530 10572 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10532 39450 10572 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10506 6042 10546 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10506 5956 10546 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10506 5870 10546 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10506 5784 10546 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10506 5698 10546 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10506 5612 10546 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10506 5526 10546 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10506 5440 10546 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10506 5354 10546 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10506 5268 10546 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10506 5182 10546 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10452 39930 10492 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10452 39850 10492 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10452 39770 10492 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10452 39690 10492 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10452 39610 10492 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10452 39530 10492 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10452 39450 10492 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10424 6042 10464 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10424 5956 10464 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10424 5870 10464 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10424 5784 10464 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10424 5698 10464 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10424 5612 10464 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10424 5526 10464 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10424 5440 10464 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10424 5354 10464 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10424 5268 10464 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10424 5182 10464 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10372 39930 10412 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10372 39850 10412 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10372 39770 10412 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10372 39690 10412 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10372 39610 10412 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10372 39530 10412 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10372 39450 10412 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 6042 10382 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5956 10382 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5870 10382 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5784 10382 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5698 10382 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5612 10382 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5526 10382 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5440 10382 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5354 10382 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5268 10382 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5182 10382 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10292 39930 10332 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10292 39850 10332 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10292 39770 10332 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10292 39690 10332 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10292 39610 10332 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10292 39530 10332 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10292 39450 10332 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10260 6042 10300 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10260 5956 10300 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10260 5870 10300 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10260 5784 10300 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10260 5698 10300 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10260 5612 10300 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10260 5526 10300 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10260 5440 10300 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10260 5354 10300 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10260 5268 10300 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10260 5182 10300 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10212 39930 10252 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10212 39850 10252 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10212 39770 10252 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10212 39690 10252 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10212 39610 10252 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10212 39530 10252 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10212 39450 10252 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10178 6042 10218 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10178 5956 10218 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10178 5870 10218 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10178 5784 10218 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10178 5698 10218 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10178 5612 10218 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10178 5526 10218 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10178 5440 10218 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10178 5354 10218 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10178 5268 10218 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10178 5182 10218 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10132 39930 10172 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10132 39850 10172 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10132 39770 10172 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10132 39690 10172 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10132 39610 10172 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10132 39530 10172 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10132 39450 10172 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10096 6042 10136 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10096 5956 10136 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10096 5870 10136 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10096 5784 10136 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10096 5698 10136 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10096 5612 10136 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10096 5526 10136 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10096 5440 10136 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10096 5354 10136 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10096 5268 10136 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10096 5182 10136 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10052 39930 10092 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10052 39850 10092 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10052 39770 10092 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10052 39690 10092 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10052 39610 10092 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10052 39530 10092 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10052 39450 10092 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9972 39930 10012 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9972 39850 10012 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9972 39770 10012 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9972 39690 10012 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9972 39610 10012 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9972 39530 10012 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9972 39450 10012 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9892 39930 9932 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9892 39850 9932 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9892 39770 9932 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9892 39690 9932 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9892 39610 9932 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9892 39530 9932 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9892 39450 9932 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9812 39930 9852 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9812 39850 9852 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9812 39770 9852 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9812 39690 9852 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9812 39610 9852 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9812 39530 9852 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9812 39450 9852 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9732 39930 9772 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9732 39850 9772 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9732 39770 9772 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9732 39690 9772 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9732 39610 9772 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9732 39530 9772 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9732 39450 9772 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9652 39930 9692 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9652 39850 9692 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9652 39770 9692 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9652 39690 9692 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9652 39610 9692 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9652 39530 9692 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9652 39450 9692 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9572 39930 9612 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9572 39850 9612 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9572 39770 9612 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9572 39690 9612 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9572 39610 9612 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9572 39530 9612 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9572 39450 9612 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9492 39930 9532 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9492 39850 9532 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9492 39770 9532 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9492 39690 9532 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9492 39610 9532 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9492 39530 9532 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9492 39450 9532 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9412 39930 9452 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9412 39850 9452 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9412 39770 9452 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9412 39690 9452 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9412 39610 9452 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9412 39530 9452 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9412 39450 9452 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9332 39930 9372 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9332 39850 9372 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9332 39770 9372 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9332 39690 9372 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9332 39610 9372 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9332 39530 9372 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9332 39450 9372 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9252 39930 9292 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9252 39850 9292 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9252 39770 9292 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9252 39690 9292 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9252 39610 9292 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9252 39530 9292 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9252 39450 9292 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9172 39930 9212 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9172 39850 9212 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9172 39770 9212 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9172 39690 9212 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9172 39610 9212 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9172 39530 9212 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9172 39450 9212 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9092 39930 9132 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9092 39850 9132 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9092 39770 9132 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9092 39690 9132 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9092 39610 9132 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9092 39530 9132 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9092 39450 9132 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9012 39930 9052 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9012 39850 9052 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9012 39770 9052 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9012 39690 9052 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9012 39610 9052 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9012 39530 9052 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9012 39450 9052 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8932 39930 8972 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8932 39850 8972 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8932 39770 8972 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8932 39690 8972 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8932 39610 8972 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8932 39530 8972 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8932 39450 8972 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8852 39930 8892 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8852 39850 8892 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8852 39770 8892 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8852 39690 8892 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8852 39610 8892 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8852 39530 8892 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8852 39450 8892 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8772 39930 8812 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8772 39850 8812 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8772 39770 8812 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8772 39690 8812 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8772 39610 8812 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8772 39530 8812 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8772 39450 8812 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8692 39930 8732 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8692 39850 8732 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8692 39770 8732 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8692 39690 8732 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8692 39610 8732 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8692 39530 8732 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8692 39450 8732 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8612 39930 8652 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8612 39850 8652 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8612 39770 8652 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8612 39690 8652 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8612 39610 8652 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8612 39530 8652 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8612 39450 8652 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8532 39930 8572 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8532 39850 8572 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8532 39770 8572 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8532 39690 8572 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8532 39610 8572 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8532 39530 8572 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8532 39450 8572 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8452 39930 8492 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8452 39850 8492 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8452 39770 8492 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8452 39690 8492 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8452 39610 8492 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8452 39530 8492 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8452 39450 8492 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8372 39930 8412 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8372 39850 8412 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8372 39770 8412 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8372 39690 8412 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8372 39610 8412 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8372 39530 8412 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8372 39450 8412 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8292 39930 8332 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8292 39850 8332 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8292 39770 8332 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8292 39690 8332 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8292 39610 8332 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8292 39530 8332 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8292 39450 8332 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8212 39930 8252 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8212 39850 8252 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8212 39770 8252 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8212 39690 8252 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8212 39610 8252 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8212 39530 8252 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8212 39450 8252 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8132 39930 8172 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8132 39850 8172 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8132 39770 8172 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8132 39690 8172 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8132 39610 8172 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8132 39530 8172 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8132 39450 8172 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8052 39930 8092 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8052 39850 8092 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8052 39770 8092 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8052 39690 8092 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8052 39610 8092 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8052 39530 8092 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8052 39450 8092 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7972 39930 8012 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7972 39850 8012 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7972 39770 8012 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7972 39690 8012 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7972 39610 8012 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7972 39530 8012 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7972 39450 8012 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7892 39930 7932 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7892 39850 7932 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7892 39770 7932 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7892 39690 7932 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7892 39610 7932 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7892 39530 7932 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7892 39450 7932 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7812 39930 7852 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7812 39850 7852 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7812 39770 7852 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7812 39690 7852 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7812 39610 7852 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7812 39530 7852 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7812 39450 7852 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7732 39930 7772 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7732 39850 7772 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7732 39770 7772 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7732 39690 7772 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7732 39610 7772 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7732 39530 7772 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7732 39450 7772 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7652 39930 7692 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7652 39850 7692 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7652 39770 7692 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7652 39690 7692 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7652 39610 7692 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7652 39530 7692 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7652 39450 7692 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7572 39930 7612 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7572 39850 7612 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7572 39770 7612 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7572 39690 7612 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7572 39610 7612 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7572 39530 7612 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7572 39450 7612 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7492 39930 7532 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7492 39850 7532 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7492 39770 7532 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7492 39690 7532 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7492 39610 7532 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7492 39530 7532 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7492 39450 7532 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7412 39930 7452 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7412 39850 7452 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7412 39770 7452 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7412 39690 7452 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7412 39610 7452 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7412 39530 7452 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7412 39450 7452 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5400 39438 7412 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7332 39850 7372 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7332 39770 7372 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7332 39690 7372 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7332 39610 7372 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7332 39530 7372 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7332 39450 7372 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7252 39930 7292 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7252 39850 7292 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7252 39770 7292 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7252 39690 7292 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7252 39610 7292 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7252 39530 7292 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7252 39450 7292 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7172 39930 7212 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7172 39850 7212 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7172 39770 7212 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7172 39690 7212 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7172 39610 7212 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7172 39530 7212 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7172 39450 7212 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7092 39930 7132 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7092 39850 7132 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7092 39770 7132 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7092 39690 7132 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7092 39610 7132 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7092 39530 7132 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7092 39450 7132 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7012 39930 7052 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7012 39850 7052 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7012 39770 7052 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7012 39690 7052 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7012 39610 7052 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7012 39530 7052 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7012 39450 7052 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6932 39930 6972 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6932 39850 6972 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6932 39770 6972 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6932 39690 6972 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6932 39610 6972 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6932 39530 6972 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6932 39450 6972 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6852 39930 6892 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6852 39850 6892 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6852 39770 6892 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6852 39690 6892 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6852 39610 6892 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6852 39530 6892 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6852 39450 6892 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6772 39930 6812 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6772 39850 6812 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6772 39770 6812 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6772 39690 6812 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6772 39610 6812 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6772 39530 6812 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6772 39450 6812 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6692 39930 6732 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6692 39850 6732 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6692 39770 6732 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6692 39690 6732 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6692 39610 6732 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6692 39530 6732 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6692 39450 6732 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6612 39930 6652 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6612 39850 6652 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6612 39770 6652 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6612 39690 6652 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6612 39610 6652 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6612 39530 6652 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6612 39450 6652 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6532 39930 6572 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6532 39850 6572 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6532 39770 6572 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6532 39690 6572 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6532 39610 6572 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6532 39530 6572 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6532 39450 6572 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6452 39930 6492 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6452 39850 6492 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6452 39770 6492 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6452 39690 6492 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6452 39610 6492 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6452 39530 6492 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6452 39450 6492 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6372 39930 6412 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6372 39850 6412 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6372 39770 6412 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6372 39690 6412 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6372 39610 6412 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6372 39530 6412 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6372 39450 6412 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6292 39930 6332 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6292 39850 6332 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6292 39770 6332 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6292 39690 6332 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6292 39610 6332 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6292 39530 6332 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6292 39450 6332 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6212 39930 6252 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6212 39850 6252 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6212 39770 6252 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6212 39690 6252 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6212 39610 6252 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6212 39530 6252 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6212 39450 6252 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6132 39930 6172 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6132 39850 6172 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6132 39770 6172 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6132 39690 6172 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6132 39610 6172 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6132 39530 6172 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6132 39450 6172 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6052 39930 6092 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6052 39850 6092 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6052 39770 6092 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6052 39690 6092 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6052 39610 6092 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6052 39530 6092 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6052 39450 6092 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5972 39930 6012 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5972 39850 6012 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5972 39770 6012 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5972 39690 6012 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5972 39610 6012 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5972 39530 6012 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5972 39450 6012 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5892 39930 5932 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5892 39850 5932 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5892 39770 5932 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5892 39690 5932 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5892 39610 5932 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5892 39530 5932 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5892 39450 5932 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5812 39930 5852 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5812 39850 5852 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5812 39770 5852 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5812 39690 5852 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5812 39610 5852 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5812 39530 5852 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5812 39450 5852 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5732 39930 5772 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5732 39850 5772 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5732 39770 5772 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5732 39690 5772 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5732 39610 5772 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5732 39530 5772 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5732 39450 5772 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5652 39930 5692 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5652 39850 5692 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5652 39770 5692 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5652 39690 5692 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5652 39610 5692 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5652 39530 5692 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5652 39450 5692 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5572 39930 5612 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5572 39850 5612 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5572 39770 5612 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5572 39690 5612 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5572 39610 5612 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5572 39530 5612 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5572 39450 5612 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5492 39930 5532 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5492 39850 5532 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5492 39770 5532 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5492 39690 5532 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5492 39610 5532 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5492 39530 5532 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5492 39450 5532 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5412 39930 5452 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5412 39850 5452 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5412 39770 5452 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5412 39690 5452 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5412 39610 5452 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5412 39530 5452 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5412 39450 5452 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5319 39918 5383 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5319 39838 5383 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5319 39758 5383 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5319 39678 5383 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5319 39598 5383 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5319 39518 5383 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5319 39438 5383 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5238 39918 5302 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5238 39838 5302 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5238 39758 5302 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5238 39678 5302 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5238 39598 5302 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5238 39518 5302 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5238 39438 5302 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5157 39918 5221 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5157 39838 5221 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5157 39758 5221 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5157 39678 5221 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5157 39598 5221 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5157 39518 5221 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5157 39438 5221 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5076 39918 5140 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5076 39838 5140 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5076 39758 5140 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5076 39678 5140 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5076 39598 5140 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5076 39518 5140 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5076 39438 5140 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4995 39918 5059 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4995 39838 5059 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4995 39758 5059 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4995 39678 5059 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4995 39598 5059 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4995 39518 5059 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4995 39438 5059 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4914 39918 4978 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4914 39838 4978 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4914 39758 4978 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4914 39678 4978 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4914 39598 4978 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4914 39518 4978 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4914 39438 4978 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4833 39918 4897 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4833 39838 4897 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4833 39758 4897 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4833 39678 4897 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4833 39598 4897 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4833 39518 4897 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4833 39438 4897 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4821 6042 4861 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4821 5956 4861 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4821 5870 4861 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4821 5784 4861 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4821 5698 4861 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4821 5612 4861 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4821 5526 4861 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4821 5440 4861 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4821 5354 4861 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4821 5268 4861 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4821 5182 4861 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4752 39918 4816 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4752 39838 4816 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4752 39758 4816 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4752 39678 4816 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4752 39598 4816 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4752 39518 4816 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4752 39438 4816 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4740 6042 4780 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4740 5956 4780 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4740 5870 4780 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4740 5784 4780 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4740 5698 4780 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4740 5612 4780 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4740 5526 4780 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4740 5440 4780 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4740 5354 4780 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4740 5268 4780 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4740 5182 4780 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4671 39918 4735 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4671 39838 4735 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4671 39758 4735 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4671 39678 4735 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4671 39598 4735 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4671 39518 4735 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4671 39438 4735 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4659 6042 4699 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4659 5956 4699 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4659 5870 4699 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4659 5784 4699 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4659 5698 4699 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4659 5612 4699 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4659 5526 4699 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4659 5440 4699 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4659 5354 4699 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4659 5268 4699 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4659 5182 4699 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4590 39918 4654 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4590 39838 4654 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4590 39758 4654 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4590 39678 4654 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4590 39598 4654 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4590 39518 4654 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4590 39438 4654 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 6042 4618 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5956 4618 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5870 4618 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5784 4618 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5698 4618 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5612 4618 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5526 4618 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5440 4618 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5354 4618 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5268 4618 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5182 4618 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4509 39918 4573 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4509 39838 4573 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4509 39758 4573 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4509 39678 4573 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4509 39598 4573 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4509 39518 4573 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4509 39438 4573 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4497 6042 4537 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4497 5956 4537 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4497 5870 4537 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4497 5784 4537 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4497 5698 4537 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4497 5612 4537 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4497 5526 4537 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4497 5440 4537 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4497 5354 4537 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4497 5268 4537 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4497 5182 4537 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4428 39918 4492 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4428 39838 4492 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4428 39758 4492 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4428 39678 4492 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4428 39598 4492 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4428 39518 4492 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4428 39438 4492 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4416 6042 4456 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4416 5956 4456 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4416 5870 4456 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4416 5784 4456 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4416 5698 4456 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4416 5612 4456 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4416 5526 4456 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4416 5440 4456 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4416 5354 4456 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4416 5268 4456 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4416 5182 4456 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4347 39918 4411 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4347 39838 4411 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4347 39758 4411 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4347 39678 4411 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4347 39598 4411 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4347 39518 4411 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4347 39438 4411 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4335 6042 4375 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4335 5956 4375 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4335 5870 4375 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4335 5784 4375 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4335 5698 4375 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4335 5612 4375 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4335 5526 4375 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4335 5440 4375 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4335 5354 4375 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4335 5268 4375 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4335 5182 4375 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4266 39918 4330 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4266 39838 4330 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4266 39758 4330 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4266 39678 4330 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4266 39598 4330 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4266 39518 4330 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4266 39438 4330 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 6042 4294 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5956 4294 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5870 4294 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5784 4294 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5698 4294 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5612 4294 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5526 4294 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5440 4294 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5354 4294 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5268 4294 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5182 4294 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4185 39918 4249 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4185 39838 4249 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4185 39758 4249 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4185 39678 4249 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4185 39598 4249 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4185 39518 4249 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4185 39438 4249 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4173 6042 4213 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4173 5956 4213 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4173 5870 4213 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4173 5784 4213 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4173 5698 4213 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4173 5612 4213 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4173 5526 4213 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4173 5440 4213 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4173 5354 4213 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4173 5268 4213 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4173 5182 4213 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4104 39918 4168 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4104 39838 4168 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4104 39758 4168 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4104 39678 4168 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4104 39598 4168 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4104 39518 4168 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4104 39438 4168 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4092 6042 4132 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4092 5956 4132 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4092 5870 4132 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4092 5784 4132 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4092 5698 4132 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4092 5612 4132 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4092 5526 4132 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4092 5440 4132 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4092 5354 4132 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4092 5268 4132 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4092 5182 4132 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4023 39918 4087 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4023 39838 4087 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4023 39758 4087 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4023 39678 4087 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4023 39598 4087 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4023 39518 4087 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4023 39438 4087 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4011 6042 4051 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4011 5956 4051 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4011 5870 4051 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4011 5784 4051 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4011 5698 4051 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4011 5612 4051 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4011 5526 4051 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4011 5440 4051 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4011 5354 4051 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4011 5268 4051 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4011 5182 4051 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3942 39918 4006 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3942 39838 4006 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3942 39758 4006 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3942 39678 4006 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3942 39598 4006 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3942 39518 4006 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3942 39438 4006 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 6042 3970 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5956 3970 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5870 3970 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5784 3970 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5698 3970 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5612 3970 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5526 3970 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5440 3970 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5354 3970 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5268 3970 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5182 3970 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3861 39918 3925 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3861 39838 3925 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3861 39758 3925 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3861 39678 3925 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3861 39598 3925 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3861 39518 3925 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3861 39438 3925 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3849 6042 3889 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3849 5956 3889 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3849 5870 3889 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3849 5784 3889 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3849 5698 3889 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3849 5612 3889 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3849 5526 3889 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3849 5440 3889 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3849 5354 3889 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3849 5268 3889 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3849 5182 3889 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3780 39918 3844 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3780 39838 3844 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3780 39758 3844 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3780 39678 3844 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3780 39598 3844 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3780 39518 3844 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3780 39438 3844 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3768 6042 3808 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3768 5956 3808 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3768 5870 3808 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3768 5784 3808 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3768 5698 3808 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3768 5612 3808 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3768 5526 3808 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3768 5440 3808 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3768 5354 3808 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3768 5268 3808 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3768 5182 3808 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3699 39918 3763 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3699 39838 3763 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3699 39758 3763 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3699 39678 3763 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3699 39598 3763 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3699 39518 3763 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3699 39438 3763 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3687 6042 3727 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3687 5956 3727 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3687 5870 3727 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3687 5784 3727 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3687 5698 3727 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3687 5612 3727 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3687 5526 3727 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3687 5440 3727 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3687 5354 3727 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3687 5268 3727 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3687 5182 3727 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3618 39918 3682 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3618 39838 3682 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3618 39758 3682 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3618 39678 3682 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3618 39598 3682 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3618 39518 3682 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3618 39438 3682 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 6042 3646 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5956 3646 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5870 3646 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5784 3646 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5698 3646 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5612 3646 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5526 3646 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5440 3646 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5354 3646 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5268 3646 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5182 3646 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3537 39918 3601 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3537 39838 3601 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3537 39758 3601 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3537 39678 3601 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3537 39598 3601 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3537 39518 3601 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3537 39438 3601 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3525 6042 3565 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3525 5956 3565 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3525 5870 3565 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3525 5784 3565 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3525 5698 3565 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3525 5612 3565 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3525 5526 3565 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3525 5440 3565 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3525 5354 3565 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3525 5268 3565 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3525 5182 3565 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3456 39918 3520 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3456 39838 3520 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3456 39758 3520 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3456 39678 3520 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3456 39598 3520 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3456 39518 3520 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3456 39438 3520 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3444 6042 3484 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3444 5956 3484 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3444 5870 3484 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3444 5784 3484 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3444 5698 3484 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3444 5612 3484 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3444 5526 3484 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3444 5440 3484 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3444 5354 3484 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3444 5268 3484 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3444 5182 3484 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3375 39918 3439 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3375 39838 3439 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3375 39758 3439 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3375 39678 3439 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3375 39598 3439 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3375 39518 3439 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3375 39438 3439 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3363 6042 3403 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3363 5956 3403 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3363 5870 3403 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3363 5784 3403 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3363 5698 3403 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3363 5612 3403 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3363 5526 3403 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3363 5440 3403 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3363 5354 3403 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3363 5268 3403 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3363 5182 3403 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3294 39918 3358 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3294 39838 3358 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3294 39758 3358 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3294 39678 3358 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3294 39598 3358 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3294 39518 3358 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3294 39438 3358 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 6042 3322 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5956 3322 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5870 3322 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5784 3322 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5698 3322 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5612 3322 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5526 3322 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5440 3322 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5354 3322 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5268 3322 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5182 3322 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3213 39918 3277 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3213 39838 3277 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3213 39758 3277 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3213 39678 3277 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3213 39598 3277 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3213 39518 3277 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3213 39438 3277 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3201 6042 3241 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3201 5956 3241 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3201 5870 3241 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3201 5784 3241 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3201 5698 3241 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3201 5612 3241 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3201 5526 3241 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3201 5440 3241 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3201 5354 3241 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3201 5268 3241 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3201 5182 3241 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3132 39918 3196 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3132 39838 3196 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3132 39758 3196 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3132 39678 3196 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3132 39598 3196 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3132 39518 3196 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3132 39438 3196 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3120 6042 3160 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3120 5956 3160 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3120 5870 3160 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3120 5784 3160 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3120 5698 3160 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3120 5612 3160 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3120 5526 3160 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3120 5440 3160 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3120 5354 3160 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3120 5268 3160 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3120 5182 3160 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3051 39918 3115 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3051 39838 3115 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3051 39758 3115 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3051 39678 3115 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3051 39598 3115 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3051 39518 3115 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3051 39438 3115 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3039 6042 3079 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3039 5956 3079 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3039 5870 3079 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3039 5784 3079 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3039 5698 3079 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3039 5612 3079 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3039 5526 3079 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3039 5440 3079 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3039 5354 3079 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3039 5268 3079 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3039 5182 3079 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2970 39918 3034 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2970 39838 3034 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2970 39758 3034 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2970 39678 3034 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2970 39598 3034 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2970 39518 3034 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2970 39438 3034 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 6042 2998 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5956 2998 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5870 2998 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5784 2998 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5698 2998 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5612 2998 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5526 2998 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5440 2998 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5354 2998 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5268 2998 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5182 2998 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2889 39918 2953 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2889 39838 2953 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2889 39758 2953 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2889 39678 2953 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2889 39598 2953 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2889 39518 2953 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2889 39438 2953 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2877 6042 2917 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2877 5956 2917 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2877 5870 2917 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2877 5784 2917 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2877 5698 2917 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2877 5612 2917 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2877 5526 2917 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2877 5440 2917 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2877 5354 2917 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2877 5268 2917 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2877 5182 2917 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2808 39918 2872 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2808 39838 2872 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2808 39758 2872 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2808 39678 2872 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2808 39598 2872 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2808 39518 2872 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2808 39438 2872 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2796 6042 2836 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2796 5956 2836 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2796 5870 2836 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2796 5784 2836 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2796 5698 2836 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2796 5612 2836 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2796 5526 2836 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2796 5440 2836 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2796 5354 2836 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2796 5268 2836 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2796 5182 2836 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2753 39329 2817 39393 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2753 39247 2817 39311 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2727 39918 2791 39982 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2727 39838 2791 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2727 39758 2791 39822 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2727 39678 2791 39742 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2727 39598 2791 39662 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2727 39518 2791 39582 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2727 39438 2791 39502 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2715 6042 2755 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2715 5956 2755 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2715 5870 2755 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2715 5784 2755 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2715 5698 2755 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2715 5612 2755 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2715 5526 2755 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2715 5440 2755 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2715 5354 2755 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2715 5268 2755 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2715 5182 2755 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 6042 2674 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5956 2674 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5870 2674 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5784 2674 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5698 2674 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5612 2674 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5526 2674 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5440 2674 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5354 2674 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5268 2674 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5182 2674 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2605 39919 2669 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2605 39838 2669 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2605 39757 2669 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2605 39676 2669 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2605 39595 2669 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2605 39514 2669 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2605 39433 2669 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2605 39352 2669 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2605 39271 2669 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2605 39190 2669 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2605 39109 2669 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2605 39028 2669 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 125 35187 2669 39011 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 38879 2657 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 38799 2657 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 38719 2657 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 38639 2657 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 38559 2657 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 38479 2657 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 38399 2657 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 38319 2657 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 38239 2657 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 38159 2657 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 38079 2657 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 37999 2657 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 37919 2657 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 37839 2657 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 37759 2657 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 37679 2657 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 37599 2657 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 37519 2657 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 37439 2657 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 37359 2657 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 37279 2657 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 37199 2657 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 37119 2657 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 37039 2657 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 36959 2657 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 36879 2657 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 36799 2657 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 36719 2657 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 36639 2657 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 36559 2657 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 36479 2657 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 36399 2657 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 36319 2657 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 36239 2657 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 36159 2657 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 36079 2657 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 35999 2657 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 35919 2657 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 35839 2657 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 35759 2657 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 35679 2657 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 35599 2657 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 35519 2657 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 35439 2657 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 35359 2657 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 35279 2657 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 35199 2657 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2553 6042 2593 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2553 5956 2593 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2553 5870 2593 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2553 5784 2593 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2553 5698 2593 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2553 5612 2593 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2553 5526 2593 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2553 5440 2593 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2553 5354 2593 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2553 5268 2593 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2553 5182 2593 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2525 39919 2589 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2525 39838 2589 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2525 39757 2589 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2525 39676 2589 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2525 39595 2589 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2525 39514 2589 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2525 39433 2589 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2525 39352 2589 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2525 39271 2589 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2525 39190 2589 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2525 39109 2589 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2525 39028 2589 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 38959 2577 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 38879 2577 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 38799 2577 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 38719 2577 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 38639 2577 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 38559 2577 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 38479 2577 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 38399 2577 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 38319 2577 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 38239 2577 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 38159 2577 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 38079 2577 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 37999 2577 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 37919 2577 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 37839 2577 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 37759 2577 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 37679 2577 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 37599 2577 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 37519 2577 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 37439 2577 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 37359 2577 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 37279 2577 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 37199 2577 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 37119 2577 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 37039 2577 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 36959 2577 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 36879 2577 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 36799 2577 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 36719 2577 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 36639 2577 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 36559 2577 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 36479 2577 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 36399 2577 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 36319 2577 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 36239 2577 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 36159 2577 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 36079 2577 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 35999 2577 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 35919 2577 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 35839 2577 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 35759 2577 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 35679 2577 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 35599 2577 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 35519 2577 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 35439 2577 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 35359 2577 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 35279 2577 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 35199 2577 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2472 6042 2512 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2472 5956 2512 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2472 5870 2512 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2472 5784 2512 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2472 5698 2512 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2472 5612 2512 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2472 5526 2512 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2472 5440 2512 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2472 5354 2512 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2472 5268 2512 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2472 5182 2512 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2445 39919 2509 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2445 39838 2509 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2445 39757 2509 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2445 39676 2509 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2445 39595 2509 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2445 39514 2509 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2445 39433 2509 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2445 39352 2509 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2445 39271 2509 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2445 39190 2509 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2445 39109 2509 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2445 39028 2509 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 38959 2497 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 38879 2497 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 38799 2497 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 38719 2497 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 38639 2497 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 38559 2497 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 38479 2497 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 38399 2497 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 38319 2497 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 38239 2497 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 38159 2497 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 38079 2497 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 37999 2497 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 37919 2497 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 37839 2497 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 37759 2497 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 37679 2497 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 37599 2497 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 37519 2497 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 37439 2497 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 37359 2497 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 37279 2497 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 37199 2497 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 37119 2497 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 37039 2497 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 36959 2497 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 36879 2497 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 36799 2497 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 36719 2497 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 36639 2497 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 36559 2497 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 36479 2497 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 36399 2497 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 36319 2497 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 36239 2497 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 36159 2497 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 36079 2497 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 35999 2497 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 35919 2497 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 35839 2497 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 35759 2497 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 35679 2497 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 35599 2497 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 35519 2497 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 35439 2497 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 35359 2497 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 35279 2497 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 35199 2497 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2391 6042 2431 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2391 5956 2431 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2391 5870 2431 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2391 5784 2431 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2391 5698 2431 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2391 5612 2431 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2391 5526 2431 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2391 5440 2431 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2391 5354 2431 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2391 5268 2431 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2391 5182 2431 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2365 39919 2429 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2365 39838 2429 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2365 39757 2429 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2365 39676 2429 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2365 39595 2429 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2365 39514 2429 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2365 39433 2429 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2365 39352 2429 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2365 39271 2429 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2365 39190 2429 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2365 39109 2429 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2365 39028 2429 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 38959 2417 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 38879 2417 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 38799 2417 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 38719 2417 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 38639 2417 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 38559 2417 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 38479 2417 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 38399 2417 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 38319 2417 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 38239 2417 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 38159 2417 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 38079 2417 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 37999 2417 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 37919 2417 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 37839 2417 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 37759 2417 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 37679 2417 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 37599 2417 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 37519 2417 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 37439 2417 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 37359 2417 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 37279 2417 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 37199 2417 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 37119 2417 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 37039 2417 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 36959 2417 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 36879 2417 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 36799 2417 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 36719 2417 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 36639 2417 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 36559 2417 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 36479 2417 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 36399 2417 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 36319 2417 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 36239 2417 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 36159 2417 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 36079 2417 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 35999 2417 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 35919 2417 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 35839 2417 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 35759 2417 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 35679 2417 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 35599 2417 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 35519 2417 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 35439 2417 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 35359 2417 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 35279 2417 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 35199 2417 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 6042 2350 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5956 2350 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5870 2350 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5784 2350 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5698 2350 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5612 2350 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5526 2350 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5440 2350 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5354 2350 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5268 2350 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5182 2350 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2285 39919 2349 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2285 39838 2349 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2285 39757 2349 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2285 39676 2349 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2285 39595 2349 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2285 39514 2349 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2285 39433 2349 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2285 39352 2349 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2285 39271 2349 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2285 39190 2349 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2285 39109 2349 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2285 39028 2349 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 38959 2337 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 38879 2337 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 38799 2337 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 38719 2337 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 38639 2337 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 38559 2337 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 38479 2337 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 38399 2337 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 38319 2337 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 38239 2337 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 38159 2337 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 38079 2337 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 37999 2337 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 37919 2337 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 37839 2337 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 37759 2337 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 37679 2337 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 37599 2337 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 37519 2337 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 37439 2337 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 37359 2337 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 37279 2337 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 37199 2337 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 37119 2337 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 37039 2337 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 36959 2337 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 36879 2337 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 36799 2337 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 36719 2337 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 36639 2337 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 36559 2337 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 36479 2337 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 36399 2337 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 36319 2337 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 36239 2337 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 36159 2337 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 36079 2337 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 35999 2337 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 35919 2337 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 35839 2337 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 35759 2337 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 35679 2337 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 35599 2337 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 35519 2337 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 35439 2337 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 35359 2337 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 35279 2337 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 35199 2337 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2229 6042 2269 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2229 5956 2269 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2229 5870 2269 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2229 5784 2269 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2229 5698 2269 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2229 5612 2269 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2229 5526 2269 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2229 5440 2269 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2229 5354 2269 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2229 5268 2269 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2229 5182 2269 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2205 39919 2269 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2205 39838 2269 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2205 39757 2269 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2205 39676 2269 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2205 39595 2269 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2205 39514 2269 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2205 39433 2269 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2205 39352 2269 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2205 39271 2269 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2205 39190 2269 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2205 39109 2269 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2205 39028 2269 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 38959 2257 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 38879 2257 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 38799 2257 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 38719 2257 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 38639 2257 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 38559 2257 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 38479 2257 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 38399 2257 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 38319 2257 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 38239 2257 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 38159 2257 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 38079 2257 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 37999 2257 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 37919 2257 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 37839 2257 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 37759 2257 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 37679 2257 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 37599 2257 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 37519 2257 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 37439 2257 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 37359 2257 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 37279 2257 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 37199 2257 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 37119 2257 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 37039 2257 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 36959 2257 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 36879 2257 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 36799 2257 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 36719 2257 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 36639 2257 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 36559 2257 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 36479 2257 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 36399 2257 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 36319 2257 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 36239 2257 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 36159 2257 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 36079 2257 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 35999 2257 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 35919 2257 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 35839 2257 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 35759 2257 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 35679 2257 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 35599 2257 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 35519 2257 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 35439 2257 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 35359 2257 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 35279 2257 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 35199 2257 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2148 6042 2188 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2148 5956 2188 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2148 5870 2188 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2148 5784 2188 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2148 5698 2188 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2148 5612 2188 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2148 5526 2188 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2148 5440 2188 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2148 5354 2188 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2148 5268 2188 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2148 5182 2188 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2125 39919 2189 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2125 39838 2189 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2125 39757 2189 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2125 39676 2189 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2125 39595 2189 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2125 39514 2189 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2125 39433 2189 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2125 39352 2189 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2125 39271 2189 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2125 39190 2189 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2125 39109 2189 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2125 39028 2189 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 38959 2177 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 38879 2177 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 38799 2177 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 38719 2177 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 38639 2177 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 38559 2177 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 38479 2177 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 38399 2177 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 38319 2177 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 38239 2177 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 38159 2177 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 38079 2177 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 37999 2177 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 37919 2177 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 37839 2177 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 37759 2177 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 37679 2177 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 37599 2177 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 37519 2177 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 37439 2177 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 37359 2177 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 37279 2177 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 37199 2177 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 37119 2177 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 37039 2177 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 36959 2177 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 36879 2177 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 36799 2177 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 36719 2177 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 36639 2177 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 36559 2177 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 36479 2177 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 36399 2177 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 36319 2177 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 36239 2177 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 36159 2177 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 36079 2177 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 35999 2177 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 35919 2177 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 35839 2177 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 35759 2177 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 35679 2177 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 35599 2177 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 35519 2177 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 35439 2177 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 35359 2177 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 35279 2177 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 35199 2177 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2067 6042 2107 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2067 5956 2107 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2067 5870 2107 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2067 5784 2107 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2067 5698 2107 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2067 5612 2107 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2067 5526 2107 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2067 5440 2107 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2067 5354 2107 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2067 5268 2107 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2067 5182 2107 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2045 39919 2109 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2045 39838 2109 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2045 39757 2109 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2045 39676 2109 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2045 39595 2109 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2045 39514 2109 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2045 39433 2109 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2045 39352 2109 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2045 39271 2109 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2045 39190 2109 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2045 39109 2109 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2045 39028 2109 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 38959 2097 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 38879 2097 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 38799 2097 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 38719 2097 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 38639 2097 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 38559 2097 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 38479 2097 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 38399 2097 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 38319 2097 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 38239 2097 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 38159 2097 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 38079 2097 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 37999 2097 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 37919 2097 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 37839 2097 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 37759 2097 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 37679 2097 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 37599 2097 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 37519 2097 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 37439 2097 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 37359 2097 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 37279 2097 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 37199 2097 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 37119 2097 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 37039 2097 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 36959 2097 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 36879 2097 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 36799 2097 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 36719 2097 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 36639 2097 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 36559 2097 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 36479 2097 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 36399 2097 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 36319 2097 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 36239 2097 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 36159 2097 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 36079 2097 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 35999 2097 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 35919 2097 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 35839 2097 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 35759 2097 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 35679 2097 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 35599 2097 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 35519 2097 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 35439 2097 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 35359 2097 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 35279 2097 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 35199 2097 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 6042 2026 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5956 2026 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5870 2026 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5784 2026 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5698 2026 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5612 2026 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5526 2026 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5440 2026 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5354 2026 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5268 2026 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5182 2026 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1965 39919 2029 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1965 39838 2029 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1965 39757 2029 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1965 39676 2029 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1965 39595 2029 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1965 39514 2029 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1965 39433 2029 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1965 39352 2029 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1965 39271 2029 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1965 39190 2029 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1965 39109 2029 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1965 39028 2029 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 38959 2017 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 38879 2017 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 38799 2017 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 38719 2017 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 38639 2017 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 38559 2017 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 38479 2017 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 38399 2017 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 38319 2017 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 38239 2017 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 38159 2017 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 38079 2017 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 37999 2017 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 37919 2017 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 37839 2017 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 37759 2017 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 37679 2017 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 37599 2017 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 37519 2017 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 37439 2017 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 37359 2017 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 37279 2017 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 37199 2017 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 37119 2017 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 37039 2017 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 36959 2017 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 36879 2017 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 36799 2017 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 36719 2017 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 36639 2017 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 36559 2017 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 36479 2017 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 36399 2017 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 36319 2017 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 36239 2017 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 36159 2017 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 36079 2017 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 35999 2017 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 35919 2017 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 35839 2017 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 35759 2017 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 35679 2017 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 35599 2017 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 35519 2017 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 35439 2017 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 35359 2017 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 35279 2017 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 35199 2017 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1905 6042 1945 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1905 5956 1945 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1905 5870 1945 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1905 5784 1945 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1905 5698 1945 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1905 5612 1945 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1905 5526 1945 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1905 5440 1945 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1905 5354 1945 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1905 5268 1945 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1905 5182 1945 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1885 39919 1949 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1885 39838 1949 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1885 39757 1949 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1885 39676 1949 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1885 39595 1949 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1885 39514 1949 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1885 39433 1949 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1885 39352 1949 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1885 39271 1949 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1885 39190 1949 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1885 39109 1949 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1885 39028 1949 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 38959 1937 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 38879 1937 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 38799 1937 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 38719 1937 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 38639 1937 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 38559 1937 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 38479 1937 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 38399 1937 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 38319 1937 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 38239 1937 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 38159 1937 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 38079 1937 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 37999 1937 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 37919 1937 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 37839 1937 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 37759 1937 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 37679 1937 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 37599 1937 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 37519 1937 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 37439 1937 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 37359 1937 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 37279 1937 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 37199 1937 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 37119 1937 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 37039 1937 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 36959 1937 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 36879 1937 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 36799 1937 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 36719 1937 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 36639 1937 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 36559 1937 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 36479 1937 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 36399 1937 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 36319 1937 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 36239 1937 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 36159 1937 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 36079 1937 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 35999 1937 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 35919 1937 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 35839 1937 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 35759 1937 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 35679 1937 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 35599 1937 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 35519 1937 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 35439 1937 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 35359 1937 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 35279 1937 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 35199 1937 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1824 6042 1864 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1824 5956 1864 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1824 5870 1864 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1824 5784 1864 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1824 5698 1864 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1824 5612 1864 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1824 5526 1864 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1824 5440 1864 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1824 5354 1864 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1824 5268 1864 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1824 5182 1864 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1805 39919 1869 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1805 39838 1869 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1805 39757 1869 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1805 39676 1869 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1805 39595 1869 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1805 39514 1869 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1805 39433 1869 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1805 39352 1869 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1805 39271 1869 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1805 39190 1869 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1805 39109 1869 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1805 39028 1869 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 38959 1857 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 38879 1857 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 38799 1857 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 38719 1857 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 38639 1857 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 38559 1857 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 38479 1857 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 38399 1857 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 38319 1857 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 38239 1857 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 38159 1857 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 38079 1857 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 37999 1857 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 37919 1857 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 37839 1857 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 37759 1857 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 37679 1857 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 37599 1857 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 37519 1857 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 37439 1857 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 37359 1857 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 37279 1857 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 37199 1857 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 37119 1857 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 37039 1857 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 36959 1857 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 36879 1857 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 36799 1857 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 36719 1857 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 36639 1857 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 36559 1857 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 36479 1857 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 36399 1857 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 36319 1857 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 36239 1857 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 36159 1857 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 36079 1857 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 35999 1857 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 35919 1857 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 35839 1857 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 35759 1857 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 35679 1857 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 35599 1857 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 35519 1857 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 35439 1857 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 35359 1857 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 35279 1857 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 35199 1857 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1743 6042 1783 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1743 5956 1783 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1743 5870 1783 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1743 5784 1783 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1743 5698 1783 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1743 5612 1783 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1743 5526 1783 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1743 5440 1783 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1743 5354 1783 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1743 5268 1783 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1743 5182 1783 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1725 39919 1789 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1725 39838 1789 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1725 39757 1789 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1725 39676 1789 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1725 39595 1789 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1725 39514 1789 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1725 39433 1789 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1725 39352 1789 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1725 39271 1789 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1725 39190 1789 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1725 39109 1789 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1725 39028 1789 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 38959 1777 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 38879 1777 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 38799 1777 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 38719 1777 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 38639 1777 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 38559 1777 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 38479 1777 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 38399 1777 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 38319 1777 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 38239 1777 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 38159 1777 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 38079 1777 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 37999 1777 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 37919 1777 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 37839 1777 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 37759 1777 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 37679 1777 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 37599 1777 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 37519 1777 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 37439 1777 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 37359 1777 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 37279 1777 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 37199 1777 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 37119 1777 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 37039 1777 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 36959 1777 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 36879 1777 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 36799 1777 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 36719 1777 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 36639 1777 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 36559 1777 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 36479 1777 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 36399 1777 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 36319 1777 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 36239 1777 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 36159 1777 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 36079 1777 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 35999 1777 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 35919 1777 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 35839 1777 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 35759 1777 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 35679 1777 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 35599 1777 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 35519 1777 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 35439 1777 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 35359 1777 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 35279 1777 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 35199 1777 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 6042 1702 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5956 1702 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5870 1702 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5784 1702 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5698 1702 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5612 1702 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5526 1702 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5440 1702 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5354 1702 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5268 1702 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5182 1702 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1645 39919 1709 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1645 39838 1709 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1645 39757 1709 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1645 39676 1709 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1645 39595 1709 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1645 39514 1709 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1645 39433 1709 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1645 39352 1709 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1645 39271 1709 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1645 39190 1709 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1645 39109 1709 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1645 39028 1709 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 38959 1697 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 38879 1697 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 38799 1697 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 38719 1697 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 38639 1697 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 38559 1697 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 38479 1697 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 38399 1697 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 38319 1697 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 38239 1697 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 38159 1697 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 38079 1697 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 37999 1697 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 37919 1697 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 37839 1697 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 37759 1697 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 37679 1697 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 37599 1697 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 37519 1697 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 37439 1697 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 37359 1697 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 37279 1697 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 37199 1697 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 37119 1697 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 37039 1697 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 36959 1697 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 36879 1697 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 36799 1697 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 36719 1697 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 36639 1697 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 36559 1697 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 36479 1697 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 36399 1697 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 36319 1697 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 36239 1697 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 36159 1697 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 36079 1697 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 35999 1697 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 35919 1697 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 35839 1697 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 35759 1697 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 35679 1697 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 35599 1697 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 35519 1697 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 35439 1697 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 35359 1697 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 35279 1697 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 35199 1697 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1581 6042 1621 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1581 5956 1621 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1581 5870 1621 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1581 5784 1621 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1581 5698 1621 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1581 5612 1621 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1581 5526 1621 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1581 5440 1621 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1581 5354 1621 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1581 5268 1621 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1581 5182 1621 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1565 39919 1629 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1565 39838 1629 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1565 39757 1629 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1565 39676 1629 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1565 39595 1629 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1565 39514 1629 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1565 39433 1629 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1565 39352 1629 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1565 39271 1629 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1565 39190 1629 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1565 39109 1629 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1565 39028 1629 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 38959 1617 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 38879 1617 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 38799 1617 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 38719 1617 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 38639 1617 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 38559 1617 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 38479 1617 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 38399 1617 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 38319 1617 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 38239 1617 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 38159 1617 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 38079 1617 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 37999 1617 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 37919 1617 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 37839 1617 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 37759 1617 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 37679 1617 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 37599 1617 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 37519 1617 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 37439 1617 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 37359 1617 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 37279 1617 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 37199 1617 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 37119 1617 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 37039 1617 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 36959 1617 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 36879 1617 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 36799 1617 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 36719 1617 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 36639 1617 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 36559 1617 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 36479 1617 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 36399 1617 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 36319 1617 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 36239 1617 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 36159 1617 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 36079 1617 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 35999 1617 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 35919 1617 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 35839 1617 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 35759 1617 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 35679 1617 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 35599 1617 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 35519 1617 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 35439 1617 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 35359 1617 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 35279 1617 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 35199 1617 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1500 6042 1540 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1500 5956 1540 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1500 5870 1540 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1500 5784 1540 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1500 5698 1540 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1500 5612 1540 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1500 5526 1540 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1500 5440 1540 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1500 5354 1540 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1500 5268 1540 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1500 5182 1540 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1485 39919 1549 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1485 39838 1549 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1485 39757 1549 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1485 39676 1549 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1485 39595 1549 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1485 39514 1549 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1485 39433 1549 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1485 39352 1549 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1485 39271 1549 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1485 39190 1549 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1485 39109 1549 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1485 39028 1549 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 38959 1537 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 38879 1537 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 38799 1537 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 38719 1537 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 38639 1537 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 38559 1537 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 38479 1537 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 38399 1537 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 38319 1537 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 38239 1537 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 38159 1537 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 38079 1537 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 37999 1537 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 37919 1537 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 37839 1537 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 37759 1537 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 37679 1537 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 37599 1537 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 37519 1537 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 37439 1537 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 37359 1537 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 37279 1537 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 37199 1537 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 37119 1537 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 37039 1537 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 36959 1537 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 36879 1537 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 36799 1537 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 36719 1537 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 36639 1537 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 36559 1537 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 36479 1537 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 36399 1537 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 36319 1537 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 36239 1537 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 36159 1537 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 36079 1537 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 35999 1537 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 35919 1537 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 35839 1537 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 35759 1537 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 35679 1537 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 35599 1537 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 35519 1537 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 35439 1537 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 35359 1537 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 35279 1537 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 35199 1537 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1419 6042 1459 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1419 5956 1459 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1419 5870 1459 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1419 5784 1459 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1419 5698 1459 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1419 5612 1459 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1419 5526 1459 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1419 5440 1459 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1419 5354 1459 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1419 5268 1459 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1419 5182 1459 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1405 39919 1469 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1405 39838 1469 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1405 39757 1469 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1405 39676 1469 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1405 39595 1469 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1405 39514 1469 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1405 39433 1469 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1405 39352 1469 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1405 39271 1469 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1405 39190 1469 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1405 39109 1469 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1405 39028 1469 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 38959 1457 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 38879 1457 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 38799 1457 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 38719 1457 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 38639 1457 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 38559 1457 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 38479 1457 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 38399 1457 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 38319 1457 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 38239 1457 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 38159 1457 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 38079 1457 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 37999 1457 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 37919 1457 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 37839 1457 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 37759 1457 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 37679 1457 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 37599 1457 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 37519 1457 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 37439 1457 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 37359 1457 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 37279 1457 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 37199 1457 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 37119 1457 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 37039 1457 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 36959 1457 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 36879 1457 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 36799 1457 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 36719 1457 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 36639 1457 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 36559 1457 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 36479 1457 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 36399 1457 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 36319 1457 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 36239 1457 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 36159 1457 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 36079 1457 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 35999 1457 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 35919 1457 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 35839 1457 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 35759 1457 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 35679 1457 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 35599 1457 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 35519 1457 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 35439 1457 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 35359 1457 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 35279 1457 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 35199 1457 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 6042 1378 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5956 1378 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5870 1378 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5784 1378 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5698 1378 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5612 1378 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5526 1378 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5440 1378 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5354 1378 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5268 1378 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5182 1378 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1325 39919 1389 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1325 39838 1389 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1325 39757 1389 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1325 39676 1389 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1325 39595 1389 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1325 39514 1389 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1325 39433 1389 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1325 39352 1389 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1325 39271 1389 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1325 39190 1389 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1325 39109 1389 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1325 39028 1389 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 38959 1377 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 38879 1377 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 38799 1377 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 38719 1377 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 38639 1377 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 38559 1377 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 38479 1377 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 38399 1377 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 38319 1377 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 38239 1377 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 38159 1377 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 38079 1377 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 37999 1377 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 37919 1377 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 37839 1377 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 37759 1377 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 37679 1377 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 37599 1377 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 37519 1377 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 37439 1377 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 37359 1377 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 37279 1377 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 37199 1377 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 37119 1377 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 37039 1377 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 36959 1377 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 36879 1377 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 36799 1377 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 36719 1377 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 36639 1377 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 36559 1377 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 36479 1377 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 36399 1377 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 36319 1377 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 36239 1377 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 36159 1377 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 36079 1377 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 35999 1377 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 35919 1377 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 35839 1377 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 35759 1377 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 35679 1377 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 35599 1377 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 35519 1377 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 35439 1377 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 35359 1377 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 35279 1377 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 35199 1377 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1245 39919 1309 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1245 39838 1309 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1245 39757 1309 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1245 39676 1309 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1245 39595 1309 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1245 39514 1309 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1245 39433 1309 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1245 39352 1309 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1245 39271 1309 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1245 39190 1309 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1245 39109 1309 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1245 39028 1309 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 38959 1297 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 38879 1297 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 38799 1297 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 38719 1297 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 38639 1297 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 38559 1297 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 38479 1297 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 38399 1297 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 38319 1297 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 38239 1297 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 38159 1297 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 38079 1297 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 37999 1297 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 37919 1297 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 37839 1297 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 37759 1297 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 37679 1297 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 37599 1297 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 37519 1297 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 37439 1297 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 37359 1297 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 37279 1297 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 37199 1297 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 37119 1297 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 37039 1297 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 36959 1297 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 36879 1297 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 36799 1297 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 36719 1297 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 36639 1297 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 36559 1297 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 36479 1297 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 36399 1297 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 36319 1297 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 36239 1297 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 36159 1297 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 36079 1297 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 35999 1297 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 35919 1297 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 35839 1297 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 35759 1297 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 35679 1297 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 35599 1297 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 35519 1297 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 35439 1297 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 35359 1297 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 35279 1297 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 35199 1297 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 6042 1297 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 5956 1297 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 5870 1297 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 5784 1297 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 5698 1297 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 5612 1297 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 5526 1297 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 5440 1297 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 5354 1297 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 5268 1297 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 5182 1297 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1165 39919 1229 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1165 39838 1229 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1165 39757 1229 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1165 39676 1229 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1165 39595 1229 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1165 39514 1229 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1165 39433 1229 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1165 39352 1229 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1165 39271 1229 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1165 39190 1229 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1165 39109 1229 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1165 39028 1229 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 38959 1217 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 38879 1217 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 38799 1217 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 38719 1217 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 38639 1217 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 38559 1217 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 38479 1217 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 38399 1217 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 38319 1217 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 38239 1217 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 38159 1217 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 38079 1217 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 37999 1217 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 37919 1217 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 37839 1217 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 37759 1217 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 37679 1217 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 37599 1217 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 37519 1217 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 37439 1217 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 37359 1217 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 37279 1217 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 37199 1217 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 37119 1217 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 37039 1217 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 36959 1217 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 36879 1217 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 36799 1217 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 36719 1217 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 36639 1217 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 36559 1217 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 36479 1217 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 36399 1217 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 36319 1217 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 36239 1217 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 36159 1217 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 36079 1217 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 35999 1217 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 35919 1217 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 35839 1217 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 35759 1217 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 35679 1217 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 35599 1217 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 35519 1217 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 35439 1217 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 35359 1217 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 35279 1217 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 35199 1217 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1176 6042 1216 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1176 5956 1216 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1176 5870 1216 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1176 5784 1216 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1176 5698 1216 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1176 5612 1216 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1176 5526 1216 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1176 5440 1216 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1176 5354 1216 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1176 5268 1216 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1176 5182 1216 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1085 39919 1149 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1085 39838 1149 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1085 39757 1149 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1085 39676 1149 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1085 39595 1149 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1085 39514 1149 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1085 39433 1149 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1085 39352 1149 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1085 39271 1149 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1085 39190 1149 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1085 39109 1149 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1085 39028 1149 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 38959 1137 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 38879 1137 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 38799 1137 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 38719 1137 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 38639 1137 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 38559 1137 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 38479 1137 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 38399 1137 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 38319 1137 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 38239 1137 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 38159 1137 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 38079 1137 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 37999 1137 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 37919 1137 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 37839 1137 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 37759 1137 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 37679 1137 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 37599 1137 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 37519 1137 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 37439 1137 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 37359 1137 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 37279 1137 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 37199 1137 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 37119 1137 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 37039 1137 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 36959 1137 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 36879 1137 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 36799 1137 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 36719 1137 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 36639 1137 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 36559 1137 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 36479 1137 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 36399 1137 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 36319 1137 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 36239 1137 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 36159 1137 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 36079 1137 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 35999 1137 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 35919 1137 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 35839 1137 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 35759 1137 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 35679 1137 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 35599 1137 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 35519 1137 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 35439 1137 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 35359 1137 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 35279 1137 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 35199 1137 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1095 6042 1135 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1095 5956 1135 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1095 5870 1135 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1095 5784 1135 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1095 5698 1135 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1095 5612 1135 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1095 5526 1135 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1095 5440 1135 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1095 5354 1135 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1095 5268 1135 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1095 5182 1135 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1005 39919 1069 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1005 39838 1069 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1005 39757 1069 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1005 39676 1069 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1005 39595 1069 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1005 39514 1069 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1005 39433 1069 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1005 39352 1069 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1005 39271 1069 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1005 39190 1069 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1005 39109 1069 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1005 39028 1069 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 38959 1057 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 38879 1057 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 38799 1057 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 38719 1057 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 38639 1057 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 38559 1057 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 38479 1057 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 38399 1057 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 38319 1057 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 38239 1057 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 38159 1057 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 38079 1057 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 37999 1057 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 37919 1057 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 37839 1057 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 37759 1057 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 37679 1057 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 37599 1057 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 37519 1057 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 37439 1057 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 37359 1057 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 37279 1057 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 37199 1057 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 37119 1057 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 37039 1057 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 36959 1057 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 36879 1057 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 36799 1057 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 36719 1057 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 36639 1057 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 36559 1057 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 36479 1057 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 36399 1057 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 36319 1057 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 36239 1057 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 36159 1057 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 36079 1057 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 35999 1057 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 35919 1057 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 35839 1057 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 35759 1057 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 35679 1057 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 35599 1057 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 35519 1057 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 35439 1057 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 35359 1057 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 35279 1057 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 35199 1057 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 6042 1054 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5956 1054 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5870 1054 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5784 1054 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5698 1054 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5612 1054 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5526 1054 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5440 1054 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5354 1054 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5268 1054 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5182 1054 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 925 39919 989 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 925 39838 989 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 925 39757 989 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 925 39676 989 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 925 39595 989 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 925 39514 989 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 925 39433 989 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 925 39352 989 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 925 39271 989 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 925 39190 989 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 925 39109 989 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 925 39028 989 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 38959 977 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 38879 977 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 38799 977 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 38719 977 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 38639 977 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 38559 977 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 38479 977 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 38399 977 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 38319 977 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 38239 977 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 38159 977 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 38079 977 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 37999 977 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 37919 977 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 37839 977 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 37759 977 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 37679 977 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 37599 977 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 37519 977 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 37439 977 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 37359 977 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 37279 977 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 37199 977 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 37119 977 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 37039 977 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 36959 977 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 36879 977 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 36799 977 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 36719 977 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 36639 977 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 36559 977 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 36479 977 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 36399 977 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 36319 977 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 36239 977 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 36159 977 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 36079 977 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 35999 977 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 35919 977 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 35839 977 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 35759 977 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 35679 977 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 35599 977 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 35519 977 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 35439 977 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 35359 977 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 35279 977 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 35199 977 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 933 6042 973 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 933 5956 973 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 933 5870 973 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 933 5784 973 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 933 5698 973 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 933 5612 973 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 933 5526 973 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 933 5440 973 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 933 5354 973 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 933 5268 973 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 933 5182 973 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 845 39919 909 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 845 39838 909 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 845 39757 909 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 845 39676 909 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 845 39595 909 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 845 39514 909 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 845 39433 909 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 845 39352 909 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 845 39271 909 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 845 39190 909 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 845 39109 909 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 845 39028 909 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 38959 897 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 38879 897 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 38799 897 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 38719 897 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 38639 897 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 38559 897 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 38479 897 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 38399 897 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 38319 897 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 38239 897 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 38159 897 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 38079 897 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 37999 897 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 37919 897 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 37839 897 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 37759 897 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 37679 897 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 37599 897 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 37519 897 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 37439 897 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 37359 897 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 37279 897 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 37199 897 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 37119 897 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 37039 897 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 36959 897 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 36879 897 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 36799 897 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 36719 897 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 36639 897 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 36559 897 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 36479 897 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 36399 897 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 36319 897 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 36239 897 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 36159 897 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 36079 897 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 35999 897 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 35919 897 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 35839 897 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 35759 897 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 35679 897 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 35599 897 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 35519 897 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 35439 897 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 35359 897 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 35279 897 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 35199 897 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 852 6042 892 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 852 5956 892 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 852 5870 892 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 852 5784 892 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 852 5698 892 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 852 5612 892 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 852 5526 892 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 852 5440 892 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 852 5354 892 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 852 5268 892 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 852 5182 892 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 765 39919 829 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 765 39838 829 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 765 39757 829 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 765 39676 829 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 765 39595 829 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 765 39514 829 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 765 39433 829 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 765 39352 829 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 765 39271 829 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 765 39190 829 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 765 39109 829 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 765 39028 829 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 38959 817 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 38879 817 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 38799 817 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 38719 817 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 38639 817 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 38559 817 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 38479 817 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 38399 817 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 38319 817 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 38239 817 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 38159 817 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 38079 817 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 37999 817 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 37919 817 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 37839 817 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 37759 817 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 37679 817 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 37599 817 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 37519 817 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 37439 817 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 37359 817 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 37279 817 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 37199 817 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 37119 817 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 37039 817 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 36959 817 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 36879 817 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 36799 817 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 36719 817 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 36639 817 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 36559 817 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 36479 817 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 36399 817 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 36319 817 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 36239 817 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 36159 817 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 36079 817 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 35999 817 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 35919 817 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 35839 817 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 35759 817 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 35679 817 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 35599 817 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 35519 817 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 35439 817 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 35359 817 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 35279 817 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 35199 817 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 771 6042 811 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 771 5956 811 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 771 5870 811 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 771 5784 811 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 771 5698 811 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 771 5612 811 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 771 5526 811 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 771 5440 811 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 771 5354 811 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 771 5268 811 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 771 5182 811 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 685 39919 749 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 685 39838 749 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 685 39757 749 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 685 39676 749 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 685 39595 749 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 685 39514 749 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 685 39433 749 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 685 39352 749 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 685 39271 749 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 685 39190 749 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 685 39109 749 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 685 39028 749 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 38959 737 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 38879 737 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 38799 737 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 38719 737 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 38639 737 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 38559 737 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 38479 737 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 38399 737 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 38319 737 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 38239 737 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 38159 737 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 38079 737 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 37999 737 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 37919 737 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 37839 737 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 37759 737 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 37679 737 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 37599 737 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 37519 737 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 37439 737 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 37359 737 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 37279 737 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 37199 737 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 37119 737 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 37039 737 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 36959 737 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 36879 737 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 36799 737 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 36719 737 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 36639 737 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 36559 737 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 36479 737 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 36399 737 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 36319 737 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 36239 737 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 36159 737 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 36079 737 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 35999 737 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 35919 737 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 35839 737 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 35759 737 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 35679 737 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 35599 737 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 35519 737 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 35439 737 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 35359 737 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 35279 737 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 35199 737 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 6042 730 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5956 730 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5870 730 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5784 730 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5698 730 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5612 730 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5526 730 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5440 730 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5354 730 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5268 730 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5182 730 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 605 39919 669 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 605 39838 669 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 605 39757 669 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 605 39676 669 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 605 39595 669 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 605 39514 669 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 605 39433 669 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 605 39352 669 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 605 39271 669 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 605 39190 669 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 605 39109 669 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 605 39028 669 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 38959 657 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 38879 657 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 38799 657 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 38719 657 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 38639 657 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 38559 657 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 38479 657 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 38399 657 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 38319 657 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 38239 657 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 38159 657 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 38079 657 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 37999 657 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 37919 657 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 37839 657 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 37759 657 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 37679 657 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 37599 657 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 37519 657 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 37439 657 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 37359 657 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 37279 657 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 37199 657 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 37119 657 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 37039 657 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 36959 657 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 36879 657 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 36799 657 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 36719 657 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 36639 657 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 36559 657 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 36479 657 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 36399 657 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 36319 657 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 36239 657 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 36159 657 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 36079 657 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 35999 657 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 35919 657 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 35839 657 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 35759 657 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 35679 657 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 35599 657 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 35519 657 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 35439 657 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 35359 657 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 35279 657 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 35199 657 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 609 6042 649 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 609 5956 649 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 609 5870 649 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 609 5784 649 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 609 5698 649 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 609 5612 649 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 609 5526 649 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 609 5440 649 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 609 5354 649 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 609 5268 649 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 609 5182 649 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 525 39919 589 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 525 39838 589 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 525 39757 589 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 525 39676 589 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 525 39595 589 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 525 39514 589 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 525 39433 589 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 525 39352 589 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 525 39271 589 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 525 39190 589 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 525 39109 589 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 525 39028 589 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 38959 577 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 38879 577 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 38799 577 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 38719 577 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 38639 577 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 38559 577 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 38479 577 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 38399 577 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 38319 577 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 38239 577 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 38159 577 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 38079 577 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 37999 577 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 37919 577 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 37839 577 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 37759 577 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 37679 577 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 37599 577 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 37519 577 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 37439 577 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 37359 577 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 37279 577 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 37199 577 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 37119 577 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 37039 577 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 36959 577 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 36879 577 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 36799 577 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 36719 577 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 36639 577 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 36559 577 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 36479 577 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 36399 577 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 36319 577 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 36239 577 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 36159 577 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 36079 577 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 35999 577 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 35919 577 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 35839 577 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 35759 577 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 35679 577 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 35599 577 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 35519 577 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 35439 577 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 35359 577 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 35279 577 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 35199 577 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 527 6042 567 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 527 5956 567 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 527 5870 567 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 527 5784 567 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 527 5698 567 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 527 5612 567 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 527 5526 567 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 527 5440 567 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 527 5354 567 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 527 5268 567 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 527 5182 567 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 39919 509 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 39838 509 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 39757 509 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 39676 509 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 39595 509 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 39514 509 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 39433 509 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 39352 509 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 39271 509 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 39190 509 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 39109 509 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 39028 509 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 38959 497 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 38879 497 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 38799 497 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 38719 497 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 38639 497 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 38559 497 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 38479 497 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 38399 497 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 38319 497 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 38239 497 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 38159 497 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 38079 497 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 37999 497 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 37919 497 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 37839 497 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 37759 497 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 37679 497 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 37599 497 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 37519 497 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 37439 497 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 37359 497 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 37279 497 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 37199 497 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 37119 497 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 37039 497 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 36959 497 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 36879 497 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 36799 497 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 36719 497 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 36639 497 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 36559 497 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 36479 497 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 36399 497 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 36319 497 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 36239 497 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 36159 497 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 36079 497 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 35999 497 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 35919 497 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 35839 497 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 35759 497 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 35679 497 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 35599 497 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 35519 497 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 35439 497 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 35359 497 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 35279 497 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 35199 497 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 6042 485 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 5956 485 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 5870 485 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 5784 485 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 5698 485 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 5612 485 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 5526 485 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 5440 485 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 5354 485 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 5268 485 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 5182 485 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 365 39919 429 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 365 39838 429 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 365 39757 429 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 365 39676 429 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 365 39595 429 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 365 39514 429 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 365 39433 429 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 365 39352 429 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 365 39271 429 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 365 39190 429 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 365 39109 429 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 365 39028 429 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 38959 417 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 38879 417 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 38799 417 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 38719 417 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 38639 417 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 38559 417 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 38479 417 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 38399 417 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 38319 417 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 38239 417 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 38159 417 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 38079 417 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 37999 417 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 37919 417 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 37839 417 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 37759 417 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 37679 417 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 37599 417 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 37519 417 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 37439 417 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 37359 417 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 37279 417 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 37199 417 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 37119 417 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 37039 417 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 36959 417 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 36879 417 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 36799 417 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 36719 417 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 36639 417 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 36559 417 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 36479 417 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 36399 417 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 36319 417 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 36239 417 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 36159 417 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 36079 417 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 35999 417 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 35919 417 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 35839 417 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 35759 417 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 35679 417 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 35599 417 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 35519 417 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 35439 417 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 35359 417 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 35279 417 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 35199 417 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 6042 403 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5956 403 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5870 403 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5784 403 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5698 403 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5612 403 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5526 403 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5440 403 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5354 403 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5268 403 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5182 403 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 285 39919 349 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 285 39838 349 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 285 39757 349 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 285 39676 349 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 285 39595 349 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 285 39514 349 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 285 39433 349 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 285 39352 349 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 285 39271 349 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 285 39190 349 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 285 39109 349 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 285 39028 349 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 38959 337 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 38879 337 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 38799 337 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 38719 337 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 38639 337 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 38559 337 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 38479 337 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 38399 337 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 38319 337 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 38239 337 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 38159 337 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 38079 337 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 37999 337 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 37919 337 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 37839 337 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 37759 337 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 37679 337 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 37599 337 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 37519 337 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 37439 337 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 37359 337 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 37279 337 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 37199 337 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 37119 337 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 37039 337 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 36959 337 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 36879 337 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 36799 337 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 36719 337 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 36639 337 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 36559 337 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 36479 337 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 36399 337 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 36319 337 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 36239 337 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 36159 337 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 36079 337 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 35999 337 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 35919 337 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 35839 337 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 35759 337 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 35679 337 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 35599 337 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 35519 337 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 35439 337 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 35359 337 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 35279 337 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 35199 337 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 281 6042 321 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 281 5956 321 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 281 5870 321 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 281 5784 321 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 281 5698 321 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 281 5612 321 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 281 5526 321 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 281 5440 321 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 281 5354 321 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 281 5268 321 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 281 5182 321 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 205 39919 269 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 205 39838 269 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 205 39757 269 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 205 39676 269 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 205 39595 269 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 205 39514 269 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 205 39433 269 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 205 39352 269 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 205 39271 269 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 205 39190 269 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 205 39109 269 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 205 39028 269 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 38959 257 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 38879 257 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 38799 257 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 38719 257 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 38639 257 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 38559 257 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 38479 257 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 38399 257 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 38319 257 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 38239 257 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 38159 257 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 38079 257 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 37999 257 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 37919 257 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 37839 257 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 37759 257 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 37679 257 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 37599 257 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 37519 257 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 37439 257 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 37359 257 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 37279 257 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 37199 257 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 37119 257 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 37039 257 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 36959 257 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 36879 257 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 36799 257 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 36719 257 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 36639 257 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 36559 257 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 36479 257 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 36399 257 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 36319 257 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 36239 257 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 36159 257 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 36079 257 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 35999 257 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 35919 257 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 35839 257 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 35759 257 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 35679 257 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 35599 257 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 35519 257 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 35439 257 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 35359 257 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 35279 257 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 35199 257 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 6042 239 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5956 239 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5870 239 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5784 239 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5698 239 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5612 239 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5526 239 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5440 239 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5354 239 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5268 239 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5182 239 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 125 39919 189 39983 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 125 39838 189 39902 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 125 39757 189 39821 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 125 39676 189 39740 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 125 39595 189 39659 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 125 39514 189 39578 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 125 39433 189 39497 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 125 39352 189 39416 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 125 39271 189 39335 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 125 39190 189 39254 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 125 39109 189 39173 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 125 39028 189 39092 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 38959 177 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 38879 177 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 38799 177 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 38719 177 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 38639 177 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 38559 177 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 38479 177 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 38399 177 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 38319 177 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 38239 177 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 38159 177 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 38079 177 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 37999 177 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 37919 177 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 37839 177 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 37759 177 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 37679 177 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 37599 177 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 37519 177 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 37439 177 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 37359 177 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 37279 177 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 37199 177 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 37119 177 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 37039 177 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 36959 177 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 36879 177 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 36799 177 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 36719 177 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 36639 177 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 36559 177 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 36479 177 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 36399 177 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 36319 177 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 36239 177 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 36159 177 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 36079 177 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 35999 177 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 35919 177 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 35839 177 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 35759 177 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 35679 177 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 35599 177 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 35519 177 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 35439 177 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 35359 177 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 35279 177 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 35199 177 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 6042 157 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5956 157 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5870 157 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5784 157 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5698 157 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5612 157 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5526 157 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5440 157 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5354 157 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5268 157 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5182 157 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10078 5168 14858 6096 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 0 39984 254 40000 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 0 35186 2695 39984 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 0 35157 254 35186 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 0 5167 4874 6097 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2719 39246 2851 39394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 2726 39434 12265 39986 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 10083 5167 15000 6097 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12136 39246 12268 39394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14746 39984 15000 40000 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 14746 35157 15000 35186 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal4 s 12301 35186 15000 39984 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 0 35157 254 40000 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 0 5187 254 6077 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 14746 35157 15000 40000 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 14746 5187 15000 6077 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 6042 14840 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5956 14840 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5870 14840 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5784 14840 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5698 14840 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5612 14840 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5526 14840 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5440 14840 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5354 14840 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5268 14840 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14800 5182 14840 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 39931 14838 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 39850 14838 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 39769 14838 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 39688 14838 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 39607 14838 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 39526 14838 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 39445 14838 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 39364 14838 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 39283 14838 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 39202 14838 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 39121 14838 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 39040 14838 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 38959 14838 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 38879 14838 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 38799 14838 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 38719 14838 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 38639 14838 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 38559 14838 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 38479 14838 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 38399 14838 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 38319 14838 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 38239 14838 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 38159 14838 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 38079 14838 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 37999 14838 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 37919 14838 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 37839 14838 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 37759 14838 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 37679 14838 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 37599 14838 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 37519 14838 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 37439 14838 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 37359 14838 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 37279 14838 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 37199 14838 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 37119 14838 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 37039 14838 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 36959 14838 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 36879 14838 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 36799 14838 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 36719 14838 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 36639 14838 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 36559 14838 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 36479 14838 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 36399 14838 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 36319 14838 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 36239 14838 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 36159 14838 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 36079 14838 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 35999 14838 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 35919 14838 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 35839 14838 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 35759 14838 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 35679 14838 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 35599 14838 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 35519 14838 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 35439 14838 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 35359 14838 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 35279 14838 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14798 35199 14838 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 6042 14759 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5956 14759 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5870 14759 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5784 14759 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5698 14759 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5612 14759 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5526 14759 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5440 14759 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5354 14759 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5268 14759 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14719 5182 14759 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 39931 14758 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 39850 14758 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 39769 14758 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 39688 14758 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 39607 14758 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 39526 14758 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 39445 14758 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 39364 14758 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 39283 14758 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 39202 14758 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 39121 14758 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 39040 14758 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 38959 14758 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 38879 14758 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 38799 14758 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 38719 14758 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 38639 14758 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 38559 14758 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 38479 14758 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 38399 14758 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 38319 14758 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 38239 14758 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 38159 14758 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 38079 14758 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 37999 14758 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 37919 14758 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 37839 14758 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 37759 14758 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 37679 14758 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 37599 14758 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 37519 14758 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 37439 14758 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 37359 14758 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 37279 14758 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 37199 14758 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 37119 14758 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 37039 14758 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 36959 14758 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 36879 14758 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 36799 14758 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 36719 14758 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 36639 14758 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 36559 14758 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 36479 14758 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 36399 14758 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 36319 14758 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 36239 14758 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 36159 14758 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 36079 14758 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 35999 14758 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 35919 14758 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 35839 14758 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 35759 14758 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 35679 14758 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 35599 14758 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 35519 14758 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 35439 14758 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 35359 14758 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 35279 14758 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14718 35199 14758 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 39931 14678 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 39850 14678 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 39769 14678 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 39688 14678 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 39607 14678 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 39526 14678 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 39445 14678 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 39364 14678 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 39283 14678 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 39202 14678 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 39121 14678 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 39040 14678 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 38959 14678 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 38879 14678 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 38799 14678 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 38719 14678 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 38639 14678 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 38559 14678 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 38479 14678 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 38399 14678 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 38319 14678 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 38239 14678 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 38159 14678 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 38079 14678 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 37999 14678 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 37919 14678 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 37839 14678 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 37759 14678 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 37679 14678 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 37599 14678 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 37519 14678 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 37439 14678 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 37359 14678 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 37279 14678 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 37199 14678 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 37119 14678 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 37039 14678 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 36959 14678 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 36879 14678 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 36799 14678 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 36719 14678 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 36639 14678 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 36559 14678 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 36479 14678 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 36399 14678 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 36319 14678 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 36239 14678 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 36159 14678 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 36079 14678 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 35999 14678 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 35919 14678 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 35839 14678 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 35759 14678 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 35679 14678 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 35599 14678 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 35519 14678 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 35439 14678 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 35359 14678 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 35279 14678 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 35199 14678 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 6042 14678 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 5956 14678 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 5870 14678 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 5784 14678 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 5698 14678 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 5612 14678 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 5526 14678 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 5440 14678 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 5354 14678 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 5268 14678 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14638 5182 14678 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 39931 14598 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 39850 14598 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 39769 14598 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 39688 14598 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 39607 14598 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 39526 14598 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 39445 14598 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 39364 14598 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 39283 14598 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 39202 14598 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 39121 14598 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 39040 14598 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 38959 14598 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 38879 14598 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 38799 14598 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 38719 14598 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 38639 14598 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 38559 14598 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 38479 14598 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 38399 14598 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 38319 14598 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 38239 14598 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 38159 14598 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 38079 14598 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 37999 14598 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 37919 14598 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 37839 14598 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 37759 14598 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 37679 14598 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 37599 14598 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 37519 14598 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 37439 14598 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 37359 14598 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 37279 14598 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 37199 14598 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 37119 14598 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 37039 14598 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 36959 14598 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 36879 14598 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 36799 14598 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 36719 14598 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 36639 14598 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 36559 14598 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 36479 14598 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 36399 14598 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 36319 14598 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 36239 14598 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 36159 14598 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 36079 14598 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 35999 14598 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 35919 14598 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 35839 14598 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 35759 14598 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 35679 14598 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 35599 14598 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 35519 14598 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 35439 14598 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 35359 14598 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 35279 14598 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14558 35199 14598 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 6042 14597 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5956 14597 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5870 14597 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5784 14597 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5698 14597 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5612 14597 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5526 14597 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5440 14597 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5354 14597 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5268 14597 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14557 5182 14597 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 39931 14518 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 39850 14518 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 39769 14518 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 39688 14518 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 39607 14518 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 39526 14518 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 39445 14518 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 39364 14518 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 39283 14518 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 39202 14518 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 39121 14518 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 39040 14518 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 38959 14518 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 38879 14518 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 38799 14518 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 38719 14518 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 38639 14518 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 38559 14518 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 38479 14518 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 38399 14518 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 38319 14518 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 38239 14518 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 38159 14518 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 38079 14518 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 37999 14518 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 37919 14518 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 37839 14518 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 37759 14518 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 37679 14518 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 37599 14518 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 37519 14518 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 37439 14518 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 37359 14518 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 37279 14518 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 37199 14518 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 37119 14518 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 37039 14518 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 36959 14518 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 36879 14518 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 36799 14518 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 36719 14518 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 36639 14518 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 36559 14518 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 36479 14518 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 36399 14518 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 36319 14518 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 36239 14518 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 36159 14518 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 36079 14518 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 35999 14518 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 35919 14518 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 35839 14518 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 35759 14518 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 35679 14518 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 35599 14518 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 35519 14518 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 35439 14518 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 35359 14518 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 35279 14518 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14478 35199 14518 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14476 6042 14516 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14476 5956 14516 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14476 5870 14516 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14476 5784 14516 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14476 5698 14516 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14476 5612 14516 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14476 5526 14516 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14476 5440 14516 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14476 5354 14516 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14476 5268 14516 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14476 5182 14516 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 39931 14438 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 39850 14438 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 39769 14438 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 39688 14438 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 39607 14438 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 39526 14438 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 39445 14438 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 39364 14438 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 39283 14438 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 39202 14438 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 39121 14438 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 39040 14438 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 38959 14438 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 38879 14438 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 38799 14438 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 38719 14438 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 38639 14438 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 38559 14438 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 38479 14438 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 38399 14438 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 38319 14438 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 38239 14438 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 38159 14438 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 38079 14438 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 37999 14438 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 37919 14438 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 37839 14438 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 37759 14438 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 37679 14438 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 37599 14438 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 37519 14438 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 37439 14438 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 37359 14438 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 37279 14438 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 37199 14438 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 37119 14438 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 37039 14438 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 36959 14438 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 36879 14438 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 36799 14438 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 36719 14438 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 36639 14438 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 36559 14438 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 36479 14438 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 36399 14438 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 36319 14438 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 36239 14438 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 36159 14438 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 36079 14438 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 35999 14438 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 35919 14438 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 35839 14438 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 35759 14438 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 35679 14438 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 35599 14438 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 35519 14438 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 35439 14438 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 35359 14438 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 35279 14438 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14398 35199 14438 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14395 6042 14435 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14395 5956 14435 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14395 5870 14435 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14395 5784 14435 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14395 5698 14435 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14395 5612 14435 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14395 5526 14435 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14395 5440 14435 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14395 5354 14435 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14395 5268 14435 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14395 5182 14435 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 39931 14358 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 39850 14358 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 39769 14358 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 39688 14358 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 39607 14358 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 39526 14358 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 39445 14358 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 39364 14358 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 39283 14358 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 39202 14358 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 39121 14358 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 39040 14358 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 38959 14358 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 38879 14358 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 38799 14358 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 38719 14358 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 38639 14358 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 38559 14358 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 38479 14358 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 38399 14358 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 38319 14358 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 38239 14358 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 38159 14358 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 38079 14358 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 37999 14358 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 37919 14358 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 37839 14358 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 37759 14358 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 37679 14358 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 37599 14358 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 37519 14358 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 37439 14358 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 37359 14358 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 37279 14358 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 37199 14358 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 37119 14358 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 37039 14358 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 36959 14358 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 36879 14358 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 36799 14358 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 36719 14358 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 36639 14358 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 36559 14358 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 36479 14358 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 36399 14358 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 36319 14358 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 36239 14358 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 36159 14358 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 36079 14358 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 35999 14358 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 35919 14358 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 35839 14358 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 35759 14358 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 35679 14358 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 35599 14358 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 35519 14358 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 35439 14358 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 35359 14358 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 35279 14358 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14318 35199 14358 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14314 6042 14354 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14314 5956 14354 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14314 5870 14354 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14314 5784 14354 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14314 5698 14354 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14314 5612 14354 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14314 5526 14354 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14314 5440 14354 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14314 5354 14354 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14314 5268 14354 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14314 5182 14354 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 39931 14278 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 39850 14278 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 39769 14278 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 39688 14278 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 39607 14278 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 39526 14278 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 39445 14278 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 39364 14278 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 39283 14278 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 39202 14278 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 39121 14278 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 39040 14278 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 38959 14278 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 38879 14278 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 38799 14278 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 38719 14278 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 38639 14278 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 38559 14278 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 38479 14278 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 38399 14278 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 38319 14278 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 38239 14278 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 38159 14278 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 38079 14278 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 37999 14278 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 37919 14278 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 37839 14278 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 37759 14278 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 37679 14278 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 37599 14278 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 37519 14278 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 37439 14278 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 37359 14278 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 37279 14278 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 37199 14278 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 37119 14278 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 37039 14278 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 36959 14278 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 36879 14278 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 36799 14278 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 36719 14278 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 36639 14278 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 36559 14278 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 36479 14278 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 36399 14278 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 36319 14278 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 36239 14278 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 36159 14278 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 36079 14278 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 35999 14278 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 35919 14278 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 35839 14278 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 35759 14278 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 35679 14278 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 35599 14278 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 35519 14278 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 35439 14278 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 35359 14278 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 35279 14278 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14238 35199 14278 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 6042 14273 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5956 14273 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5870 14273 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5784 14273 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5698 14273 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5612 14273 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5526 14273 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5440 14273 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5354 14273 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5268 14273 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14233 5182 14273 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 39931 14198 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 39850 14198 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 39769 14198 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 39688 14198 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 39607 14198 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 39526 14198 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 39445 14198 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 39364 14198 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 39283 14198 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 39202 14198 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 39121 14198 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 39040 14198 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 38959 14198 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 38879 14198 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 38799 14198 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 38719 14198 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 38639 14198 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 38559 14198 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 38479 14198 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 38399 14198 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 38319 14198 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 38239 14198 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 38159 14198 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 38079 14198 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 37999 14198 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 37919 14198 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 37839 14198 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 37759 14198 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 37679 14198 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 37599 14198 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 37519 14198 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 37439 14198 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 37359 14198 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 37279 14198 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 37199 14198 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 37119 14198 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 37039 14198 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 36959 14198 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 36879 14198 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 36799 14198 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 36719 14198 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 36639 14198 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 36559 14198 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 36479 14198 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 36399 14198 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 36319 14198 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 36239 14198 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 36159 14198 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 36079 14198 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 35999 14198 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 35919 14198 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 35839 14198 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 35759 14198 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 35679 14198 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 35599 14198 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 35519 14198 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 35439 14198 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 35359 14198 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 35279 14198 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14158 35199 14198 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14152 6042 14192 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14152 5956 14192 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14152 5870 14192 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14152 5784 14192 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14152 5698 14192 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14152 5612 14192 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14152 5526 14192 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14152 5440 14192 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14152 5354 14192 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14152 5268 14192 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14152 5182 14192 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 39931 14118 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 39850 14118 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 39769 14118 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 39688 14118 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 39607 14118 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 39526 14118 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 39445 14118 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 39364 14118 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 39283 14118 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 39202 14118 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 39121 14118 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 39040 14118 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 38959 14118 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 38879 14118 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 38799 14118 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 38719 14118 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 38639 14118 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 38559 14118 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 38479 14118 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 38399 14118 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 38319 14118 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 38239 14118 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 38159 14118 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 38079 14118 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 37999 14118 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 37919 14118 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 37839 14118 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 37759 14118 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 37679 14118 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 37599 14118 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 37519 14118 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 37439 14118 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 37359 14118 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 37279 14118 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 37199 14118 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 37119 14118 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 37039 14118 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 36959 14118 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 36879 14118 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 36799 14118 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 36719 14118 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 36639 14118 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 36559 14118 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 36479 14118 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 36399 14118 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 36319 14118 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 36239 14118 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 36159 14118 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 36079 14118 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 35999 14118 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 35919 14118 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 35839 14118 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 35759 14118 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 35679 14118 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 35599 14118 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 35519 14118 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 35439 14118 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 35359 14118 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 35279 14118 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14078 35199 14118 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14071 6042 14111 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14071 5956 14111 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14071 5870 14111 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14071 5784 14111 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14071 5698 14111 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14071 5612 14111 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14071 5526 14111 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14071 5440 14111 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14071 5354 14111 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14071 5268 14111 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 14071 5182 14111 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 39931 14038 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 39850 14038 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 39769 14038 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 39688 14038 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 39607 14038 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 39526 14038 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 39445 14038 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 39364 14038 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 39283 14038 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 39202 14038 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 39121 14038 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 39040 14038 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 38959 14038 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 38879 14038 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 38799 14038 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 38719 14038 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 38639 14038 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 38559 14038 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 38479 14038 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 38399 14038 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 38319 14038 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 38239 14038 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 38159 14038 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 38079 14038 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 37999 14038 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 37919 14038 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 37839 14038 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 37759 14038 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 37679 14038 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 37599 14038 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 37519 14038 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 37439 14038 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 37359 14038 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 37279 14038 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 37199 14038 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 37119 14038 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 37039 14038 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 36959 14038 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 36879 14038 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 36799 14038 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 36719 14038 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 36639 14038 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 36559 14038 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 36479 14038 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 36399 14038 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 36319 14038 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 36239 14038 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 36159 14038 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 36079 14038 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 35999 14038 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 35919 14038 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 35839 14038 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 35759 14038 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 35679 14038 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 35599 14038 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 35519 14038 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 35439 14038 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 35359 14038 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 35279 14038 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13998 35199 14038 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13990 6042 14030 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13990 5956 14030 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13990 5870 14030 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13990 5784 14030 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13990 5698 14030 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13990 5612 14030 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13990 5526 14030 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13990 5440 14030 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13990 5354 14030 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13990 5268 14030 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13990 5182 14030 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 39931 13958 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 39850 13958 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 39769 13958 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 39688 13958 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 39607 13958 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 39526 13958 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 39445 13958 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 39364 13958 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 39283 13958 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 39202 13958 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 39121 13958 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 39040 13958 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 38959 13958 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 38879 13958 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 38799 13958 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 38719 13958 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 38639 13958 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 38559 13958 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 38479 13958 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 38399 13958 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 38319 13958 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 38239 13958 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 38159 13958 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 38079 13958 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 37999 13958 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 37919 13958 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 37839 13958 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 37759 13958 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 37679 13958 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 37599 13958 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 37519 13958 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 37439 13958 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 37359 13958 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 37279 13958 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 37199 13958 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 37119 13958 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 37039 13958 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 36959 13958 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 36879 13958 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 36799 13958 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 36719 13958 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 36639 13958 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 36559 13958 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 36479 13958 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 36399 13958 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 36319 13958 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 36239 13958 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 36159 13958 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 36079 13958 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 35999 13958 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 35919 13958 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 35839 13958 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 35759 13958 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 35679 13958 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 35599 13958 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 35519 13958 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 35439 13958 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 35359 13958 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 35279 13958 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13918 35199 13958 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 6042 13949 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5956 13949 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5870 13949 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5784 13949 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5698 13949 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5612 13949 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5526 13949 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5440 13949 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5354 13949 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5268 13949 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13909 5182 13949 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 39931 13878 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 39850 13878 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 39769 13878 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 39688 13878 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 39607 13878 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 39526 13878 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 39445 13878 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 39364 13878 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 39283 13878 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 39202 13878 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 39121 13878 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 39040 13878 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 38959 13878 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 38879 13878 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 38799 13878 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 38719 13878 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 38639 13878 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 38559 13878 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 38479 13878 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 38399 13878 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 38319 13878 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 38239 13878 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 38159 13878 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 38079 13878 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 37999 13878 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 37919 13878 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 37839 13878 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 37759 13878 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 37679 13878 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 37599 13878 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 37519 13878 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 37439 13878 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 37359 13878 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 37279 13878 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 37199 13878 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 37119 13878 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 37039 13878 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 36959 13878 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 36879 13878 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 36799 13878 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 36719 13878 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 36639 13878 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 36559 13878 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 36479 13878 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 36399 13878 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 36319 13878 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 36239 13878 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 36159 13878 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 36079 13878 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 35999 13878 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 35919 13878 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 35839 13878 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 35759 13878 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 35679 13878 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 35599 13878 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 35519 13878 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 35439 13878 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 35359 13878 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 35279 13878 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13838 35199 13878 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13828 6042 13868 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13828 5956 13868 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13828 5870 13868 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13828 5784 13868 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13828 5698 13868 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13828 5612 13868 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13828 5526 13868 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13828 5440 13868 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13828 5354 13868 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13828 5268 13868 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13828 5182 13868 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 39931 13798 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 39850 13798 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 39769 13798 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 39688 13798 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 39607 13798 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 39526 13798 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 39445 13798 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 39364 13798 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 39283 13798 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 39202 13798 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 39121 13798 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 39040 13798 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 38959 13798 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 38879 13798 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 38799 13798 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 38719 13798 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 38639 13798 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 38559 13798 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 38479 13798 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 38399 13798 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 38319 13798 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 38239 13798 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 38159 13798 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 38079 13798 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 37999 13798 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 37919 13798 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 37839 13798 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 37759 13798 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 37679 13798 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 37599 13798 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 37519 13798 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 37439 13798 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 37359 13798 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 37279 13798 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 37199 13798 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 37119 13798 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 37039 13798 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 36959 13798 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 36879 13798 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 36799 13798 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 36719 13798 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 36639 13798 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 36559 13798 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 36479 13798 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 36399 13798 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 36319 13798 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 36239 13798 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 36159 13798 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 36079 13798 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 35999 13798 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 35919 13798 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 35839 13798 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 35759 13798 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 35679 13798 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 35599 13798 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 35519 13798 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 35439 13798 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 35359 13798 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 35279 13798 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13758 35199 13798 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13747 6042 13787 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13747 5956 13787 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13747 5870 13787 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13747 5784 13787 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13747 5698 13787 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13747 5612 13787 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13747 5526 13787 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13747 5440 13787 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13747 5354 13787 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13747 5268 13787 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13747 5182 13787 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 39931 13718 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 39850 13718 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 39769 13718 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 39688 13718 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 39607 13718 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 39526 13718 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 39445 13718 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 39364 13718 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 39283 13718 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 39202 13718 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 39121 13718 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 39040 13718 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 38959 13718 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 38879 13718 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 38799 13718 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 38719 13718 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 38639 13718 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 38559 13718 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 38479 13718 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 38399 13718 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 38319 13718 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 38239 13718 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 38159 13718 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 38079 13718 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 37999 13718 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 37919 13718 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 37839 13718 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 37759 13718 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 37679 13718 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 37599 13718 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 37519 13718 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 37439 13718 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 37359 13718 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 37279 13718 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 37199 13718 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 37119 13718 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 37039 13718 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 36959 13718 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 36879 13718 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 36799 13718 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 36719 13718 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 36639 13718 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 36559 13718 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 36479 13718 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 36399 13718 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 36319 13718 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 36239 13718 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 36159 13718 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 36079 13718 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 35999 13718 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 35919 13718 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 35839 13718 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 35759 13718 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 35679 13718 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 35599 13718 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 35519 13718 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 35439 13718 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 35359 13718 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 35279 13718 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13678 35199 13718 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 6042 13706 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 5956 13706 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 5870 13706 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 5784 13706 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 5698 13706 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 5612 13706 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 5526 13706 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 5440 13706 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 5354 13706 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 5268 13706 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13666 5182 13706 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 39931 13638 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 39850 13638 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 39769 13638 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 39688 13638 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 39607 13638 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 39526 13638 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 39445 13638 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 39364 13638 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 39283 13638 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 39202 13638 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 39121 13638 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 39040 13638 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 38959 13638 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 38879 13638 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 38799 13638 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 38719 13638 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 38639 13638 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 38559 13638 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 38479 13638 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 38399 13638 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 38319 13638 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 38239 13638 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 38159 13638 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 38079 13638 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 37999 13638 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 37919 13638 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 37839 13638 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 37759 13638 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 37679 13638 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 37599 13638 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 37519 13638 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 37439 13638 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 37359 13638 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 37279 13638 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 37199 13638 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 37119 13638 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 37039 13638 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 36959 13638 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 36879 13638 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 36799 13638 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 36719 13638 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 36639 13638 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 36559 13638 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 36479 13638 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 36399 13638 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 36319 13638 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 36239 13638 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 36159 13638 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 36079 13638 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 35999 13638 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 35919 13638 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 35839 13638 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 35759 13638 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 35679 13638 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 35599 13638 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 35519 13638 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 35439 13638 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 35359 13638 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 35279 13638 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13598 35199 13638 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 6042 13625 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5956 13625 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5870 13625 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5784 13625 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5698 13625 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5612 13625 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5526 13625 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5440 13625 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5354 13625 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5268 13625 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13585 5182 13625 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 39931 13558 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 39850 13558 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 39769 13558 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 39688 13558 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 39607 13558 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 39526 13558 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 39445 13558 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 39364 13558 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 39283 13558 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 39202 13558 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 39121 13558 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 39040 13558 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 38959 13558 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 38879 13558 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 38799 13558 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 38719 13558 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 38639 13558 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 38559 13558 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 38479 13558 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 38399 13558 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 38319 13558 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 38239 13558 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 38159 13558 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 38079 13558 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 37999 13558 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 37919 13558 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 37839 13558 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 37759 13558 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 37679 13558 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 37599 13558 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 37519 13558 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 37439 13558 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 37359 13558 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 37279 13558 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 37199 13558 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 37119 13558 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 37039 13558 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 36959 13558 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 36879 13558 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 36799 13558 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 36719 13558 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 36639 13558 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 36559 13558 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 36479 13558 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 36399 13558 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 36319 13558 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 36239 13558 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 36159 13558 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 36079 13558 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 35999 13558 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 35919 13558 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 35839 13558 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 35759 13558 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 35679 13558 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 35599 13558 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 35519 13558 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 35439 13558 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 35359 13558 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 35279 13558 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13518 35199 13558 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13504 6042 13544 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13504 5956 13544 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13504 5870 13544 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13504 5784 13544 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13504 5698 13544 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13504 5612 13544 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13504 5526 13544 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13504 5440 13544 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13504 5354 13544 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13504 5268 13544 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13504 5182 13544 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 39931 13478 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 39850 13478 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 39769 13478 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 39688 13478 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 39607 13478 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 39526 13478 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 39445 13478 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 39364 13478 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 39283 13478 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 39202 13478 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 39121 13478 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 39040 13478 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 38959 13478 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 38879 13478 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 38799 13478 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 38719 13478 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 38639 13478 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 38559 13478 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 38479 13478 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 38399 13478 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 38319 13478 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 38239 13478 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 38159 13478 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 38079 13478 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 37999 13478 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 37919 13478 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 37839 13478 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 37759 13478 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 37679 13478 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 37599 13478 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 37519 13478 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 37439 13478 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 37359 13478 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 37279 13478 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 37199 13478 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 37119 13478 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 37039 13478 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 36959 13478 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 36879 13478 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 36799 13478 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 36719 13478 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 36639 13478 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 36559 13478 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 36479 13478 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 36399 13478 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 36319 13478 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 36239 13478 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 36159 13478 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 36079 13478 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 35999 13478 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 35919 13478 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 35839 13478 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 35759 13478 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 35679 13478 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 35599 13478 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 35519 13478 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 35439 13478 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 35359 13478 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 35279 13478 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13438 35199 13478 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13423 6042 13463 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13423 5956 13463 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13423 5870 13463 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13423 5784 13463 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13423 5698 13463 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13423 5612 13463 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13423 5526 13463 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13423 5440 13463 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13423 5354 13463 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13423 5268 13463 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13423 5182 13463 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 39931 13398 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 39850 13398 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 39769 13398 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 39688 13398 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 39607 13398 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 39526 13398 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 39445 13398 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 39364 13398 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 39283 13398 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 39202 13398 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 39121 13398 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 39040 13398 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 38959 13398 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 38879 13398 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 38799 13398 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 38719 13398 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 38639 13398 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 38559 13398 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 38479 13398 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 38399 13398 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 38319 13398 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 38239 13398 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 38159 13398 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 38079 13398 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 37999 13398 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 37919 13398 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 37839 13398 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 37759 13398 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 37679 13398 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 37599 13398 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 37519 13398 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 37439 13398 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 37359 13398 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 37279 13398 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 37199 13398 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 37119 13398 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 37039 13398 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 36959 13398 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 36879 13398 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 36799 13398 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 36719 13398 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 36639 13398 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 36559 13398 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 36479 13398 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 36399 13398 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 36319 13398 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 36239 13398 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 36159 13398 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 36079 13398 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 35999 13398 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 35919 13398 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 35839 13398 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 35759 13398 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 35679 13398 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 35599 13398 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 35519 13398 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 35439 13398 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 35359 13398 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 35279 13398 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13358 35199 13398 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13342 6042 13382 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13342 5956 13382 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13342 5870 13382 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13342 5784 13382 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13342 5698 13382 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13342 5612 13382 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13342 5526 13382 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13342 5440 13382 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13342 5354 13382 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13342 5268 13382 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13342 5182 13382 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 39931 13318 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 39850 13318 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 39769 13318 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 39688 13318 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 39607 13318 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 39526 13318 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 39445 13318 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 39364 13318 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 39283 13318 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 39202 13318 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 39121 13318 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 39040 13318 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 38959 13318 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 38879 13318 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 38799 13318 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 38719 13318 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 38639 13318 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 38559 13318 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 38479 13318 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 38399 13318 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 38319 13318 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 38239 13318 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 38159 13318 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 38079 13318 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 37999 13318 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 37919 13318 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 37839 13318 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 37759 13318 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 37679 13318 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 37599 13318 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 37519 13318 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 37439 13318 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 37359 13318 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 37279 13318 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 37199 13318 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 37119 13318 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 37039 13318 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 36959 13318 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 36879 13318 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 36799 13318 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 36719 13318 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 36639 13318 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 36559 13318 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 36479 13318 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 36399 13318 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 36319 13318 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 36239 13318 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 36159 13318 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 36079 13318 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 35999 13318 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 35919 13318 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 35839 13318 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 35759 13318 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 35679 13318 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 35599 13318 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 35519 13318 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 35439 13318 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 35359 13318 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 35279 13318 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13278 35199 13318 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 6042 13301 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5956 13301 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5870 13301 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5784 13301 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5698 13301 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5612 13301 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5526 13301 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5440 13301 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5354 13301 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5268 13301 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13261 5182 13301 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 39931 13238 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 39850 13238 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 39769 13238 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 39688 13238 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 39607 13238 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 39526 13238 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 39445 13238 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 39364 13238 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 39283 13238 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 39202 13238 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 39121 13238 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 39040 13238 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 38959 13238 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 38879 13238 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 38799 13238 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 38719 13238 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 38639 13238 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 38559 13238 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 38479 13238 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 38399 13238 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 38319 13238 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 38239 13238 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 38159 13238 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 38079 13238 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 37999 13238 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 37919 13238 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 37839 13238 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 37759 13238 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 37679 13238 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 37599 13238 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 37519 13238 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 37439 13238 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 37359 13238 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 37279 13238 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 37199 13238 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 37119 13238 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 37039 13238 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 36959 13238 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 36879 13238 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 36799 13238 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 36719 13238 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 36639 13238 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 36559 13238 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 36479 13238 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 36399 13238 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 36319 13238 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 36239 13238 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 36159 13238 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 36079 13238 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 35999 13238 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 35919 13238 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 35839 13238 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 35759 13238 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 35679 13238 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 35599 13238 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 35519 13238 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 35439 13238 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 35359 13238 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 35279 13238 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13198 35199 13238 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13180 6042 13220 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13180 5956 13220 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13180 5870 13220 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13180 5784 13220 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13180 5698 13220 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13180 5612 13220 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13180 5526 13220 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13180 5440 13220 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13180 5354 13220 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13180 5268 13220 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13180 5182 13220 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 39931 13158 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 39850 13158 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 39769 13158 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 39688 13158 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 39607 13158 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 39526 13158 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 39445 13158 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 39364 13158 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 39283 13158 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 39202 13158 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 39121 13158 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 39040 13158 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 38959 13158 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 38879 13158 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 38799 13158 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 38719 13158 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 38639 13158 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 38559 13158 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 38479 13158 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 38399 13158 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 38319 13158 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 38239 13158 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 38159 13158 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 38079 13158 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 37999 13158 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 37919 13158 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 37839 13158 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 37759 13158 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 37679 13158 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 37599 13158 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 37519 13158 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 37439 13158 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 37359 13158 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 37279 13158 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 37199 13158 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 37119 13158 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 37039 13158 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 36959 13158 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 36879 13158 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 36799 13158 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 36719 13158 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 36639 13158 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 36559 13158 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 36479 13158 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 36399 13158 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 36319 13158 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 36239 13158 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 36159 13158 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 36079 13158 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 35999 13158 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 35919 13158 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 35839 13158 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 35759 13158 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 35679 13158 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 35599 13158 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 35519 13158 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 35439 13158 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 35359 13158 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 35279 13158 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13118 35199 13158 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13099 6042 13139 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13099 5956 13139 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13099 5870 13139 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13099 5784 13139 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13099 5698 13139 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13099 5612 13139 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13099 5526 13139 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13099 5440 13139 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13099 5354 13139 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13099 5268 13139 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13099 5182 13139 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 39931 13078 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 39850 13078 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 39769 13078 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 39688 13078 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 39607 13078 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 39526 13078 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 39445 13078 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 39364 13078 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 39283 13078 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 39202 13078 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 39121 13078 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 39040 13078 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 38959 13078 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 38879 13078 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 38799 13078 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 38719 13078 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 38639 13078 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 38559 13078 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 38479 13078 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 38399 13078 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 38319 13078 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 38239 13078 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 38159 13078 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 38079 13078 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 37999 13078 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 37919 13078 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 37839 13078 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 37759 13078 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 37679 13078 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 37599 13078 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 37519 13078 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 37439 13078 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 37359 13078 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 37279 13078 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 37199 13078 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 37119 13078 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 37039 13078 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 36959 13078 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 36879 13078 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 36799 13078 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 36719 13078 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 36639 13078 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 36559 13078 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 36479 13078 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 36399 13078 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 36319 13078 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 36239 13078 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 36159 13078 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 36079 13078 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 35999 13078 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 35919 13078 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 35839 13078 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 35759 13078 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 35679 13078 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 35599 13078 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 35519 13078 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 35439 13078 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 35359 13078 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 35279 13078 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13038 35199 13078 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13018 6042 13058 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13018 5956 13058 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13018 5870 13058 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13018 5784 13058 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13018 5698 13058 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13018 5612 13058 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13018 5526 13058 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13018 5440 13058 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13018 5354 13058 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13018 5268 13058 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 13018 5182 13058 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 39931 12998 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 39850 12998 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 39769 12998 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 39688 12998 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 39607 12998 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 39526 12998 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 39445 12998 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 39364 12998 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 39283 12998 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 39202 12998 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 39121 12998 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 39040 12998 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 38959 12998 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 38879 12998 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 38799 12998 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 38719 12998 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 38639 12998 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 38559 12998 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 38479 12998 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 38399 12998 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 38319 12998 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 38239 12998 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 38159 12998 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 38079 12998 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 37999 12998 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 37919 12998 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 37839 12998 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 37759 12998 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 37679 12998 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 37599 12998 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 37519 12998 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 37439 12998 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 37359 12998 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 37279 12998 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 37199 12998 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 37119 12998 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 37039 12998 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 36959 12998 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 36879 12998 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 36799 12998 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 36719 12998 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 36639 12998 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 36559 12998 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 36479 12998 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 36399 12998 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 36319 12998 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 36239 12998 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 36159 12998 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 36079 12998 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 35999 12998 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 35919 12998 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 35839 12998 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 35759 12998 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 35679 12998 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 35599 12998 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 35519 12998 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 35439 12998 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 35359 12998 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 35279 12998 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12958 35199 12998 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 6042 12977 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5956 12977 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5870 12977 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5784 12977 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5698 12977 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5612 12977 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5526 12977 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5440 12977 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5354 12977 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5268 12977 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12937 5182 12977 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 39931 12918 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 39850 12918 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 39769 12918 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 39688 12918 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 39607 12918 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 39526 12918 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 39445 12918 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 39364 12918 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 39283 12918 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 39202 12918 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 39121 12918 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 39040 12918 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 38959 12918 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 38879 12918 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 38799 12918 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 38719 12918 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 38639 12918 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 38559 12918 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 38479 12918 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 38399 12918 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 38319 12918 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 38239 12918 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 38159 12918 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 38079 12918 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 37999 12918 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 37919 12918 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 37839 12918 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 37759 12918 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 37679 12918 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 37599 12918 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 37519 12918 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 37439 12918 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 37359 12918 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 37279 12918 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 37199 12918 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 37119 12918 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 37039 12918 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 36959 12918 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 36879 12918 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 36799 12918 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 36719 12918 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 36639 12918 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 36559 12918 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 36479 12918 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 36399 12918 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 36319 12918 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 36239 12918 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 36159 12918 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 36079 12918 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 35999 12918 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 35919 12918 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 35839 12918 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 35759 12918 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 35679 12918 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 35599 12918 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 35519 12918 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 35439 12918 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 35359 12918 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 35279 12918 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12878 35199 12918 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12856 6042 12896 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12856 5956 12896 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12856 5870 12896 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12856 5784 12896 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12856 5698 12896 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12856 5612 12896 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12856 5526 12896 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12856 5440 12896 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12856 5354 12896 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12856 5268 12896 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12856 5182 12896 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 39931 12838 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 39850 12838 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 39769 12838 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 39688 12838 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 39607 12838 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 39526 12838 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 39445 12838 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 39364 12838 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 39283 12838 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 39202 12838 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 39121 12838 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 39040 12838 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 38959 12838 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 38879 12838 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 38799 12838 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 38719 12838 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 38639 12838 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 38559 12838 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 38479 12838 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 38399 12838 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 38319 12838 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 38239 12838 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 38159 12838 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 38079 12838 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 37999 12838 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 37919 12838 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 37839 12838 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 37759 12838 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 37679 12838 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 37599 12838 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 37519 12838 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 37439 12838 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 37359 12838 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 37279 12838 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 37199 12838 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 37119 12838 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 37039 12838 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 36959 12838 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 36879 12838 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 36799 12838 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 36719 12838 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 36639 12838 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 36559 12838 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 36479 12838 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 36399 12838 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 36319 12838 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 36239 12838 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 36159 12838 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 36079 12838 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 35999 12838 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 35919 12838 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 35839 12838 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 35759 12838 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 35679 12838 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 35599 12838 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 35519 12838 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 35439 12838 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 35359 12838 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 35279 12838 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12798 35199 12838 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12775 6042 12815 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12775 5956 12815 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12775 5870 12815 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12775 5784 12815 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12775 5698 12815 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12775 5612 12815 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12775 5526 12815 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12775 5440 12815 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12775 5354 12815 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12775 5268 12815 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12775 5182 12815 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 39931 12758 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 39850 12758 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 39769 12758 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 39688 12758 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 39607 12758 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 39526 12758 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 39445 12758 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 39364 12758 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 39283 12758 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 39202 12758 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 39121 12758 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 39040 12758 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 38959 12758 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 38879 12758 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 38799 12758 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 38719 12758 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 38639 12758 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 38559 12758 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 38479 12758 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 38399 12758 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 38319 12758 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 38239 12758 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 38159 12758 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 38079 12758 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 37999 12758 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 37919 12758 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 37839 12758 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 37759 12758 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 37679 12758 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 37599 12758 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 37519 12758 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 37439 12758 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 37359 12758 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 37279 12758 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 37199 12758 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 37119 12758 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 37039 12758 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 36959 12758 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 36879 12758 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 36799 12758 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 36719 12758 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 36639 12758 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 36559 12758 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 36479 12758 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 36399 12758 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 36319 12758 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 36239 12758 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 36159 12758 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 36079 12758 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 35999 12758 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 35919 12758 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 35839 12758 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 35759 12758 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 35679 12758 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 35599 12758 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 35519 12758 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 35439 12758 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 35359 12758 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 35279 12758 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12718 35199 12758 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12694 6042 12734 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12694 5956 12734 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12694 5870 12734 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12694 5784 12734 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12694 5698 12734 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12694 5612 12734 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12694 5526 12734 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12694 5440 12734 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12694 5354 12734 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12694 5268 12734 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12694 5182 12734 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 39931 12678 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 39850 12678 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 39769 12678 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 39688 12678 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 39607 12678 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 39526 12678 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 39445 12678 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 39364 12678 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 39283 12678 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 39202 12678 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 39121 12678 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 39040 12678 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 38959 12678 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 38879 12678 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 38799 12678 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 38719 12678 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 38639 12678 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 38559 12678 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 38479 12678 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 38399 12678 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 38319 12678 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 38239 12678 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 38159 12678 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 38079 12678 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 37999 12678 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 37919 12678 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 37839 12678 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 37759 12678 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 37679 12678 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 37599 12678 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 37519 12678 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 37439 12678 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 37359 12678 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 37279 12678 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 37199 12678 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 37119 12678 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 37039 12678 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 36959 12678 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 36879 12678 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 36799 12678 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 36719 12678 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 36639 12678 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 36559 12678 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 36479 12678 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 36399 12678 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 36319 12678 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 36239 12678 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 36159 12678 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 36079 12678 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 35999 12678 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 35919 12678 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 35839 12678 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 35759 12678 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 35679 12678 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 35599 12678 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 35519 12678 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 35439 12678 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 35359 12678 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 35279 12678 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12638 35199 12678 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 6042 12653 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5956 12653 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5870 12653 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5784 12653 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5698 12653 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5612 12653 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5526 12653 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5440 12653 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5354 12653 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5268 12653 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12613 5182 12653 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 39931 12598 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 39850 12598 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 39769 12598 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 39688 12598 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 39607 12598 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 39526 12598 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 39445 12598 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 39364 12598 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 39283 12598 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 39202 12598 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 39121 12598 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 39040 12598 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 38959 12598 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 38879 12598 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 38799 12598 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 38719 12598 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 38639 12598 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 38559 12598 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 38479 12598 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 38399 12598 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 38319 12598 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 38239 12598 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 38159 12598 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 38079 12598 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 37999 12598 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 37919 12598 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 37839 12598 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 37759 12598 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 37679 12598 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 37599 12598 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 37519 12598 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 37439 12598 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 37359 12598 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 37279 12598 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 37199 12598 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 37119 12598 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 37039 12598 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 36959 12598 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 36879 12598 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 36799 12598 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 36719 12598 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 36639 12598 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 36559 12598 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 36479 12598 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 36399 12598 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 36319 12598 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 36239 12598 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 36159 12598 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 36079 12598 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 35999 12598 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 35919 12598 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 35839 12598 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 35759 12598 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 35679 12598 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 35599 12598 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 35519 12598 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 35439 12598 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 35359 12598 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 35279 12598 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12558 35199 12598 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12532 6042 12572 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12532 5956 12572 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12532 5870 12572 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12532 5784 12572 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12532 5698 12572 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12532 5612 12572 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12532 5526 12572 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12532 5440 12572 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12532 5354 12572 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12532 5268 12572 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12532 5182 12572 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 39931 12518 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 39850 12518 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 39769 12518 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 39688 12518 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 39607 12518 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 39526 12518 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 39445 12518 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 39364 12518 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 39283 12518 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 39202 12518 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 39121 12518 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 39040 12518 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 38959 12518 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 38879 12518 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 38799 12518 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 38719 12518 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 38639 12518 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 38559 12518 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 38479 12518 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 38399 12518 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 38319 12518 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 38239 12518 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 38159 12518 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 38079 12518 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 37999 12518 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 37919 12518 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 37839 12518 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 37759 12518 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 37679 12518 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 37599 12518 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 37519 12518 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 37439 12518 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 37359 12518 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 37279 12518 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 37199 12518 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 37119 12518 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 37039 12518 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 36959 12518 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 36879 12518 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 36799 12518 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 36719 12518 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 36639 12518 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 36559 12518 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 36479 12518 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 36399 12518 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 36319 12518 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 36239 12518 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 36159 12518 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 36079 12518 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 35999 12518 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 35919 12518 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 35839 12518 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 35759 12518 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 35679 12518 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 35599 12518 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 35519 12518 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 35439 12518 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 35359 12518 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 35279 12518 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12478 35199 12518 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12451 6042 12491 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12451 5956 12491 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12451 5870 12491 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12451 5784 12491 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12451 5698 12491 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12451 5612 12491 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12451 5526 12491 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12451 5440 12491 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12451 5354 12491 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12451 5268 12491 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12451 5182 12491 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 39931 12438 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 39850 12438 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 39769 12438 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 39688 12438 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 39607 12438 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 39526 12438 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 39445 12438 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 39364 12438 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 39283 12438 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 39202 12438 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 39121 12438 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 39040 12438 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 38959 12438 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 38879 12438 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 38799 12438 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 38719 12438 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 38639 12438 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 38559 12438 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 38479 12438 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 38399 12438 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 38319 12438 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 38239 12438 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 38159 12438 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 38079 12438 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 37999 12438 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 37919 12438 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 37839 12438 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 37759 12438 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 37679 12438 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 37599 12438 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 37519 12438 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 37439 12438 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 37359 12438 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 37279 12438 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 37199 12438 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 37119 12438 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 37039 12438 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 36959 12438 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 36879 12438 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 36799 12438 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 36719 12438 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 36639 12438 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 36559 12438 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 36479 12438 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 36399 12438 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 36319 12438 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 36239 12438 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 36159 12438 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 36079 12438 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 35999 12438 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 35919 12438 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 35839 12438 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 35759 12438 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 35679 12438 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 35599 12438 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 35519 12438 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 35439 12438 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 35359 12438 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 35279 12438 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12398 35199 12438 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12370 6042 12410 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12370 5956 12410 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12370 5870 12410 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12370 5784 12410 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12370 5698 12410 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12370 5612 12410 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12370 5526 12410 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12370 5440 12410 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12370 5354 12410 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12370 5268 12410 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12370 5182 12410 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 39931 12358 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 39850 12358 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 39769 12358 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 39688 12358 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 39607 12358 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 39526 12358 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 39445 12358 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 39364 12358 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 39283 12358 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 39202 12358 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 39121 12358 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 39040 12358 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 38959 12358 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 38879 12358 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 38799 12358 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 38719 12358 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 38639 12358 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 38559 12358 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 38479 12358 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 38399 12358 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 38319 12358 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 38239 12358 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 38159 12358 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 38079 12358 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 37999 12358 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 37919 12358 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 37839 12358 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 37759 12358 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 37679 12358 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 37599 12358 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 37519 12358 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 37439 12358 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 37359 12358 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 37279 12358 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 37199 12358 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 37119 12358 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 37039 12358 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 36959 12358 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 36879 12358 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 36799 12358 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 36719 12358 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 36639 12358 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 36559 12358 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 36479 12358 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 36399 12358 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 36319 12358 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 36239 12358 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 36159 12358 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 36079 12358 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 35999 12358 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 35919 12358 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 35839 12358 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 35759 12358 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 35679 12358 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 35599 12358 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 35519 12358 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 35439 12358 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 35359 12358 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 35279 12358 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12318 35199 12358 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 6042 12329 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5956 12329 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5870 12329 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5784 12329 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5698 12329 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5612 12329 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5526 12329 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5440 12329 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5354 12329 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5268 12329 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12289 5182 12329 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12212 39930 12252 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12212 39850 12252 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12212 39770 12252 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12212 39690 12252 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12212 39610 12252 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12212 39530 12252 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12212 39450 12252 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12208 6042 12248 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12208 5956 12248 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12208 5870 12248 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12208 5784 12248 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12208 5698 12248 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12208 5612 12248 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12208 5526 12248 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12208 5440 12248 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12208 5354 12248 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12208 5268 12248 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12208 5182 12248 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12182 39341 12222 39381 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12182 39259 12222 39299 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12132 39930 12172 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12132 39850 12172 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12132 39770 12172 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12132 39690 12172 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12132 39610 12172 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12132 39530 12172 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12132 39450 12172 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12127 6042 12167 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12127 5956 12167 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12127 5870 12167 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12127 5784 12167 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12127 5698 12167 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12127 5612 12167 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12127 5526 12167 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12127 5440 12167 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12127 5354 12167 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12127 5268 12167 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12127 5182 12167 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12052 39930 12092 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12052 39850 12092 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12052 39770 12092 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12052 39690 12092 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12052 39610 12092 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12052 39530 12092 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12052 39450 12092 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12046 6042 12086 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12046 5956 12086 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12046 5870 12086 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12046 5784 12086 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12046 5698 12086 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12046 5612 12086 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12046 5526 12086 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12046 5440 12086 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12046 5354 12086 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12046 5268 12086 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 12046 5182 12086 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11972 39930 12012 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11972 39850 12012 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11972 39770 12012 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11972 39690 12012 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11972 39610 12012 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11972 39530 12012 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11972 39450 12012 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 6042 12005 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5956 12005 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5870 12005 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5784 12005 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5698 12005 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5612 12005 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5526 12005 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5440 12005 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5354 12005 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5268 12005 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11965 5182 12005 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11892 39930 11932 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11892 39850 11932 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11892 39770 11932 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11892 39690 11932 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11892 39610 11932 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11892 39530 11932 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11892 39450 11932 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11884 6042 11924 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11884 5956 11924 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11884 5870 11924 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11884 5784 11924 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11884 5698 11924 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11884 5612 11924 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11884 5526 11924 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11884 5440 11924 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11884 5354 11924 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11884 5268 11924 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11884 5182 11924 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11812 39930 11852 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11812 39850 11852 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11812 39770 11852 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11812 39690 11852 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11812 39610 11852 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11812 39530 11852 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11812 39450 11852 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11803 6042 11843 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11803 5956 11843 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11803 5870 11843 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11803 5784 11843 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11803 5698 11843 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11803 5612 11843 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11803 5526 11843 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11803 5440 11843 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11803 5354 11843 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11803 5268 11843 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11803 5182 11843 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11732 39930 11772 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11732 39850 11772 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11732 39770 11772 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11732 39690 11772 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11732 39610 11772 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11732 39530 11772 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11732 39450 11772 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11722 6042 11762 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11722 5956 11762 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11722 5870 11762 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11722 5784 11762 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11722 5698 11762 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11722 5612 11762 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11722 5526 11762 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11722 5440 11762 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11722 5354 11762 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11722 5268 11762 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11722 5182 11762 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11652 39930 11692 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11652 39850 11692 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11652 39770 11692 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11652 39690 11692 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11652 39610 11692 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11652 39530 11692 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11652 39450 11692 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 6042 11681 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5956 11681 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5870 11681 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5784 11681 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5698 11681 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5612 11681 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5526 11681 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5440 11681 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5354 11681 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5268 11681 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11641 5182 11681 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11572 39930 11612 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11572 39850 11612 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11572 39770 11612 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11572 39690 11612 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11572 39610 11612 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11572 39530 11612 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11572 39450 11612 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11560 6042 11600 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11560 5956 11600 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11560 5870 11600 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11560 5784 11600 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11560 5698 11600 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11560 5612 11600 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11560 5526 11600 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11560 5440 11600 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11560 5354 11600 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11560 5268 11600 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11560 5182 11600 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11492 39930 11532 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11492 39850 11532 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11492 39770 11532 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11492 39690 11532 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11492 39610 11532 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11492 39530 11532 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11492 39450 11532 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11479 6042 11519 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11479 5956 11519 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11479 5870 11519 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11479 5784 11519 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11479 5698 11519 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11479 5612 11519 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11479 5526 11519 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11479 5440 11519 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11479 5354 11519 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11479 5268 11519 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11479 5182 11519 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11412 39930 11452 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11412 39850 11452 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11412 39770 11452 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11412 39690 11452 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11412 39610 11452 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11412 39530 11452 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11412 39450 11452 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11398 6042 11438 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11398 5956 11438 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11398 5870 11438 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11398 5784 11438 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11398 5698 11438 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11398 5612 11438 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11398 5526 11438 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11398 5440 11438 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11398 5354 11438 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11398 5268 11438 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11398 5182 11438 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11332 39930 11372 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11332 39850 11372 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11332 39770 11372 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11332 39690 11372 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11332 39610 11372 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11332 39530 11372 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11332 39450 11372 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 6042 11357 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5956 11357 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5870 11357 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5784 11357 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5698 11357 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5612 11357 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5526 11357 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5440 11357 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5354 11357 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5268 11357 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11317 5182 11357 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11252 39930 11292 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11252 39850 11292 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11252 39770 11292 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11252 39690 11292 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11252 39610 11292 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11252 39530 11292 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11252 39450 11292 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11236 6042 11276 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11236 5956 11276 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11236 5870 11276 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11236 5784 11276 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11236 5698 11276 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11236 5612 11276 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11236 5526 11276 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11236 5440 11276 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11236 5354 11276 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11236 5268 11276 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11236 5182 11276 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11172 39930 11212 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11172 39850 11212 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11172 39770 11212 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11172 39690 11212 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11172 39610 11212 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11172 39530 11212 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11172 39450 11212 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11155 6042 11195 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11155 5956 11195 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11155 5870 11195 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11155 5784 11195 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11155 5698 11195 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11155 5612 11195 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11155 5526 11195 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11155 5440 11195 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11155 5354 11195 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11155 5268 11195 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11155 5182 11195 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11092 39930 11132 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11092 39850 11132 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11092 39770 11132 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11092 39690 11132 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11092 39610 11132 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11092 39530 11132 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11092 39450 11132 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11074 6042 11114 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11074 5956 11114 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11074 5870 11114 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11074 5784 11114 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11074 5698 11114 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11074 5612 11114 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11074 5526 11114 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11074 5440 11114 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11074 5354 11114 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11074 5268 11114 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11074 5182 11114 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11012 39930 11052 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11012 39850 11052 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11012 39770 11052 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11012 39690 11052 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11012 39610 11052 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11012 39530 11052 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 11012 39450 11052 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 6042 11033 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5956 11033 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5870 11033 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5784 11033 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5698 11033 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5612 11033 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5526 11033 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5440 11033 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5354 11033 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5268 11033 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10993 5182 11033 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10932 39930 10972 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10932 39850 10972 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10932 39770 10972 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10932 39690 10972 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10932 39610 10972 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10932 39530 10972 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10932 39450 10972 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10912 6042 10952 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10912 5956 10952 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10912 5870 10952 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10912 5784 10952 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10912 5698 10952 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10912 5612 10952 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10912 5526 10952 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10912 5440 10952 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10912 5354 10952 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10912 5268 10952 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10912 5182 10952 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10852 39930 10892 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10852 39850 10892 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10852 39770 10892 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10852 39690 10892 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10852 39610 10892 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10852 39530 10892 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10852 39450 10892 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10831 6042 10871 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10831 5956 10871 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10831 5870 10871 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10831 5784 10871 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10831 5698 10871 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10831 5612 10871 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10831 5526 10871 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10831 5440 10871 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10831 5354 10871 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10831 5268 10871 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10831 5182 10871 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10772 39930 10812 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10772 39850 10812 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10772 39770 10812 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10772 39690 10812 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10772 39610 10812 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10772 39530 10812 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10772 39450 10812 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10750 6042 10790 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10750 5956 10790 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10750 5870 10790 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10750 5784 10790 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10750 5698 10790 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10750 5612 10790 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10750 5526 10790 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10750 5440 10790 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10750 5354 10790 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10750 5268 10790 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10750 5182 10790 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10692 39930 10732 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10692 39850 10732 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10692 39770 10732 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10692 39690 10732 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10692 39610 10732 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10692 39530 10732 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10692 39450 10732 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 6042 10709 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5956 10709 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5870 10709 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5784 10709 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5698 10709 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5612 10709 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5526 10709 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5440 10709 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5354 10709 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5268 10709 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10669 5182 10709 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10612 39930 10652 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10612 39850 10652 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10612 39770 10652 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10612 39690 10652 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10612 39610 10652 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10612 39530 10652 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10612 39450 10652 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10588 6042 10628 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10588 5956 10628 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10588 5870 10628 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10588 5784 10628 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10588 5698 10628 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10588 5612 10628 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10588 5526 10628 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10588 5440 10628 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10588 5354 10628 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10588 5268 10628 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10588 5182 10628 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10532 39930 10572 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10532 39850 10572 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10532 39770 10572 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10532 39690 10572 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10532 39610 10572 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10532 39530 10572 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10532 39450 10572 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10506 6042 10546 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10506 5956 10546 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10506 5870 10546 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10506 5784 10546 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10506 5698 10546 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10506 5612 10546 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10506 5526 10546 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10506 5440 10546 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10506 5354 10546 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10506 5268 10546 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10506 5182 10546 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10452 39930 10492 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10452 39850 10492 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10452 39770 10492 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10452 39690 10492 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10452 39610 10492 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10452 39530 10492 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10452 39450 10492 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10424 6042 10464 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10424 5956 10464 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10424 5870 10464 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10424 5784 10464 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10424 5698 10464 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10424 5612 10464 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10424 5526 10464 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10424 5440 10464 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10424 5354 10464 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10424 5268 10464 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10424 5182 10464 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10372 39930 10412 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10372 39850 10412 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10372 39770 10412 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10372 39690 10412 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10372 39610 10412 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10372 39530 10412 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10372 39450 10412 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 6042 10382 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5956 10382 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5870 10382 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5784 10382 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5698 10382 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5612 10382 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5526 10382 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5440 10382 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5354 10382 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5268 10382 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10342 5182 10382 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10292 39930 10332 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10292 39850 10332 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10292 39770 10332 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10292 39690 10332 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10292 39610 10332 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10292 39530 10332 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10292 39450 10332 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10260 6042 10300 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10260 5956 10300 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10260 5870 10300 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10260 5784 10300 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10260 5698 10300 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10260 5612 10300 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10260 5526 10300 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10260 5440 10300 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10260 5354 10300 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10260 5268 10300 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10260 5182 10300 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10212 39930 10252 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10212 39850 10252 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10212 39770 10252 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10212 39690 10252 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10212 39610 10252 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10212 39530 10252 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10212 39450 10252 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10178 6042 10218 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10178 5956 10218 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10178 5870 10218 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10178 5784 10218 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10178 5698 10218 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10178 5612 10218 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10178 5526 10218 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10178 5440 10218 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10178 5354 10218 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10178 5268 10218 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10178 5182 10218 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10132 39930 10172 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10132 39850 10172 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10132 39770 10172 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10132 39690 10172 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10132 39610 10172 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10132 39530 10172 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10132 39450 10172 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10096 6042 10136 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10096 5956 10136 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10096 5870 10136 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10096 5784 10136 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10096 5698 10136 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10096 5612 10136 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10096 5526 10136 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10096 5440 10136 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10096 5354 10136 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10096 5268 10136 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10096 5182 10136 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10052 39930 10092 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10052 39850 10092 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10052 39770 10092 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10052 39690 10092 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10052 39610 10092 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10052 39530 10092 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 10052 39450 10092 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9972 39930 10012 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9972 39850 10012 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9972 39770 10012 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9972 39690 10012 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9972 39610 10012 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9972 39530 10012 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9972 39450 10012 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9892 39930 9932 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9892 39850 9932 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9892 39770 9932 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9892 39690 9932 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9892 39610 9932 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9892 39530 9932 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9892 39450 9932 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9812 39930 9852 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9812 39850 9852 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9812 39770 9852 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9812 39690 9852 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9812 39610 9852 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9812 39530 9852 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9812 39450 9852 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9732 39930 9772 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9732 39850 9772 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9732 39770 9772 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9732 39690 9772 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9732 39610 9772 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9732 39530 9772 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9732 39450 9772 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9652 39930 9692 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9652 39850 9692 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9652 39770 9692 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9652 39690 9692 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9652 39610 9692 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9652 39530 9692 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9652 39450 9692 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9572 39930 9612 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9572 39850 9612 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9572 39770 9612 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9572 39690 9612 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9572 39610 9612 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9572 39530 9612 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9572 39450 9612 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9492 39930 9532 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9492 39850 9532 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9492 39770 9532 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9492 39690 9532 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9492 39610 9532 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9492 39530 9532 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9492 39450 9532 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9412 39930 9452 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9412 39850 9452 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9412 39770 9452 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9412 39690 9452 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9412 39610 9452 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9412 39530 9452 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9412 39450 9452 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9332 39930 9372 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9332 39850 9372 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9332 39770 9372 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9332 39690 9372 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9332 39610 9372 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9332 39530 9372 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9332 39450 9372 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9252 39930 9292 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9252 39850 9292 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9252 39770 9292 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9252 39690 9292 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9252 39610 9292 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9252 39530 9292 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9252 39450 9292 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9172 39930 9212 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9172 39850 9212 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9172 39770 9212 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9172 39690 9212 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9172 39610 9212 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9172 39530 9212 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9172 39450 9212 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9092 39930 9132 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9092 39850 9132 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9092 39770 9132 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9092 39690 9132 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9092 39610 9132 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9092 39530 9132 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9092 39450 9132 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9012 39930 9052 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9012 39850 9052 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9012 39770 9052 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9012 39690 9052 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9012 39610 9052 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9012 39530 9052 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 9012 39450 9052 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8932 39930 8972 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8932 39850 8972 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8932 39770 8972 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8932 39690 8972 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8932 39610 8972 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8932 39530 8972 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8932 39450 8972 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8852 39930 8892 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8852 39850 8892 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8852 39770 8892 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8852 39690 8892 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8852 39610 8892 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8852 39530 8892 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8852 39450 8892 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8772 39930 8812 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8772 39850 8812 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8772 39770 8812 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8772 39690 8812 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8772 39610 8812 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8772 39530 8812 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8772 39450 8812 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8692 39930 8732 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8692 39850 8732 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8692 39770 8732 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8692 39690 8732 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8692 39610 8732 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8692 39530 8732 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8692 39450 8732 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8612 39930 8652 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8612 39850 8652 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8612 39770 8652 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8612 39690 8652 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8612 39610 8652 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8612 39530 8652 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8612 39450 8652 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8532 39930 8572 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8532 39850 8572 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8532 39770 8572 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8532 39690 8572 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8532 39610 8572 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8532 39530 8572 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8532 39450 8572 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8452 39930 8492 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8452 39850 8492 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8452 39770 8492 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8452 39690 8492 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8452 39610 8492 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8452 39530 8492 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8452 39450 8492 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8372 39930 8412 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8372 39850 8412 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8372 39770 8412 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8372 39690 8412 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8372 39610 8412 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8372 39530 8412 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8372 39450 8412 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8292 39930 8332 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8292 39850 8332 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8292 39770 8332 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8292 39690 8332 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8292 39610 8332 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8292 39530 8332 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8292 39450 8332 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8212 39930 8252 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8212 39850 8252 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8212 39770 8252 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8212 39690 8252 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8212 39610 8252 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8212 39530 8252 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8212 39450 8252 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8132 39930 8172 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8132 39850 8172 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8132 39770 8172 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8132 39690 8172 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8132 39610 8172 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8132 39530 8172 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8132 39450 8172 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8052 39930 8092 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8052 39850 8092 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8052 39770 8092 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8052 39690 8092 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8052 39610 8092 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8052 39530 8092 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 8052 39450 8092 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7972 39930 8012 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7972 39850 8012 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7972 39770 8012 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7972 39690 8012 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7972 39610 8012 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7972 39530 8012 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7972 39450 8012 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7892 39930 7932 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7892 39850 7932 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7892 39770 7932 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7892 39690 7932 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7892 39610 7932 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7892 39530 7932 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7892 39450 7932 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7812 39930 7852 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7812 39850 7852 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7812 39770 7852 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7812 39690 7852 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7812 39610 7852 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7812 39530 7852 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7812 39450 7852 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7732 39930 7772 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7732 39850 7772 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7732 39770 7772 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7732 39690 7772 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7732 39610 7772 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7732 39530 7772 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7732 39450 7772 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7652 39930 7692 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7652 39850 7692 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7652 39770 7692 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7652 39690 7692 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7652 39610 7692 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7652 39530 7692 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7652 39450 7692 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7572 39930 7612 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7572 39850 7612 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7572 39770 7612 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7572 39690 7612 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7572 39610 7612 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7572 39530 7612 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7572 39450 7612 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7492 39930 7532 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7492 39850 7532 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7492 39770 7532 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7492 39690 7532 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7492 39610 7532 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7492 39530 7532 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7492 39450 7532 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7412 39930 7452 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7412 39850 7452 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7412 39770 7452 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7412 39690 7452 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7412 39610 7452 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7412 39530 7452 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7412 39450 7452 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7332 39930 7372 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7332 39850 7372 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7332 39770 7372 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7332 39690 7372 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7332 39610 7372 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7332 39530 7372 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7332 39450 7372 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7252 39930 7292 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7252 39850 7292 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7252 39770 7292 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7252 39690 7292 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7252 39610 7292 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7252 39530 7292 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7252 39450 7292 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7172 39930 7212 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7172 39850 7212 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7172 39770 7212 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7172 39690 7212 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7172 39610 7212 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7172 39530 7212 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7172 39450 7212 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7092 39930 7132 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7092 39850 7132 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7092 39770 7132 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7092 39690 7132 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7092 39610 7132 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7092 39530 7132 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7092 39450 7132 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7012 39930 7052 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7012 39850 7052 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7012 39770 7052 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7012 39690 7052 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7012 39610 7052 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7012 39530 7052 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 7012 39450 7052 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6932 39930 6972 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6932 39850 6972 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6932 39770 6972 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6932 39690 6972 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6932 39610 6972 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6932 39530 6972 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6932 39450 6972 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6852 39930 6892 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6852 39850 6892 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6852 39770 6892 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6852 39690 6892 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6852 39610 6892 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6852 39530 6892 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6852 39450 6892 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6772 39930 6812 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6772 39850 6812 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6772 39770 6812 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6772 39690 6812 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6772 39610 6812 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6772 39530 6812 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6772 39450 6812 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6692 39930 6732 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6692 39850 6732 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6692 39770 6732 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6692 39690 6732 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6692 39610 6732 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6692 39530 6732 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6692 39450 6732 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6612 39930 6652 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6612 39850 6652 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6612 39770 6652 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6612 39690 6652 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6612 39610 6652 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6612 39530 6652 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6612 39450 6652 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6532 39930 6572 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6532 39850 6572 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6532 39770 6572 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6532 39690 6572 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6532 39610 6572 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6532 39530 6572 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6532 39450 6572 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6452 39930 6492 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6452 39850 6492 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6452 39770 6492 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6452 39690 6492 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6452 39610 6492 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6452 39530 6492 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6452 39450 6492 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6372 39930 6412 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6372 39850 6412 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6372 39770 6412 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6372 39690 6412 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6372 39610 6412 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6372 39530 6412 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6372 39450 6412 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6292 39930 6332 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6292 39850 6332 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6292 39770 6332 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6292 39690 6332 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6292 39610 6332 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6292 39530 6332 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6292 39450 6332 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6212 39930 6252 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6212 39850 6252 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6212 39770 6252 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6212 39690 6252 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6212 39610 6252 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6212 39530 6252 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6212 39450 6252 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6132 39930 6172 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6132 39850 6172 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6132 39770 6172 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6132 39690 6172 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6132 39610 6172 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6132 39530 6172 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6132 39450 6172 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6052 39930 6092 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6052 39850 6092 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6052 39770 6092 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6052 39690 6092 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6052 39610 6092 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6052 39530 6092 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 6052 39450 6092 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5972 39930 6012 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5972 39850 6012 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5972 39770 6012 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5972 39690 6012 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5972 39610 6012 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5972 39530 6012 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5972 39450 6012 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5892 39930 5932 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5892 39850 5932 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5892 39770 5932 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5892 39690 5932 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5892 39610 5932 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5892 39530 5932 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5892 39450 5932 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5812 39930 5852 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5812 39850 5852 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5812 39770 5852 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5812 39690 5852 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5812 39610 5852 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5812 39530 5852 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5812 39450 5852 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5732 39930 5772 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5732 39850 5772 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5732 39770 5772 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5732 39690 5772 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5732 39610 5772 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5732 39530 5772 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5732 39450 5772 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5652 39930 5692 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5652 39850 5692 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5652 39770 5692 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5652 39690 5692 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5652 39610 5692 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5652 39530 5692 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5652 39450 5692 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5572 39930 5612 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5572 39850 5612 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5572 39770 5612 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5572 39690 5612 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5572 39610 5612 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5572 39530 5612 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5572 39450 5612 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5492 39930 5532 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5492 39850 5532 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5492 39770 5532 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5492 39690 5532 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5492 39610 5532 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5492 39530 5532 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5492 39450 5532 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5412 39930 5452 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5412 39850 5452 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5412 39770 5452 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5412 39690 5452 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5412 39610 5452 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5412 39530 5452 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5412 39450 5452 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5331 39930 5371 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5331 39850 5371 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5331 39770 5371 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5331 39690 5371 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5331 39610 5371 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5331 39530 5371 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5331 39450 5371 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5250 39930 5290 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5250 39850 5290 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5250 39770 5290 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5250 39690 5290 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5250 39610 5290 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5250 39530 5290 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5250 39450 5290 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5169 39930 5209 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5169 39850 5209 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5169 39770 5209 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5169 39690 5209 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5169 39610 5209 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5169 39530 5209 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5169 39450 5209 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5088 39930 5128 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5088 39850 5128 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5088 39770 5128 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5088 39690 5128 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5088 39610 5128 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5088 39530 5128 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5088 39450 5128 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5007 39930 5047 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5007 39850 5047 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5007 39770 5047 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5007 39690 5047 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5007 39610 5047 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5007 39530 5047 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 5007 39450 5047 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4926 39930 4966 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4926 39850 4966 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4926 39770 4966 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4926 39690 4966 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4926 39610 4966 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4926 39530 4966 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4926 39450 4966 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4845 39930 4885 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4845 39850 4885 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4845 39770 4885 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4845 39690 4885 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4845 39610 4885 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4845 39530 4885 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4845 39450 4885 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4821 6042 4861 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4821 5956 4861 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4821 5870 4861 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4821 5784 4861 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4821 5698 4861 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4821 5612 4861 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4821 5526 4861 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4821 5440 4861 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4821 5354 4861 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4821 5268 4861 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4821 5182 4861 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4764 39930 4804 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4764 39850 4804 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4764 39770 4804 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4764 39690 4804 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4764 39610 4804 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4764 39530 4804 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4764 39450 4804 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4740 6042 4780 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4740 5956 4780 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4740 5870 4780 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4740 5784 4780 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4740 5698 4780 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4740 5612 4780 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4740 5526 4780 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4740 5440 4780 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4740 5354 4780 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4740 5268 4780 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4740 5182 4780 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4683 39930 4723 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4683 39850 4723 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4683 39770 4723 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4683 39690 4723 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4683 39610 4723 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4683 39530 4723 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4683 39450 4723 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4659 6042 4699 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4659 5956 4699 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4659 5870 4699 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4659 5784 4699 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4659 5698 4699 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4659 5612 4699 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4659 5526 4699 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4659 5440 4699 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4659 5354 4699 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4659 5268 4699 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4659 5182 4699 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4602 39930 4642 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4602 39850 4642 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4602 39770 4642 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4602 39690 4642 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4602 39610 4642 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4602 39530 4642 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4602 39450 4642 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 6042 4618 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5956 4618 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5870 4618 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5784 4618 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5698 4618 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5612 4618 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5526 4618 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5440 4618 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5354 4618 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5268 4618 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4578 5182 4618 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4521 39930 4561 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4521 39850 4561 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4521 39770 4561 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4521 39690 4561 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4521 39610 4561 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4521 39530 4561 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4521 39450 4561 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4497 6042 4537 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4497 5956 4537 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4497 5870 4537 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4497 5784 4537 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4497 5698 4537 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4497 5612 4537 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4497 5526 4537 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4497 5440 4537 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4497 5354 4537 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4497 5268 4537 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4497 5182 4537 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4440 39930 4480 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4440 39850 4480 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4440 39770 4480 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4440 39690 4480 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4440 39610 4480 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4440 39530 4480 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4440 39450 4480 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4416 6042 4456 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4416 5956 4456 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4416 5870 4456 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4416 5784 4456 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4416 5698 4456 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4416 5612 4456 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4416 5526 4456 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4416 5440 4456 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4416 5354 4456 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4416 5268 4456 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4416 5182 4456 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4359 39930 4399 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4359 39850 4399 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4359 39770 4399 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4359 39690 4399 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4359 39610 4399 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4359 39530 4399 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4359 39450 4399 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4335 6042 4375 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4335 5956 4375 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4335 5870 4375 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4335 5784 4375 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4335 5698 4375 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4335 5612 4375 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4335 5526 4375 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4335 5440 4375 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4335 5354 4375 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4335 5268 4375 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4335 5182 4375 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4278 39930 4318 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4278 39850 4318 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4278 39770 4318 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4278 39690 4318 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4278 39610 4318 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4278 39530 4318 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4278 39450 4318 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 6042 4294 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5956 4294 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5870 4294 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5784 4294 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5698 4294 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5612 4294 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5526 4294 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5440 4294 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5354 4294 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5268 4294 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4254 5182 4294 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4197 39930 4237 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4197 39850 4237 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4197 39770 4237 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4197 39690 4237 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4197 39610 4237 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4197 39530 4237 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4197 39450 4237 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4173 6042 4213 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4173 5956 4213 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4173 5870 4213 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4173 5784 4213 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4173 5698 4213 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4173 5612 4213 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4173 5526 4213 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4173 5440 4213 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4173 5354 4213 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4173 5268 4213 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4173 5182 4213 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4116 39930 4156 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4116 39850 4156 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4116 39770 4156 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4116 39690 4156 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4116 39610 4156 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4116 39530 4156 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4116 39450 4156 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4092 6042 4132 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4092 5956 4132 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4092 5870 4132 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4092 5784 4132 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4092 5698 4132 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4092 5612 4132 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4092 5526 4132 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4092 5440 4132 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4092 5354 4132 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4092 5268 4132 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4092 5182 4132 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4035 39930 4075 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4035 39850 4075 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4035 39770 4075 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4035 39690 4075 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4035 39610 4075 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4035 39530 4075 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4035 39450 4075 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4011 6042 4051 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4011 5956 4051 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4011 5870 4051 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4011 5784 4051 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4011 5698 4051 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4011 5612 4051 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4011 5526 4051 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4011 5440 4051 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4011 5354 4051 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4011 5268 4051 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 4011 5182 4051 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3954 39930 3994 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3954 39850 3994 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3954 39770 3994 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3954 39690 3994 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3954 39610 3994 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3954 39530 3994 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3954 39450 3994 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 6042 3970 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5956 3970 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5870 3970 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5784 3970 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5698 3970 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5612 3970 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5526 3970 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5440 3970 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5354 3970 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5268 3970 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3930 5182 3970 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3873 39930 3913 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3873 39850 3913 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3873 39770 3913 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3873 39690 3913 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3873 39610 3913 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3873 39530 3913 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3873 39450 3913 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3849 6042 3889 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3849 5956 3889 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3849 5870 3889 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3849 5784 3889 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3849 5698 3889 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3849 5612 3889 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3849 5526 3889 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3849 5440 3889 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3849 5354 3889 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3849 5268 3889 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3849 5182 3889 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3792 39930 3832 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3792 39850 3832 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3792 39770 3832 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3792 39690 3832 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3792 39610 3832 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3792 39530 3832 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3792 39450 3832 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3768 6042 3808 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3768 5956 3808 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3768 5870 3808 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3768 5784 3808 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3768 5698 3808 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3768 5612 3808 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3768 5526 3808 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3768 5440 3808 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3768 5354 3808 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3768 5268 3808 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3768 5182 3808 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3711 39930 3751 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3711 39850 3751 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3711 39770 3751 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3711 39690 3751 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3711 39610 3751 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3711 39530 3751 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3711 39450 3751 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3687 6042 3727 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3687 5956 3727 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3687 5870 3727 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3687 5784 3727 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3687 5698 3727 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3687 5612 3727 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3687 5526 3727 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3687 5440 3727 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3687 5354 3727 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3687 5268 3727 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3687 5182 3727 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3630 39930 3670 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3630 39850 3670 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3630 39770 3670 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3630 39690 3670 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3630 39610 3670 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3630 39530 3670 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3630 39450 3670 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 6042 3646 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5956 3646 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5870 3646 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5784 3646 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5698 3646 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5612 3646 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5526 3646 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5440 3646 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5354 3646 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5268 3646 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3606 5182 3646 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3549 39930 3589 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3549 39850 3589 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3549 39770 3589 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3549 39690 3589 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3549 39610 3589 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3549 39530 3589 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3549 39450 3589 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3525 6042 3565 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3525 5956 3565 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3525 5870 3565 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3525 5784 3565 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3525 5698 3565 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3525 5612 3565 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3525 5526 3565 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3525 5440 3565 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3525 5354 3565 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3525 5268 3565 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3525 5182 3565 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3468 39930 3508 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3468 39850 3508 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3468 39770 3508 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3468 39690 3508 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3468 39610 3508 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3468 39530 3508 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3468 39450 3508 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3444 6042 3484 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3444 5956 3484 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3444 5870 3484 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3444 5784 3484 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3444 5698 3484 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3444 5612 3484 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3444 5526 3484 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3444 5440 3484 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3444 5354 3484 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3444 5268 3484 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3444 5182 3484 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3387 39930 3427 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3387 39850 3427 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3387 39770 3427 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3387 39690 3427 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3387 39610 3427 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3387 39530 3427 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3387 39450 3427 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3363 6042 3403 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3363 5956 3403 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3363 5870 3403 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3363 5784 3403 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3363 5698 3403 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3363 5612 3403 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3363 5526 3403 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3363 5440 3403 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3363 5354 3403 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3363 5268 3403 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3363 5182 3403 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3306 39930 3346 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3306 39850 3346 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3306 39770 3346 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3306 39690 3346 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3306 39610 3346 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3306 39530 3346 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3306 39450 3346 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 6042 3322 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5956 3322 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5870 3322 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5784 3322 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5698 3322 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5612 3322 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5526 3322 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5440 3322 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5354 3322 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5268 3322 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3282 5182 3322 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3225 39930 3265 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3225 39850 3265 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3225 39770 3265 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3225 39690 3265 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3225 39610 3265 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3225 39530 3265 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3225 39450 3265 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3201 6042 3241 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3201 5956 3241 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3201 5870 3241 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3201 5784 3241 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3201 5698 3241 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3201 5612 3241 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3201 5526 3241 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3201 5440 3241 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3201 5354 3241 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3201 5268 3241 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3201 5182 3241 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3144 39930 3184 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3144 39850 3184 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3144 39770 3184 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3144 39690 3184 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3144 39610 3184 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3144 39530 3184 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3144 39450 3184 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3120 6042 3160 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3120 5956 3160 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3120 5870 3160 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3120 5784 3160 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3120 5698 3160 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3120 5612 3160 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3120 5526 3160 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3120 5440 3160 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3120 5354 3160 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3120 5268 3160 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3120 5182 3160 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3063 39930 3103 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3063 39850 3103 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3063 39770 3103 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3063 39690 3103 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3063 39610 3103 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3063 39530 3103 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3063 39450 3103 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3039 6042 3079 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3039 5956 3079 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3039 5870 3079 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3039 5784 3079 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3039 5698 3079 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3039 5612 3079 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3039 5526 3079 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3039 5440 3079 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3039 5354 3079 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3039 5268 3079 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 3039 5182 3079 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2982 39930 3022 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2982 39850 3022 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2982 39770 3022 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2982 39690 3022 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2982 39610 3022 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2982 39530 3022 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2982 39450 3022 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 6042 2998 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5956 2998 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5870 2998 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5784 2998 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5698 2998 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5612 2998 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5526 2998 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5440 2998 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5354 2998 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5268 2998 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2958 5182 2998 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2901 39930 2941 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2901 39850 2941 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2901 39770 2941 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2901 39690 2941 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2901 39610 2941 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2901 39530 2941 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2901 39450 2941 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2877 6042 2917 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2877 5956 2917 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2877 5870 2917 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2877 5784 2917 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2877 5698 2917 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2877 5612 2917 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2877 5526 2917 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2877 5440 2917 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2877 5354 2917 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2877 5268 2917 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2877 5182 2917 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2820 39930 2860 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2820 39850 2860 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2820 39770 2860 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2820 39690 2860 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2820 39610 2860 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2820 39530 2860 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2820 39450 2860 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2796 6042 2836 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2796 5956 2836 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2796 5870 2836 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2796 5784 2836 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2796 5698 2836 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2796 5612 2836 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2796 5526 2836 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2796 5440 2836 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2796 5354 2836 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2796 5268 2836 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2796 5182 2836 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2765 39341 2805 39381 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2765 39259 2805 39299 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2739 39930 2779 39970 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2739 39850 2779 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2739 39770 2779 39810 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2739 39690 2779 39730 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2739 39610 2779 39650 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2739 39530 2779 39570 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2739 39450 2779 39490 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2715 6042 2755 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2715 5956 2755 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2715 5870 2755 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2715 5784 2755 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2715 5698 2755 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2715 5612 2755 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2715 5526 2755 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2715 5440 2755 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2715 5354 2755 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2715 5268 2755 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2715 5182 2755 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 6042 2674 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5956 2674 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5870 2674 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5784 2674 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5698 2674 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5612 2674 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5526 2674 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5440 2674 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5354 2674 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5268 2674 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2634 5182 2674 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 39931 2657 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 39850 2657 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 39769 2657 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 39688 2657 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 39607 2657 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 39526 2657 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 39445 2657 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 39364 2657 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 39283 2657 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 39202 2657 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 39121 2657 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 39040 2657 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 38959 2657 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 38879 2657 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 38799 2657 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 38719 2657 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 38639 2657 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 38559 2657 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 38479 2657 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 38399 2657 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 38319 2657 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 38239 2657 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 38159 2657 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 38079 2657 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 37999 2657 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 37919 2657 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 37839 2657 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 37759 2657 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 37679 2657 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 37599 2657 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 37519 2657 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 37439 2657 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 37359 2657 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 37279 2657 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 37199 2657 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 37119 2657 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 37039 2657 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 36959 2657 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 36879 2657 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 36799 2657 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 36719 2657 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 36639 2657 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 36559 2657 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 36479 2657 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 36399 2657 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 36319 2657 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 36239 2657 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 36159 2657 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 36079 2657 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 35999 2657 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 35919 2657 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 35839 2657 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 35759 2657 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 35679 2657 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 35599 2657 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 35519 2657 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 35439 2657 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 35359 2657 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 35279 2657 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2617 35199 2657 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2553 6042 2593 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2553 5956 2593 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2553 5870 2593 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2553 5784 2593 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2553 5698 2593 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2553 5612 2593 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2553 5526 2593 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2553 5440 2593 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2553 5354 2593 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2553 5268 2593 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2553 5182 2593 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 39931 2577 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 39850 2577 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 39769 2577 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 39688 2577 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 39607 2577 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 39526 2577 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 39445 2577 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 39364 2577 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 39283 2577 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 39202 2577 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 39121 2577 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 39040 2577 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 38959 2577 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 38879 2577 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 38799 2577 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 38719 2577 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 38639 2577 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 38559 2577 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 38479 2577 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 38399 2577 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 38319 2577 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 38239 2577 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 38159 2577 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 38079 2577 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 37999 2577 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 37919 2577 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 37839 2577 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 37759 2577 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 37679 2577 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 37599 2577 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 37519 2577 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 37439 2577 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 37359 2577 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 37279 2577 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 37199 2577 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 37119 2577 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 37039 2577 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 36959 2577 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 36879 2577 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 36799 2577 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 36719 2577 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 36639 2577 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 36559 2577 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 36479 2577 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 36399 2577 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 36319 2577 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 36239 2577 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 36159 2577 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 36079 2577 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 35999 2577 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 35919 2577 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 35839 2577 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 35759 2577 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 35679 2577 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 35599 2577 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 35519 2577 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 35439 2577 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 35359 2577 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 35279 2577 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2537 35199 2577 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2472 6042 2512 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2472 5956 2512 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2472 5870 2512 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2472 5784 2512 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2472 5698 2512 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2472 5612 2512 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2472 5526 2512 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2472 5440 2512 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2472 5354 2512 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2472 5268 2512 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2472 5182 2512 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 39931 2497 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 39850 2497 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 39769 2497 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 39688 2497 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 39607 2497 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 39526 2497 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 39445 2497 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 39364 2497 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 39283 2497 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 39202 2497 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 39121 2497 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 39040 2497 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 38959 2497 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 38879 2497 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 38799 2497 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 38719 2497 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 38639 2497 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 38559 2497 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 38479 2497 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 38399 2497 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 38319 2497 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 38239 2497 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 38159 2497 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 38079 2497 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 37999 2497 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 37919 2497 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 37839 2497 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 37759 2497 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 37679 2497 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 37599 2497 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 37519 2497 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 37439 2497 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 37359 2497 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 37279 2497 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 37199 2497 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 37119 2497 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 37039 2497 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 36959 2497 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 36879 2497 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 36799 2497 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 36719 2497 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 36639 2497 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 36559 2497 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 36479 2497 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 36399 2497 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 36319 2497 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 36239 2497 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 36159 2497 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 36079 2497 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 35999 2497 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 35919 2497 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 35839 2497 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 35759 2497 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 35679 2497 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 35599 2497 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 35519 2497 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 35439 2497 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 35359 2497 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 35279 2497 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2457 35199 2497 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2391 6042 2431 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2391 5956 2431 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2391 5870 2431 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2391 5784 2431 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2391 5698 2431 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2391 5612 2431 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2391 5526 2431 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2391 5440 2431 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2391 5354 2431 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2391 5268 2431 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2391 5182 2431 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 39931 2417 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 39850 2417 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 39769 2417 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 39688 2417 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 39607 2417 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 39526 2417 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 39445 2417 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 39364 2417 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 39283 2417 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 39202 2417 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 39121 2417 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 39040 2417 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 38959 2417 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 38879 2417 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 38799 2417 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 38719 2417 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 38639 2417 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 38559 2417 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 38479 2417 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 38399 2417 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 38319 2417 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 38239 2417 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 38159 2417 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 38079 2417 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 37999 2417 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 37919 2417 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 37839 2417 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 37759 2417 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 37679 2417 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 37599 2417 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 37519 2417 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 37439 2417 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 37359 2417 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 37279 2417 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 37199 2417 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 37119 2417 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 37039 2417 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 36959 2417 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 36879 2417 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 36799 2417 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 36719 2417 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 36639 2417 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 36559 2417 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 36479 2417 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 36399 2417 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 36319 2417 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 36239 2417 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 36159 2417 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 36079 2417 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 35999 2417 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 35919 2417 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 35839 2417 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 35759 2417 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 35679 2417 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 35599 2417 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 35519 2417 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 35439 2417 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 35359 2417 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 35279 2417 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2377 35199 2417 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 6042 2350 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5956 2350 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5870 2350 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5784 2350 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5698 2350 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5612 2350 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5526 2350 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5440 2350 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5354 2350 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5268 2350 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2310 5182 2350 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 39931 2337 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 39850 2337 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 39769 2337 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 39688 2337 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 39607 2337 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 39526 2337 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 39445 2337 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 39364 2337 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 39283 2337 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 39202 2337 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 39121 2337 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 39040 2337 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 38959 2337 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 38879 2337 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 38799 2337 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 38719 2337 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 38639 2337 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 38559 2337 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 38479 2337 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 38399 2337 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 38319 2337 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 38239 2337 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 38159 2337 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 38079 2337 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 37999 2337 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 37919 2337 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 37839 2337 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 37759 2337 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 37679 2337 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 37599 2337 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 37519 2337 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 37439 2337 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 37359 2337 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 37279 2337 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 37199 2337 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 37119 2337 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 37039 2337 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 36959 2337 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 36879 2337 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 36799 2337 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 36719 2337 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 36639 2337 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 36559 2337 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 36479 2337 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 36399 2337 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 36319 2337 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 36239 2337 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 36159 2337 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 36079 2337 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 35999 2337 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 35919 2337 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 35839 2337 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 35759 2337 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 35679 2337 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 35599 2337 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 35519 2337 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 35439 2337 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 35359 2337 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 35279 2337 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2297 35199 2337 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2229 6042 2269 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2229 5956 2269 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2229 5870 2269 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2229 5784 2269 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2229 5698 2269 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2229 5612 2269 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2229 5526 2269 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2229 5440 2269 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2229 5354 2269 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2229 5268 2269 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2229 5182 2269 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 39931 2257 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 39850 2257 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 39769 2257 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 39688 2257 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 39607 2257 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 39526 2257 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 39445 2257 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 39364 2257 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 39283 2257 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 39202 2257 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 39121 2257 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 39040 2257 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 38959 2257 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 38879 2257 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 38799 2257 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 38719 2257 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 38639 2257 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 38559 2257 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 38479 2257 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 38399 2257 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 38319 2257 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 38239 2257 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 38159 2257 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 38079 2257 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 37999 2257 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 37919 2257 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 37839 2257 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 37759 2257 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 37679 2257 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 37599 2257 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 37519 2257 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 37439 2257 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 37359 2257 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 37279 2257 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 37199 2257 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 37119 2257 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 37039 2257 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 36959 2257 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 36879 2257 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 36799 2257 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 36719 2257 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 36639 2257 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 36559 2257 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 36479 2257 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 36399 2257 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 36319 2257 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 36239 2257 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 36159 2257 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 36079 2257 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 35999 2257 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 35919 2257 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 35839 2257 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 35759 2257 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 35679 2257 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 35599 2257 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 35519 2257 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 35439 2257 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 35359 2257 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 35279 2257 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2217 35199 2257 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2148 6042 2188 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2148 5956 2188 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2148 5870 2188 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2148 5784 2188 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2148 5698 2188 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2148 5612 2188 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2148 5526 2188 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2148 5440 2188 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2148 5354 2188 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2148 5268 2188 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2148 5182 2188 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 39931 2177 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 39850 2177 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 39769 2177 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 39688 2177 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 39607 2177 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 39526 2177 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 39445 2177 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 39364 2177 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 39283 2177 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 39202 2177 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 39121 2177 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 39040 2177 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 38959 2177 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 38879 2177 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 38799 2177 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 38719 2177 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 38639 2177 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 38559 2177 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 38479 2177 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 38399 2177 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 38319 2177 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 38239 2177 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 38159 2177 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 38079 2177 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 37999 2177 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 37919 2177 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 37839 2177 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 37759 2177 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 37679 2177 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 37599 2177 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 37519 2177 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 37439 2177 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 37359 2177 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 37279 2177 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 37199 2177 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 37119 2177 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 37039 2177 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 36959 2177 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 36879 2177 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 36799 2177 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 36719 2177 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 36639 2177 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 36559 2177 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 36479 2177 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 36399 2177 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 36319 2177 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 36239 2177 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 36159 2177 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 36079 2177 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 35999 2177 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 35919 2177 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 35839 2177 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 35759 2177 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 35679 2177 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 35599 2177 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 35519 2177 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 35439 2177 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 35359 2177 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 35279 2177 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2137 35199 2177 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2067 6042 2107 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2067 5956 2107 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2067 5870 2107 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2067 5784 2107 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2067 5698 2107 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2067 5612 2107 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2067 5526 2107 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2067 5440 2107 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2067 5354 2107 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2067 5268 2107 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2067 5182 2107 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 39931 2097 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 39850 2097 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 39769 2097 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 39688 2097 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 39607 2097 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 39526 2097 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 39445 2097 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 39364 2097 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 39283 2097 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 39202 2097 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 39121 2097 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 39040 2097 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 38959 2097 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 38879 2097 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 38799 2097 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 38719 2097 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 38639 2097 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 38559 2097 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 38479 2097 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 38399 2097 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 38319 2097 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 38239 2097 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 38159 2097 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 38079 2097 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 37999 2097 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 37919 2097 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 37839 2097 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 37759 2097 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 37679 2097 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 37599 2097 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 37519 2097 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 37439 2097 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 37359 2097 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 37279 2097 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 37199 2097 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 37119 2097 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 37039 2097 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 36959 2097 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 36879 2097 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 36799 2097 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 36719 2097 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 36639 2097 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 36559 2097 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 36479 2097 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 36399 2097 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 36319 2097 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 36239 2097 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 36159 2097 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 36079 2097 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 35999 2097 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 35919 2097 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 35839 2097 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 35759 2097 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 35679 2097 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 35599 2097 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 35519 2097 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 35439 2097 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 35359 2097 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 35279 2097 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 2057 35199 2097 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 6042 2026 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5956 2026 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5870 2026 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5784 2026 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5698 2026 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5612 2026 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5526 2026 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5440 2026 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5354 2026 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5268 2026 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1986 5182 2026 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 39931 2017 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 39850 2017 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 39769 2017 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 39688 2017 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 39607 2017 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 39526 2017 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 39445 2017 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 39364 2017 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 39283 2017 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 39202 2017 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 39121 2017 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 39040 2017 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 38959 2017 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 38879 2017 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 38799 2017 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 38719 2017 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 38639 2017 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 38559 2017 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 38479 2017 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 38399 2017 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 38319 2017 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 38239 2017 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 38159 2017 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 38079 2017 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 37999 2017 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 37919 2017 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 37839 2017 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 37759 2017 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 37679 2017 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 37599 2017 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 37519 2017 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 37439 2017 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 37359 2017 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 37279 2017 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 37199 2017 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 37119 2017 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 37039 2017 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 36959 2017 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 36879 2017 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 36799 2017 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 36719 2017 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 36639 2017 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 36559 2017 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 36479 2017 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 36399 2017 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 36319 2017 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 36239 2017 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 36159 2017 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 36079 2017 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 35999 2017 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 35919 2017 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 35839 2017 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 35759 2017 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 35679 2017 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 35599 2017 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 35519 2017 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 35439 2017 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 35359 2017 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 35279 2017 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1977 35199 2017 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1905 6042 1945 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1905 5956 1945 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1905 5870 1945 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1905 5784 1945 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1905 5698 1945 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1905 5612 1945 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1905 5526 1945 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1905 5440 1945 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1905 5354 1945 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1905 5268 1945 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1905 5182 1945 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 39931 1937 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 39850 1937 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 39769 1937 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 39688 1937 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 39607 1937 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 39526 1937 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 39445 1937 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 39364 1937 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 39283 1937 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 39202 1937 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 39121 1937 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 39040 1937 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 38959 1937 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 38879 1937 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 38799 1937 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 38719 1937 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 38639 1937 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 38559 1937 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 38479 1937 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 38399 1937 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 38319 1937 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 38239 1937 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 38159 1937 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 38079 1937 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 37999 1937 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 37919 1937 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 37839 1937 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 37759 1937 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 37679 1937 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 37599 1937 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 37519 1937 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 37439 1937 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 37359 1937 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 37279 1937 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 37199 1937 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 37119 1937 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 37039 1937 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 36959 1937 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 36879 1937 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 36799 1937 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 36719 1937 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 36639 1937 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 36559 1937 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 36479 1937 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 36399 1937 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 36319 1937 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 36239 1937 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 36159 1937 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 36079 1937 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 35999 1937 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 35919 1937 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 35839 1937 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 35759 1937 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 35679 1937 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 35599 1937 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 35519 1937 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 35439 1937 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 35359 1937 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 35279 1937 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1897 35199 1937 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1824 6042 1864 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1824 5956 1864 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1824 5870 1864 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1824 5784 1864 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1824 5698 1864 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1824 5612 1864 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1824 5526 1864 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1824 5440 1864 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1824 5354 1864 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1824 5268 1864 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1824 5182 1864 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 39931 1857 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 39850 1857 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 39769 1857 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 39688 1857 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 39607 1857 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 39526 1857 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 39445 1857 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 39364 1857 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 39283 1857 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 39202 1857 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 39121 1857 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 39040 1857 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 38959 1857 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 38879 1857 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 38799 1857 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 38719 1857 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 38639 1857 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 38559 1857 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 38479 1857 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 38399 1857 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 38319 1857 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 38239 1857 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 38159 1857 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 38079 1857 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 37999 1857 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 37919 1857 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 37839 1857 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 37759 1857 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 37679 1857 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 37599 1857 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 37519 1857 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 37439 1857 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 37359 1857 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 37279 1857 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 37199 1857 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 37119 1857 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 37039 1857 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 36959 1857 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 36879 1857 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 36799 1857 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 36719 1857 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 36639 1857 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 36559 1857 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 36479 1857 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 36399 1857 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 36319 1857 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 36239 1857 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 36159 1857 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 36079 1857 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 35999 1857 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 35919 1857 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 35839 1857 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 35759 1857 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 35679 1857 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 35599 1857 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 35519 1857 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 35439 1857 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 35359 1857 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 35279 1857 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1817 35199 1857 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1743 6042 1783 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1743 5956 1783 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1743 5870 1783 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1743 5784 1783 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1743 5698 1783 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1743 5612 1783 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1743 5526 1783 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1743 5440 1783 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1743 5354 1783 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1743 5268 1783 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1743 5182 1783 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 39931 1777 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 39850 1777 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 39769 1777 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 39688 1777 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 39607 1777 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 39526 1777 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 39445 1777 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 39364 1777 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 39283 1777 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 39202 1777 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 39121 1777 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 39040 1777 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 38959 1777 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 38879 1777 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 38799 1777 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 38719 1777 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 38639 1777 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 38559 1777 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 38479 1777 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 38399 1777 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 38319 1777 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 38239 1777 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 38159 1777 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 38079 1777 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 37999 1777 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 37919 1777 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 37839 1777 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 37759 1777 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 37679 1777 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 37599 1777 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 37519 1777 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 37439 1777 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 37359 1777 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 37279 1777 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 37199 1777 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 37119 1777 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 37039 1777 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 36959 1777 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 36879 1777 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 36799 1777 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 36719 1777 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 36639 1777 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 36559 1777 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 36479 1777 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 36399 1777 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 36319 1777 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 36239 1777 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 36159 1777 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 36079 1777 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 35999 1777 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 35919 1777 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 35839 1777 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 35759 1777 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 35679 1777 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 35599 1777 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 35519 1777 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 35439 1777 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 35359 1777 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 35279 1777 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1737 35199 1777 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 6042 1702 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5956 1702 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5870 1702 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5784 1702 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5698 1702 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5612 1702 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5526 1702 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5440 1702 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5354 1702 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5268 1702 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1662 5182 1702 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 39931 1697 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 39850 1697 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 39769 1697 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 39688 1697 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 39607 1697 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 39526 1697 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 39445 1697 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 39364 1697 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 39283 1697 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 39202 1697 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 39121 1697 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 39040 1697 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 38959 1697 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 38879 1697 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 38799 1697 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 38719 1697 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 38639 1697 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 38559 1697 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 38479 1697 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 38399 1697 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 38319 1697 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 38239 1697 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 38159 1697 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 38079 1697 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 37999 1697 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 37919 1697 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 37839 1697 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 37759 1697 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 37679 1697 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 37599 1697 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 37519 1697 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 37439 1697 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 37359 1697 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 37279 1697 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 37199 1697 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 37119 1697 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 37039 1697 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 36959 1697 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 36879 1697 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 36799 1697 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 36719 1697 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 36639 1697 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 36559 1697 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 36479 1697 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 36399 1697 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 36319 1697 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 36239 1697 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 36159 1697 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 36079 1697 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 35999 1697 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 35919 1697 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 35839 1697 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 35759 1697 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 35679 1697 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 35599 1697 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 35519 1697 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 35439 1697 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 35359 1697 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 35279 1697 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1657 35199 1697 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1581 6042 1621 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1581 5956 1621 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1581 5870 1621 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1581 5784 1621 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1581 5698 1621 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1581 5612 1621 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1581 5526 1621 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1581 5440 1621 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1581 5354 1621 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1581 5268 1621 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1581 5182 1621 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 39931 1617 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 39850 1617 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 39769 1617 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 39688 1617 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 39607 1617 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 39526 1617 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 39445 1617 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 39364 1617 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 39283 1617 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 39202 1617 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 39121 1617 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 39040 1617 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 38959 1617 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 38879 1617 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 38799 1617 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 38719 1617 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 38639 1617 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 38559 1617 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 38479 1617 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 38399 1617 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 38319 1617 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 38239 1617 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 38159 1617 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 38079 1617 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 37999 1617 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 37919 1617 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 37839 1617 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 37759 1617 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 37679 1617 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 37599 1617 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 37519 1617 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 37439 1617 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 37359 1617 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 37279 1617 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 37199 1617 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 37119 1617 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 37039 1617 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 36959 1617 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 36879 1617 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 36799 1617 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 36719 1617 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 36639 1617 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 36559 1617 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 36479 1617 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 36399 1617 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 36319 1617 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 36239 1617 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 36159 1617 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 36079 1617 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 35999 1617 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 35919 1617 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 35839 1617 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 35759 1617 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 35679 1617 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 35599 1617 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 35519 1617 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 35439 1617 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 35359 1617 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 35279 1617 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1577 35199 1617 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1500 6042 1540 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1500 5956 1540 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1500 5870 1540 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1500 5784 1540 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1500 5698 1540 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1500 5612 1540 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1500 5526 1540 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1500 5440 1540 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1500 5354 1540 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1500 5268 1540 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1500 5182 1540 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 39931 1537 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 39850 1537 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 39769 1537 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 39688 1537 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 39607 1537 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 39526 1537 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 39445 1537 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 39364 1537 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 39283 1537 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 39202 1537 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 39121 1537 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 39040 1537 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 38959 1537 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 38879 1537 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 38799 1537 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 38719 1537 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 38639 1537 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 38559 1537 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 38479 1537 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 38399 1537 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 38319 1537 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 38239 1537 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 38159 1537 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 38079 1537 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 37999 1537 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 37919 1537 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 37839 1537 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 37759 1537 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 37679 1537 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 37599 1537 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 37519 1537 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 37439 1537 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 37359 1537 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 37279 1537 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 37199 1537 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 37119 1537 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 37039 1537 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 36959 1537 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 36879 1537 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 36799 1537 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 36719 1537 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 36639 1537 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 36559 1537 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 36479 1537 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 36399 1537 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 36319 1537 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 36239 1537 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 36159 1537 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 36079 1537 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 35999 1537 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 35919 1537 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 35839 1537 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 35759 1537 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 35679 1537 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 35599 1537 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 35519 1537 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 35439 1537 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 35359 1537 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 35279 1537 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1497 35199 1537 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1419 6042 1459 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1419 5956 1459 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1419 5870 1459 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1419 5784 1459 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1419 5698 1459 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1419 5612 1459 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1419 5526 1459 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1419 5440 1459 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1419 5354 1459 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1419 5268 1459 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1419 5182 1459 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 39931 1457 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 39850 1457 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 39769 1457 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 39688 1457 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 39607 1457 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 39526 1457 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 39445 1457 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 39364 1457 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 39283 1457 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 39202 1457 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 39121 1457 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 39040 1457 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 38959 1457 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 38879 1457 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 38799 1457 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 38719 1457 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 38639 1457 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 38559 1457 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 38479 1457 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 38399 1457 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 38319 1457 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 38239 1457 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 38159 1457 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 38079 1457 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 37999 1457 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 37919 1457 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 37839 1457 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 37759 1457 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 37679 1457 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 37599 1457 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 37519 1457 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 37439 1457 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 37359 1457 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 37279 1457 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 37199 1457 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 37119 1457 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 37039 1457 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 36959 1457 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 36879 1457 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 36799 1457 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 36719 1457 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 36639 1457 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 36559 1457 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 36479 1457 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 36399 1457 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 36319 1457 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 36239 1457 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 36159 1457 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 36079 1457 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 35999 1457 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 35919 1457 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 35839 1457 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 35759 1457 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 35679 1457 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 35599 1457 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 35519 1457 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 35439 1457 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 35359 1457 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 35279 1457 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1417 35199 1457 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 6042 1378 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5956 1378 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5870 1378 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5784 1378 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5698 1378 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5612 1378 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5526 1378 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5440 1378 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5354 1378 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5268 1378 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1338 5182 1378 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 39931 1377 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 39850 1377 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 39769 1377 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 39688 1377 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 39607 1377 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 39526 1377 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 39445 1377 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 39364 1377 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 39283 1377 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 39202 1377 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 39121 1377 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 39040 1377 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 38959 1377 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 38879 1377 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 38799 1377 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 38719 1377 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 38639 1377 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 38559 1377 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 38479 1377 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 38399 1377 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 38319 1377 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 38239 1377 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 38159 1377 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 38079 1377 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 37999 1377 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 37919 1377 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 37839 1377 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 37759 1377 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 37679 1377 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 37599 1377 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 37519 1377 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 37439 1377 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 37359 1377 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 37279 1377 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 37199 1377 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 37119 1377 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 37039 1377 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 36959 1377 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 36879 1377 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 36799 1377 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 36719 1377 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 36639 1377 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 36559 1377 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 36479 1377 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 36399 1377 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 36319 1377 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 36239 1377 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 36159 1377 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 36079 1377 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 35999 1377 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 35919 1377 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 35839 1377 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 35759 1377 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 35679 1377 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 35599 1377 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 35519 1377 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 35439 1377 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 35359 1377 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 35279 1377 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1337 35199 1377 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 39931 1297 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 39850 1297 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 39769 1297 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 39688 1297 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 39607 1297 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 39526 1297 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 39445 1297 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 39364 1297 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 39283 1297 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 39202 1297 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 39121 1297 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 39040 1297 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 38959 1297 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 38879 1297 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 38799 1297 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 38719 1297 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 38639 1297 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 38559 1297 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 38479 1297 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 38399 1297 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 38319 1297 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 38239 1297 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 38159 1297 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 38079 1297 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 37999 1297 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 37919 1297 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 37839 1297 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 37759 1297 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 37679 1297 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 37599 1297 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 37519 1297 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 37439 1297 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 37359 1297 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 37279 1297 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 37199 1297 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 37119 1297 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 37039 1297 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 36959 1297 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 36879 1297 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 36799 1297 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 36719 1297 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 36639 1297 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 36559 1297 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 36479 1297 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 36399 1297 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 36319 1297 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 36239 1297 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 36159 1297 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 36079 1297 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 35999 1297 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 35919 1297 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 35839 1297 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 35759 1297 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 35679 1297 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 35599 1297 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 35519 1297 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 35439 1297 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 35359 1297 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 35279 1297 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 35199 1297 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 6042 1297 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 5956 1297 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 5870 1297 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 5784 1297 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 5698 1297 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 5612 1297 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 5526 1297 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 5440 1297 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 5354 1297 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 5268 1297 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1257 5182 1297 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 39931 1217 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 39850 1217 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 39769 1217 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 39688 1217 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 39607 1217 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 39526 1217 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 39445 1217 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 39364 1217 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 39283 1217 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 39202 1217 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 39121 1217 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 39040 1217 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 38959 1217 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 38879 1217 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 38799 1217 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 38719 1217 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 38639 1217 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 38559 1217 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 38479 1217 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 38399 1217 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 38319 1217 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 38239 1217 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 38159 1217 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 38079 1217 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 37999 1217 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 37919 1217 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 37839 1217 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 37759 1217 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 37679 1217 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 37599 1217 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 37519 1217 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 37439 1217 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 37359 1217 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 37279 1217 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 37199 1217 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 37119 1217 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 37039 1217 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 36959 1217 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 36879 1217 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 36799 1217 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 36719 1217 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 36639 1217 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 36559 1217 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 36479 1217 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 36399 1217 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 36319 1217 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 36239 1217 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 36159 1217 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 36079 1217 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 35999 1217 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 35919 1217 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 35839 1217 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 35759 1217 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 35679 1217 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 35599 1217 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 35519 1217 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 35439 1217 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 35359 1217 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 35279 1217 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1177 35199 1217 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1176 6042 1216 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1176 5956 1216 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1176 5870 1216 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1176 5784 1216 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1176 5698 1216 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1176 5612 1216 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1176 5526 1216 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1176 5440 1216 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1176 5354 1216 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1176 5268 1216 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1176 5182 1216 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 39931 1137 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 39850 1137 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 39769 1137 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 39688 1137 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 39607 1137 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 39526 1137 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 39445 1137 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 39364 1137 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 39283 1137 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 39202 1137 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 39121 1137 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 39040 1137 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 38959 1137 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 38879 1137 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 38799 1137 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 38719 1137 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 38639 1137 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 38559 1137 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 38479 1137 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 38399 1137 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 38319 1137 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 38239 1137 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 38159 1137 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 38079 1137 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 37999 1137 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 37919 1137 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 37839 1137 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 37759 1137 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 37679 1137 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 37599 1137 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 37519 1137 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 37439 1137 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 37359 1137 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 37279 1137 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 37199 1137 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 37119 1137 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 37039 1137 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 36959 1137 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 36879 1137 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 36799 1137 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 36719 1137 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 36639 1137 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 36559 1137 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 36479 1137 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 36399 1137 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 36319 1137 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 36239 1137 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 36159 1137 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 36079 1137 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 35999 1137 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 35919 1137 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 35839 1137 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 35759 1137 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 35679 1137 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 35599 1137 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 35519 1137 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 35439 1137 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 35359 1137 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 35279 1137 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1097 35199 1137 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1095 6042 1135 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1095 5956 1135 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1095 5870 1135 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1095 5784 1135 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1095 5698 1135 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1095 5612 1135 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1095 5526 1135 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1095 5440 1135 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1095 5354 1135 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1095 5268 1135 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1095 5182 1135 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 39931 1057 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 39850 1057 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 39769 1057 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 39688 1057 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 39607 1057 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 39526 1057 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 39445 1057 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 39364 1057 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 39283 1057 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 39202 1057 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 39121 1057 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 39040 1057 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 38959 1057 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 38879 1057 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 38799 1057 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 38719 1057 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 38639 1057 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 38559 1057 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 38479 1057 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 38399 1057 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 38319 1057 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 38239 1057 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 38159 1057 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 38079 1057 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 37999 1057 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 37919 1057 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 37839 1057 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 37759 1057 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 37679 1057 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 37599 1057 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 37519 1057 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 37439 1057 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 37359 1057 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 37279 1057 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 37199 1057 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 37119 1057 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 37039 1057 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 36959 1057 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 36879 1057 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 36799 1057 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 36719 1057 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 36639 1057 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 36559 1057 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 36479 1057 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 36399 1057 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 36319 1057 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 36239 1057 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 36159 1057 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 36079 1057 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 35999 1057 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 35919 1057 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 35839 1057 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 35759 1057 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 35679 1057 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 35599 1057 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 35519 1057 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 35439 1057 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 35359 1057 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 35279 1057 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1017 35199 1057 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 6042 1054 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5956 1054 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5870 1054 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5784 1054 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5698 1054 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5612 1054 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5526 1054 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5440 1054 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5354 1054 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5268 1054 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 1014 5182 1054 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 39931 977 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 39850 977 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 39769 977 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 39688 977 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 39607 977 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 39526 977 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 39445 977 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 39364 977 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 39283 977 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 39202 977 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 39121 977 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 39040 977 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 38959 977 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 38879 977 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 38799 977 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 38719 977 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 38639 977 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 38559 977 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 38479 977 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 38399 977 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 38319 977 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 38239 977 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 38159 977 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 38079 977 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 37999 977 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 37919 977 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 37839 977 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 37759 977 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 37679 977 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 37599 977 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 37519 977 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 37439 977 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 37359 977 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 37279 977 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 37199 977 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 37119 977 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 37039 977 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 36959 977 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 36879 977 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 36799 977 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 36719 977 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 36639 977 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 36559 977 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 36479 977 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 36399 977 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 36319 977 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 36239 977 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 36159 977 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 36079 977 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 35999 977 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 35919 977 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 35839 977 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 35759 977 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 35679 977 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 35599 977 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 35519 977 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 35439 977 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 35359 977 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 35279 977 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 937 35199 977 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 933 6042 973 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 933 5956 973 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 933 5870 973 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 933 5784 973 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 933 5698 973 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 933 5612 973 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 933 5526 973 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 933 5440 973 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 933 5354 973 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 933 5268 973 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 933 5182 973 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 39931 897 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 39850 897 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 39769 897 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 39688 897 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 39607 897 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 39526 897 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 39445 897 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 39364 897 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 39283 897 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 39202 897 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 39121 897 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 39040 897 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 38959 897 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 38879 897 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 38799 897 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 38719 897 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 38639 897 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 38559 897 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 38479 897 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 38399 897 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 38319 897 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 38239 897 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 38159 897 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 38079 897 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 37999 897 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 37919 897 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 37839 897 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 37759 897 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 37679 897 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 37599 897 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 37519 897 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 37439 897 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 37359 897 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 37279 897 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 37199 897 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 37119 897 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 37039 897 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 36959 897 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 36879 897 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 36799 897 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 36719 897 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 36639 897 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 36559 897 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 36479 897 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 36399 897 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 36319 897 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 36239 897 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 36159 897 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 36079 897 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 35999 897 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 35919 897 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 35839 897 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 35759 897 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 35679 897 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 35599 897 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 35519 897 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 35439 897 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 35359 897 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 35279 897 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 857 35199 897 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 852 6042 892 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 852 5956 892 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 852 5870 892 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 852 5784 892 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 852 5698 892 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 852 5612 892 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 852 5526 892 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 852 5440 892 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 852 5354 892 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 852 5268 892 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 852 5182 892 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 39931 817 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 39850 817 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 39769 817 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 39688 817 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 39607 817 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 39526 817 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 39445 817 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 39364 817 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 39283 817 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 39202 817 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 39121 817 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 39040 817 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 38959 817 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 38879 817 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 38799 817 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 38719 817 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 38639 817 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 38559 817 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 38479 817 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 38399 817 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 38319 817 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 38239 817 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 38159 817 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 38079 817 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 37999 817 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 37919 817 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 37839 817 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 37759 817 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 37679 817 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 37599 817 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 37519 817 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 37439 817 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 37359 817 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 37279 817 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 37199 817 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 37119 817 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 37039 817 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 36959 817 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 36879 817 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 36799 817 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 36719 817 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 36639 817 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 36559 817 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 36479 817 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 36399 817 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 36319 817 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 36239 817 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 36159 817 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 36079 817 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 35999 817 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 35919 817 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 35839 817 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 35759 817 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 35679 817 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 35599 817 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 35519 817 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 35439 817 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 35359 817 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 35279 817 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 777 35199 817 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 771 6042 811 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 771 5956 811 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 771 5870 811 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 771 5784 811 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 771 5698 811 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 771 5612 811 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 771 5526 811 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 771 5440 811 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 771 5354 811 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 771 5268 811 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 771 5182 811 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 39931 737 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 39850 737 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 39769 737 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 39688 737 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 39607 737 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 39526 737 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 39445 737 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 39364 737 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 39283 737 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 39202 737 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 39121 737 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 39040 737 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 38959 737 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 38879 737 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 38799 737 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 38719 737 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 38639 737 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 38559 737 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 38479 737 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 38399 737 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 38319 737 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 38239 737 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 38159 737 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 38079 737 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 37999 737 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 37919 737 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 37839 737 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 37759 737 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 37679 737 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 37599 737 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 37519 737 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 37439 737 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 37359 737 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 37279 737 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 37199 737 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 37119 737 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 37039 737 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 36959 737 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 36879 737 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 36799 737 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 36719 737 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 36639 737 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 36559 737 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 36479 737 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 36399 737 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 36319 737 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 36239 737 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 36159 737 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 36079 737 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 35999 737 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 35919 737 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 35839 737 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 35759 737 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 35679 737 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 35599 737 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 35519 737 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 35439 737 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 35359 737 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 35279 737 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 697 35199 737 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 6042 730 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5956 730 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5870 730 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5784 730 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5698 730 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5612 730 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5526 730 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5440 730 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5354 730 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5268 730 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 690 5182 730 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 39931 657 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 39850 657 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 39769 657 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 39688 657 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 39607 657 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 39526 657 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 39445 657 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 39364 657 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 39283 657 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 39202 657 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 39121 657 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 39040 657 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 38959 657 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 38879 657 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 38799 657 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 38719 657 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 38639 657 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 38559 657 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 38479 657 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 38399 657 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 38319 657 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 38239 657 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 38159 657 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 38079 657 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 37999 657 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 37919 657 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 37839 657 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 37759 657 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 37679 657 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 37599 657 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 37519 657 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 37439 657 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 37359 657 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 37279 657 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 37199 657 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 37119 657 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 37039 657 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 36959 657 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 36879 657 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 36799 657 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 36719 657 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 36639 657 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 36559 657 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 36479 657 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 36399 657 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 36319 657 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 36239 657 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 36159 657 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 36079 657 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 35999 657 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 35919 657 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 35839 657 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 35759 657 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 35679 657 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 35599 657 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 35519 657 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 35439 657 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 35359 657 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 35279 657 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 617 35199 657 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 609 6042 649 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 609 5956 649 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 609 5870 649 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 609 5784 649 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 609 5698 649 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 609 5612 649 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 609 5526 649 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 609 5440 649 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 609 5354 649 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 609 5268 649 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 609 5182 649 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 39931 577 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 39850 577 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 39769 577 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 39688 577 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 39607 577 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 39526 577 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 39445 577 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 39364 577 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 39283 577 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 39202 577 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 39121 577 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 39040 577 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 38959 577 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 38879 577 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 38799 577 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 38719 577 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 38639 577 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 38559 577 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 38479 577 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 38399 577 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 38319 577 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 38239 577 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 38159 577 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 38079 577 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 37999 577 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 37919 577 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 37839 577 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 37759 577 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 37679 577 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 37599 577 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 37519 577 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 37439 577 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 37359 577 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 37279 577 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 37199 577 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 37119 577 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 37039 577 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 36959 577 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 36879 577 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 36799 577 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 36719 577 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 36639 577 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 36559 577 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 36479 577 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 36399 577 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 36319 577 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 36239 577 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 36159 577 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 36079 577 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 35999 577 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 35919 577 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 35839 577 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 35759 577 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 35679 577 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 35599 577 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 35519 577 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 35439 577 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 35359 577 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 35279 577 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 537 35199 577 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 527 6042 567 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 527 5956 567 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 527 5870 567 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 527 5784 567 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 527 5698 567 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 527 5612 567 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 527 5526 567 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 527 5440 567 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 527 5354 567 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 527 5268 567 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 527 5182 567 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 39931 497 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 39850 497 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 39769 497 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 39688 497 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 39607 497 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 39526 497 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 39445 497 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 39364 497 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 39283 497 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 39202 497 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 39121 497 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 39040 497 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 38959 497 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 38879 497 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 38799 497 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 38719 497 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 38639 497 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 38559 497 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 38479 497 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 38399 497 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 38319 497 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 38239 497 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 38159 497 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 38079 497 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 37999 497 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 37919 497 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 37839 497 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 37759 497 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 37679 497 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 37599 497 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 37519 497 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 37439 497 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 37359 497 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 37279 497 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 37199 497 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 37119 497 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 37039 497 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 36959 497 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 36879 497 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 36799 497 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 36719 497 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 36639 497 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 36559 497 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 36479 497 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 36399 497 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 36319 497 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 36239 497 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 36159 497 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 36079 497 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 35999 497 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 35919 497 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 35839 497 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 35759 497 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 35679 497 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 35599 497 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 35519 497 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 35439 497 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 35359 497 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 35279 497 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 457 35199 497 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 6042 485 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 5956 485 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 5870 485 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 5784 485 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 5698 485 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 5612 485 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 5526 485 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 5440 485 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 5354 485 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 5268 485 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 445 5182 485 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 39931 417 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 39850 417 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 39769 417 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 39688 417 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 39607 417 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 39526 417 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 39445 417 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 39364 417 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 39283 417 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 39202 417 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 39121 417 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 39040 417 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 38959 417 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 38879 417 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 38799 417 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 38719 417 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 38639 417 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 38559 417 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 38479 417 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 38399 417 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 38319 417 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 38239 417 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 38159 417 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 38079 417 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 37999 417 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 37919 417 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 37839 417 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 37759 417 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 37679 417 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 37599 417 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 37519 417 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 37439 417 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 37359 417 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 37279 417 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 37199 417 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 37119 417 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 37039 417 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 36959 417 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 36879 417 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 36799 417 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 36719 417 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 36639 417 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 36559 417 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 36479 417 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 36399 417 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 36319 417 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 36239 417 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 36159 417 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 36079 417 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 35999 417 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 35919 417 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 35839 417 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 35759 417 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 35679 417 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 35599 417 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 35519 417 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 35439 417 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 35359 417 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 35279 417 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 377 35199 417 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 6042 403 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5956 403 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5870 403 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5784 403 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5698 403 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5612 403 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5526 403 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5440 403 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5354 403 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5268 403 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 363 5182 403 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 39931 337 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 39850 337 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 39769 337 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 39688 337 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 39607 337 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 39526 337 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 39445 337 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 39364 337 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 39283 337 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 39202 337 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 39121 337 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 39040 337 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 38959 337 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 38879 337 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 38799 337 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 38719 337 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 38639 337 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 38559 337 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 38479 337 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 38399 337 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 38319 337 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 38239 337 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 38159 337 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 38079 337 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 37999 337 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 37919 337 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 37839 337 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 37759 337 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 37679 337 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 37599 337 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 37519 337 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 37439 337 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 37359 337 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 37279 337 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 37199 337 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 37119 337 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 37039 337 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 36959 337 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 36879 337 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 36799 337 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 36719 337 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 36639 337 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 36559 337 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 36479 337 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 36399 337 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 36319 337 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 36239 337 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 36159 337 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 36079 337 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 35999 337 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 35919 337 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 35839 337 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 35759 337 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 35679 337 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 35599 337 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 35519 337 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 35439 337 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 35359 337 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 35279 337 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 297 35199 337 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 281 6042 321 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 281 5956 321 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 281 5870 321 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 281 5784 321 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 281 5698 321 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 281 5612 321 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 281 5526 321 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 281 5440 321 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 281 5354 321 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 281 5268 321 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 281 5182 321 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 39931 257 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 39850 257 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 39769 257 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 39688 257 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 39607 257 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 39526 257 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 39445 257 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 39364 257 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 39283 257 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 39202 257 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 39121 257 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 39040 257 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 38959 257 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 38879 257 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 38799 257 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 38719 257 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 38639 257 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 38559 257 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 38479 257 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 38399 257 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 38319 257 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 38239 257 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 38159 257 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 38079 257 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 37999 257 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 37919 257 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 37839 257 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 37759 257 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 37679 257 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 37599 257 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 37519 257 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 37439 257 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 37359 257 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 37279 257 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 37199 257 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 37119 257 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 37039 257 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 36959 257 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 36879 257 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 36799 257 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 36719 257 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 36639 257 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 36559 257 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 36479 257 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 36399 257 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 36319 257 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 36239 257 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 36159 257 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 36079 257 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 35999 257 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 35919 257 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 35839 257 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 35759 257 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 35679 257 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 35599 257 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 35519 257 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 35439 257 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 35359 257 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 35279 257 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 217 35199 257 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 6042 239 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5956 239 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5870 239 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5784 239 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5698 239 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5612 239 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5526 239 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5440 239 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5354 239 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5268 239 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 199 5182 239 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 39931 177 39971 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 39850 177 39890 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 39769 177 39809 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 39688 177 39728 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 39607 177 39647 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 39526 177 39566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 39445 177 39485 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 39364 177 39404 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 39283 177 39323 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 39202 177 39242 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 39121 177 39161 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 39040 177 39080 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 38959 177 38999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 38879 177 38919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 38799 177 38839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 38719 177 38759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 38639 177 38679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 38559 177 38599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 38479 177 38519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 38399 177 38439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 38319 177 38359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 38239 177 38279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 38159 177 38199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 38079 177 38119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 37999 177 38039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 37919 177 37959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 37839 177 37879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 37759 177 37799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 37679 177 37719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 37599 177 37639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 37519 177 37559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 37439 177 37479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 37359 177 37399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 37279 177 37319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 37199 177 37239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 37119 177 37159 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 37039 177 37079 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 36959 177 36999 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 36879 177 36919 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 36799 177 36839 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 36719 177 36759 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 36639 177 36679 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 36559 177 36599 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 36479 177 36519 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 36399 177 36439 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 36319 177 36359 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 36239 177 36279 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 36159 177 36199 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 36079 177 36119 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 35999 177 36039 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 35919 177 35959 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 35839 177 35879 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 35759 177 35799 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 35679 177 35719 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 35599 177 35639 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 35519 177 35559 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 35439 177 35479 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 35359 177 35399 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 35279 177 35319 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 137 35199 177 35239 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 6042 157 6082 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5956 157 5996 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5870 157 5910 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5784 157 5824 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5698 157 5738 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5612 157 5652 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5526 157 5566 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5440 157 5480 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5354 157 5394 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5268 157 5308 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal3 s 117 5182 157 5222 6 VSSIO
port 5 nsew ground bidirectional
rlabel metal5 s 0 6397 254 7047 6 VSWITCH
port 6 nsew power bidirectional
rlabel metal5 s 14746 6397 15000 7047 6 VSWITCH
port 6 nsew power bidirectional
rlabel metal4 s 0 6377 254 7067 6 VSWITCH
port 6 nsew power bidirectional
rlabel metal4 s 14746 6377 15000 7067 6 VSWITCH
port 6 nsew power bidirectional
rlabel metal4 s 14746 6377 15000 7067 6 VSWITCH
port 6 nsew power bidirectional
rlabel metal5 s 0 6397 254 7047 6 VSWITCH
port 6 nsew power bidirectional
rlabel metal5 s 14746 6397 15000 7047 6 VSWITCH
port 6 nsew power bidirectional
rlabel metal4 s 14746 6377 15000 7067 6 VSWITCH
port 6 nsew power bidirectional
rlabel metal5 s 0 6397 254 7047 6 VSWITCH
port 6 nsew power bidirectional
rlabel metal5 s 14746 6397 15000 7047 6 VSWITCH
port 6 nsew power bidirectional
rlabel metal5 s 0 11667 254 12517 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal5 s 14746 11667 15000 12517 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 0 11647 254 12537 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 14746 11647 15000 12537 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10078 11648 14858 12536 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 0 11647 4874 12537 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10083 11647 15000 12537 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal5 s 0 11667 254 12517 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal5 s 14746 11667 15000 12517 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14800 12482 14840 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14800 12400 14840 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14800 12318 14840 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14800 12236 14840 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14800 12154 14840 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14800 12072 14840 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14800 11990 14840 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14800 11908 14840 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14800 11826 14840 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14800 11744 14840 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14800 11662 14840 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14719 12482 14759 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14719 12400 14759 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14719 12318 14759 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14719 12236 14759 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14719 12154 14759 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14719 12072 14759 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14719 11990 14759 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14719 11908 14759 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14719 11826 14759 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14719 11744 14759 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14719 11662 14759 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14638 12482 14678 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14638 12400 14678 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14638 12318 14678 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14638 12236 14678 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14638 12154 14678 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14638 12072 14678 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14638 11990 14678 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14638 11908 14678 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14638 11826 14678 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14638 11744 14678 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14638 11662 14678 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14557 12482 14597 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14557 12400 14597 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14557 12318 14597 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14557 12236 14597 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14557 12154 14597 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14557 12072 14597 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14557 11990 14597 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14557 11908 14597 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14557 11826 14597 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14557 11744 14597 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14557 11662 14597 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14476 12482 14516 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14476 12400 14516 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14476 12318 14516 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14476 12236 14516 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14476 12154 14516 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14476 12072 14516 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14476 11990 14516 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14476 11908 14516 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14476 11826 14516 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14476 11744 14516 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14476 11662 14516 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14395 12482 14435 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14395 12400 14435 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14395 12318 14435 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14395 12236 14435 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14395 12154 14435 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14395 12072 14435 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14395 11990 14435 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14395 11908 14435 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14395 11826 14435 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14395 11744 14435 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14395 11662 14435 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14314 12482 14354 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14314 12400 14354 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14314 12318 14354 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14314 12236 14354 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14314 12154 14354 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14314 12072 14354 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14314 11990 14354 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14314 11908 14354 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14314 11826 14354 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14314 11744 14354 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14314 11662 14354 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14233 12482 14273 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14233 12400 14273 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14233 12318 14273 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14233 12236 14273 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14233 12154 14273 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14233 12072 14273 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14233 11990 14273 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14233 11908 14273 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14233 11826 14273 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14233 11744 14273 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14233 11662 14273 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14152 12482 14192 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14152 12400 14192 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14152 12318 14192 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14152 12236 14192 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14152 12154 14192 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14152 12072 14192 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14152 11990 14192 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14152 11908 14192 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14152 11826 14192 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14152 11744 14192 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14152 11662 14192 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14071 12482 14111 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14071 12400 14111 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14071 12318 14111 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14071 12236 14111 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14071 12154 14111 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14071 12072 14111 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14071 11990 14111 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14071 11908 14111 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14071 11826 14111 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14071 11744 14111 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14071 11662 14111 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13990 12482 14030 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13990 12400 14030 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13990 12318 14030 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13990 12236 14030 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13990 12154 14030 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13990 12072 14030 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13990 11990 14030 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13990 11908 14030 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13990 11826 14030 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13990 11744 14030 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13990 11662 14030 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13909 12482 13949 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13909 12400 13949 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13909 12318 13949 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13909 12236 13949 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13909 12154 13949 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13909 12072 13949 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13909 11990 13949 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13909 11908 13949 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13909 11826 13949 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13909 11744 13949 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13909 11662 13949 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13828 12482 13868 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13828 12400 13868 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13828 12318 13868 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13828 12236 13868 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13828 12154 13868 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13828 12072 13868 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13828 11990 13868 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13828 11908 13868 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13828 11826 13868 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13828 11744 13868 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13828 11662 13868 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13747 12482 13787 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13747 12400 13787 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13747 12318 13787 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13747 12236 13787 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13747 12154 13787 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13747 12072 13787 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13747 11990 13787 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13747 11908 13787 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13747 11826 13787 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13747 11744 13787 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13747 11662 13787 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13666 12482 13706 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13666 12400 13706 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13666 12318 13706 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13666 12236 13706 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13666 12154 13706 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13666 12072 13706 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13666 11990 13706 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13666 11908 13706 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13666 11826 13706 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13666 11744 13706 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13666 11662 13706 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13585 12482 13625 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13585 12400 13625 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13585 12318 13625 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13585 12236 13625 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13585 12154 13625 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13585 12072 13625 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13585 11990 13625 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13585 11908 13625 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13585 11826 13625 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13585 11744 13625 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13585 11662 13625 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13504 12482 13544 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13504 12400 13544 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13504 12318 13544 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13504 12236 13544 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13504 12154 13544 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13504 12072 13544 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13504 11990 13544 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13504 11908 13544 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13504 11826 13544 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13504 11744 13544 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13504 11662 13544 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13423 12482 13463 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13423 12400 13463 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13423 12318 13463 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13423 12236 13463 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13423 12154 13463 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13423 12072 13463 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13423 11990 13463 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13423 11908 13463 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13423 11826 13463 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13423 11744 13463 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13423 11662 13463 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13342 12482 13382 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13342 12400 13382 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13342 12318 13382 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13342 12236 13382 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13342 12154 13382 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13342 12072 13382 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13342 11990 13382 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13342 11908 13382 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13342 11826 13382 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13342 11744 13382 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13342 11662 13382 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13261 12482 13301 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13261 12400 13301 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13261 12318 13301 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13261 12236 13301 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13261 12154 13301 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13261 12072 13301 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13261 11990 13301 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13261 11908 13301 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13261 11826 13301 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13261 11744 13301 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13261 11662 13301 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13180 12482 13220 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13180 12400 13220 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13180 12318 13220 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13180 12236 13220 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13180 12154 13220 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13180 12072 13220 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13180 11990 13220 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13180 11908 13220 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13180 11826 13220 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13180 11744 13220 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13180 11662 13220 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13099 12482 13139 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13099 12400 13139 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13099 12318 13139 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13099 12236 13139 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13099 12154 13139 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13099 12072 13139 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13099 11990 13139 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13099 11908 13139 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13099 11826 13139 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13099 11744 13139 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13099 11662 13139 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13018 12482 13058 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13018 12400 13058 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13018 12318 13058 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13018 12236 13058 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13018 12154 13058 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13018 12072 13058 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13018 11990 13058 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13018 11908 13058 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13018 11826 13058 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13018 11744 13058 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13018 11662 13058 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12937 12482 12977 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12937 12400 12977 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12937 12318 12977 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12937 12236 12977 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12937 12154 12977 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12937 12072 12977 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12937 11990 12977 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12937 11908 12977 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12937 11826 12977 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12937 11744 12977 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12937 11662 12977 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12856 12482 12896 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12856 12400 12896 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12856 12318 12896 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12856 12236 12896 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12856 12154 12896 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12856 12072 12896 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12856 11990 12896 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12856 11908 12896 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12856 11826 12896 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12856 11744 12896 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12856 11662 12896 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12775 12482 12815 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12775 12400 12815 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12775 12318 12815 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12775 12236 12815 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12775 12154 12815 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12775 12072 12815 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12775 11990 12815 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12775 11908 12815 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12775 11826 12815 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12775 11744 12815 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12775 11662 12815 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12694 12482 12734 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12694 12400 12734 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12694 12318 12734 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12694 12236 12734 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12694 12154 12734 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12694 12072 12734 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12694 11990 12734 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12694 11908 12734 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12694 11826 12734 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12694 11744 12734 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12694 11662 12734 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12613 12482 12653 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12613 12400 12653 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12613 12318 12653 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12613 12236 12653 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12613 12154 12653 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12613 12072 12653 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12613 11990 12653 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12613 11908 12653 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12613 11826 12653 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12613 11744 12653 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12613 11662 12653 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12532 12482 12572 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12532 12400 12572 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12532 12318 12572 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12532 12236 12572 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12532 12154 12572 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12532 12072 12572 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12532 11990 12572 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12532 11908 12572 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12532 11826 12572 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12532 11744 12572 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12532 11662 12572 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12451 12482 12491 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12451 12400 12491 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12451 12318 12491 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12451 12236 12491 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12451 12154 12491 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12451 12072 12491 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12451 11990 12491 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12451 11908 12491 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12451 11826 12491 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12451 11744 12491 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12451 11662 12491 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12370 12482 12410 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12370 12400 12410 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12370 12318 12410 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12370 12236 12410 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12370 12154 12410 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12370 12072 12410 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12370 11990 12410 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12370 11908 12410 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12370 11826 12410 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12370 11744 12410 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12370 11662 12410 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12289 12482 12329 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12289 12400 12329 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12289 12318 12329 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12289 12236 12329 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12289 12154 12329 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12289 12072 12329 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12289 11990 12329 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12289 11908 12329 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12289 11826 12329 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12289 11744 12329 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12289 11662 12329 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12208 12482 12248 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12208 12400 12248 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12208 12318 12248 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12208 12236 12248 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12208 12154 12248 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12208 12072 12248 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12208 11990 12248 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12208 11908 12248 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12208 11826 12248 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12208 11744 12248 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12208 11662 12248 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12127 12482 12167 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12127 12400 12167 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12127 12318 12167 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12127 12236 12167 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12127 12154 12167 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12127 12072 12167 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12127 11990 12167 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12127 11908 12167 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12127 11826 12167 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12127 11744 12167 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12127 11662 12167 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12046 12482 12086 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12046 12400 12086 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12046 12318 12086 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12046 12236 12086 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12046 12154 12086 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12046 12072 12086 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12046 11990 12086 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12046 11908 12086 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12046 11826 12086 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12046 11744 12086 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12046 11662 12086 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11965 12482 12005 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11965 12400 12005 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11965 12318 12005 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11965 12236 12005 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11965 12154 12005 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11965 12072 12005 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11965 11990 12005 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11965 11908 12005 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11965 11826 12005 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11965 11744 12005 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11965 11662 12005 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11884 12482 11924 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11884 12400 11924 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11884 12318 11924 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11884 12236 11924 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11884 12154 11924 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11884 12072 11924 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11884 11990 11924 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11884 11908 11924 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11884 11826 11924 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11884 11744 11924 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11884 11662 11924 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11803 12482 11843 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11803 12400 11843 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11803 12318 11843 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11803 12236 11843 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11803 12154 11843 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11803 12072 11843 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11803 11990 11843 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11803 11908 11843 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11803 11826 11843 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11803 11744 11843 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11803 11662 11843 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11722 12482 11762 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11722 12400 11762 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11722 12318 11762 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11722 12236 11762 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11722 12154 11762 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11722 12072 11762 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11722 11990 11762 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11722 11908 11762 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11722 11826 11762 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11722 11744 11762 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11722 11662 11762 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11641 12482 11681 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11641 12400 11681 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11641 12318 11681 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11641 12236 11681 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11641 12154 11681 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11641 12072 11681 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11641 11990 11681 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11641 11908 11681 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11641 11826 11681 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11641 11744 11681 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11641 11662 11681 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11560 12482 11600 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11560 12400 11600 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11560 12318 11600 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11560 12236 11600 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11560 12154 11600 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11560 12072 11600 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11560 11990 11600 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11560 11908 11600 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11560 11826 11600 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11560 11744 11600 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11560 11662 11600 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11479 12482 11519 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11479 12400 11519 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11479 12318 11519 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11479 12236 11519 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11479 12154 11519 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11479 12072 11519 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11479 11990 11519 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11479 11908 11519 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11479 11826 11519 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11479 11744 11519 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11479 11662 11519 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11398 12482 11438 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11398 12400 11438 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11398 12318 11438 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11398 12236 11438 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11398 12154 11438 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11398 12072 11438 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11398 11990 11438 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11398 11908 11438 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11398 11826 11438 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11398 11744 11438 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11398 11662 11438 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11317 12482 11357 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11317 12400 11357 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11317 12318 11357 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11317 12236 11357 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11317 12154 11357 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11317 12072 11357 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11317 11990 11357 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11317 11908 11357 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11317 11826 11357 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11317 11744 11357 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11317 11662 11357 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11236 12482 11276 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11236 12400 11276 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11236 12318 11276 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11236 12236 11276 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11236 12154 11276 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11236 12072 11276 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11236 11990 11276 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11236 11908 11276 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11236 11826 11276 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11236 11744 11276 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11236 11662 11276 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11155 12482 11195 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11155 12400 11195 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11155 12318 11195 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11155 12236 11195 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11155 12154 11195 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11155 12072 11195 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11155 11990 11195 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11155 11908 11195 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11155 11826 11195 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11155 11744 11195 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11155 11662 11195 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11074 12482 11114 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11074 12400 11114 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11074 12318 11114 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11074 12236 11114 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11074 12154 11114 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11074 12072 11114 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11074 11990 11114 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11074 11908 11114 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11074 11826 11114 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11074 11744 11114 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11074 11662 11114 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10993 12482 11033 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10993 12400 11033 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10993 12318 11033 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10993 12236 11033 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10993 12154 11033 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10993 12072 11033 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10993 11990 11033 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10993 11908 11033 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10993 11826 11033 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10993 11744 11033 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10993 11662 11033 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10912 12482 10952 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10912 12400 10952 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10912 12318 10952 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10912 12236 10952 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10912 12154 10952 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10912 12072 10952 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10912 11990 10952 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10912 11908 10952 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10912 11826 10952 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10912 11744 10952 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10912 11662 10952 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10831 12482 10871 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10831 12400 10871 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10831 12318 10871 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10831 12236 10871 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10831 12154 10871 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10831 12072 10871 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10831 11990 10871 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10831 11908 10871 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10831 11826 10871 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10831 11744 10871 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10831 11662 10871 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10750 12482 10790 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10750 12400 10790 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10750 12318 10790 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10750 12236 10790 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10750 12154 10790 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10750 12072 10790 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10750 11990 10790 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10750 11908 10790 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10750 11826 10790 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10750 11744 10790 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10750 11662 10790 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10669 12482 10709 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10669 12400 10709 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10669 12318 10709 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10669 12236 10709 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10669 12154 10709 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10669 12072 10709 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10669 11990 10709 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10669 11908 10709 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10669 11826 10709 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10669 11744 10709 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10669 11662 10709 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10588 12482 10628 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10588 12400 10628 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10588 12318 10628 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10588 12236 10628 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10588 12154 10628 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10588 12072 10628 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10588 11990 10628 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10588 11908 10628 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10588 11826 10628 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10588 11744 10628 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10588 11662 10628 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10506 12482 10546 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10506 12400 10546 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10506 12318 10546 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10506 12236 10546 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10506 12154 10546 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10506 12072 10546 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10506 11990 10546 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10506 11908 10546 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10506 11826 10546 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10506 11744 10546 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10506 11662 10546 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10424 12482 10464 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10424 12400 10464 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10424 12318 10464 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10424 12236 10464 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10424 12154 10464 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10424 12072 10464 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10424 11990 10464 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10424 11908 10464 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10424 11826 10464 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10424 11744 10464 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10424 11662 10464 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10342 12482 10382 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10342 12400 10382 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10342 12318 10382 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10342 12236 10382 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10342 12154 10382 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10342 12072 10382 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10342 11990 10382 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10342 11908 10382 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10342 11826 10382 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10342 11744 10382 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10342 11662 10382 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10260 12482 10300 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10260 12400 10300 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10260 12318 10300 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10260 12236 10300 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10260 12154 10300 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10260 12072 10300 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10260 11990 10300 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10260 11908 10300 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10260 11826 10300 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10260 11744 10300 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10260 11662 10300 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10178 12482 10218 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10178 12400 10218 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10178 12318 10218 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10178 12236 10218 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10178 12154 10218 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10178 12072 10218 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10178 11990 10218 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10178 11908 10218 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10178 11826 10218 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10178 11744 10218 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10178 11662 10218 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10096 12482 10136 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10096 12400 10136 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10096 12318 10136 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10096 12236 10136 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10096 12154 10136 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10096 12072 10136 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10096 11990 10136 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10096 11908 10136 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10096 11826 10136 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10096 11744 10136 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10096 11662 10136 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4809 12470 4873 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4809 12388 4873 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4809 12306 4873 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4809 12224 4873 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4809 12142 4873 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4809 12060 4873 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4809 11978 4873 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4809 11896 4873 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4809 11814 4873 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4809 11732 4873 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4809 11650 4873 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4728 12470 4792 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4728 12388 4792 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4728 12306 4792 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4728 12224 4792 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4728 12142 4792 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4728 12060 4792 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4728 11978 4792 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4728 11896 4792 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4728 11814 4792 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4728 11732 4792 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4728 11650 4792 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4647 12470 4711 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4647 12388 4711 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4647 12306 4711 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4647 12224 4711 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4647 12142 4711 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4647 12060 4711 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4647 11978 4711 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4647 11896 4711 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4647 11814 4711 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4647 11732 4711 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4647 11650 4711 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4566 12470 4630 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4566 12388 4630 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4566 12306 4630 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4566 12224 4630 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4566 12142 4630 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4566 12060 4630 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4566 11978 4630 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4566 11896 4630 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4566 11814 4630 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4566 11732 4630 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4566 11650 4630 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4485 12470 4549 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4485 12388 4549 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4485 12306 4549 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4485 12224 4549 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4485 12142 4549 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4485 12060 4549 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4485 11978 4549 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4485 11896 4549 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4485 11814 4549 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4485 11732 4549 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4485 11650 4549 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4404 12470 4468 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4404 12388 4468 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4404 12306 4468 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4404 12224 4468 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4404 12142 4468 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4404 12060 4468 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4404 11978 4468 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4404 11896 4468 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4404 11814 4468 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4404 11732 4468 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4404 11650 4468 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4323 12470 4387 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4323 12388 4387 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4323 12306 4387 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4323 12224 4387 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4323 12142 4387 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4323 12060 4387 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4323 11978 4387 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4323 11896 4387 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4323 11814 4387 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4323 11732 4387 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4323 11650 4387 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4242 12470 4306 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4242 12388 4306 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4242 12306 4306 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4242 12224 4306 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4242 12142 4306 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4242 12060 4306 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4242 11978 4306 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4242 11896 4306 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4242 11814 4306 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4242 11732 4306 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4242 11650 4306 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4161 12470 4225 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4161 12388 4225 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4161 12306 4225 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4161 12224 4225 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4161 12142 4225 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4161 12060 4225 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4161 11978 4225 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4161 11896 4225 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4161 11814 4225 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4161 11732 4225 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4161 11650 4225 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4080 12470 4144 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4080 12388 4144 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4080 12306 4144 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4080 12224 4144 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4080 12142 4144 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4080 12060 4144 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4080 11978 4144 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4080 11896 4144 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4080 11814 4144 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4080 11732 4144 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4080 11650 4144 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3999 12470 4063 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3999 12388 4063 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3999 12306 4063 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3999 12224 4063 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3999 12142 4063 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3999 12060 4063 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3999 11978 4063 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3999 11896 4063 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3999 11814 4063 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3999 11732 4063 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3999 11650 4063 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3918 12470 3982 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3918 12388 3982 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3918 12306 3982 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3918 12224 3982 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3918 12142 3982 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3918 12060 3982 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3918 11978 3982 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3918 11896 3982 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3918 11814 3982 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3918 11732 3982 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3918 11650 3982 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3837 12470 3901 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3837 12388 3901 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3837 12306 3901 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3837 12224 3901 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3837 12142 3901 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3837 12060 3901 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3837 11978 3901 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3837 11896 3901 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3837 11814 3901 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3837 11732 3901 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3837 11650 3901 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3756 12470 3820 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3756 12388 3820 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3756 12306 3820 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3756 12224 3820 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3756 12142 3820 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3756 12060 3820 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3756 11978 3820 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3756 11896 3820 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3756 11814 3820 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3756 11732 3820 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3756 11650 3820 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3675 12470 3739 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3675 12388 3739 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3675 12306 3739 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3675 12224 3739 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3675 12142 3739 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3675 12060 3739 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3675 11978 3739 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3675 11896 3739 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3675 11814 3739 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3675 11732 3739 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3675 11650 3739 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3594 12470 3658 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3594 12388 3658 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3594 12306 3658 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3594 12224 3658 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3594 12142 3658 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3594 12060 3658 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3594 11978 3658 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3594 11896 3658 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3594 11814 3658 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3594 11732 3658 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3594 11650 3658 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3513 12470 3577 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3513 12388 3577 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3513 12306 3577 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3513 12224 3577 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3513 12142 3577 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3513 12060 3577 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3513 11978 3577 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3513 11896 3577 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3513 11814 3577 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3513 11732 3577 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3513 11650 3577 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3432 12470 3496 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3432 12388 3496 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3432 12306 3496 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3432 12224 3496 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3432 12142 3496 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3432 12060 3496 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3432 11978 3496 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3432 11896 3496 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3432 11814 3496 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3432 11732 3496 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3432 11650 3496 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3351 12470 3415 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3351 12388 3415 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3351 12306 3415 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3351 12224 3415 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3351 12142 3415 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3351 12060 3415 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3351 11978 3415 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3351 11896 3415 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3351 11814 3415 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3351 11732 3415 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3351 11650 3415 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3270 12470 3334 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3270 12388 3334 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3270 12306 3334 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3270 12224 3334 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3270 12142 3334 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3270 12060 3334 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3270 11978 3334 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3270 11896 3334 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3270 11814 3334 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3270 11732 3334 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3270 11650 3334 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3189 12470 3253 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3189 12388 3253 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3189 12306 3253 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3189 12224 3253 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3189 12142 3253 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3189 12060 3253 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3189 11978 3253 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3189 11896 3253 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3189 11814 3253 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3189 11732 3253 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3189 11650 3253 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3108 12470 3172 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3108 12388 3172 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3108 12306 3172 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3108 12224 3172 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3108 12142 3172 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3108 12060 3172 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3108 11978 3172 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3108 11896 3172 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3108 11814 3172 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3108 11732 3172 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3108 11650 3172 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3027 12470 3091 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3027 12388 3091 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3027 12306 3091 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3027 12224 3091 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3027 12142 3091 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3027 12060 3091 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3027 11978 3091 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3027 11896 3091 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3027 11814 3091 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3027 11732 3091 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3027 11650 3091 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2946 12470 3010 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2946 12388 3010 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2946 12306 3010 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2946 12224 3010 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2946 12142 3010 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2946 12060 3010 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2946 11978 3010 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2946 11896 3010 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2946 11814 3010 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2946 11732 3010 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2946 11650 3010 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2865 12470 2929 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2865 12388 2929 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2865 12306 2929 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2865 12224 2929 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2865 12142 2929 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2865 12060 2929 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2865 11978 2929 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2865 11896 2929 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2865 11814 2929 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2865 11732 2929 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2865 11650 2929 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2784 12470 2848 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2784 12388 2848 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2784 12306 2848 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2784 12224 2848 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2784 12142 2848 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2784 12060 2848 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2784 11978 2848 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2784 11896 2848 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2784 11814 2848 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2784 11732 2848 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2784 11650 2848 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2703 12470 2767 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2703 12388 2767 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2703 12306 2767 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2703 12224 2767 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2703 12142 2767 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2703 12060 2767 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2703 11978 2767 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2703 11896 2767 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2703 11814 2767 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2703 11732 2767 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2703 11650 2767 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2622 12470 2686 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2622 12388 2686 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2622 12306 2686 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2622 12224 2686 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2622 12142 2686 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2622 12060 2686 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2622 11978 2686 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2622 11896 2686 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2622 11814 2686 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2622 11732 2686 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2622 11650 2686 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2541 12470 2605 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2541 12388 2605 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2541 12306 2605 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2541 12224 2605 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2541 12142 2605 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2541 12060 2605 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2541 11978 2605 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2541 11896 2605 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2541 11814 2605 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2541 11732 2605 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2541 11650 2605 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2460 12470 2524 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2460 12388 2524 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2460 12306 2524 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2460 12224 2524 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2460 12142 2524 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2460 12060 2524 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2460 11978 2524 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2460 11896 2524 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2460 11814 2524 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2460 11732 2524 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2460 11650 2524 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2379 12470 2443 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2379 12388 2443 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2379 12306 2443 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2379 12224 2443 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2379 12142 2443 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2379 12060 2443 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2379 11978 2443 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2379 11896 2443 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2379 11814 2443 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2379 11732 2443 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2379 11650 2443 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2298 12470 2362 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2298 12388 2362 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2298 12306 2362 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2298 12224 2362 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2298 12142 2362 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2298 12060 2362 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2298 11978 2362 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2298 11896 2362 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2298 11814 2362 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2298 11732 2362 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2298 11650 2362 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2217 12470 2281 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2217 12388 2281 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2217 12306 2281 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2217 12224 2281 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2217 12142 2281 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2217 12060 2281 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2217 11978 2281 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2217 11896 2281 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2217 11814 2281 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2217 11732 2281 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2217 11650 2281 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2136 12470 2200 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2136 12388 2200 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2136 12306 2200 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2136 12224 2200 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2136 12142 2200 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2136 12060 2200 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2136 11978 2200 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2136 11896 2200 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2136 11814 2200 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2136 11732 2200 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2136 11650 2200 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2055 12470 2119 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2055 12388 2119 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2055 12306 2119 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2055 12224 2119 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2055 12142 2119 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2055 12060 2119 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2055 11978 2119 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2055 11896 2119 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2055 11814 2119 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2055 11732 2119 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2055 11650 2119 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1974 12470 2038 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1974 12388 2038 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1974 12306 2038 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1974 12224 2038 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1974 12142 2038 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1974 12060 2038 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1974 11978 2038 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1974 11896 2038 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1974 11814 2038 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1974 11732 2038 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1974 11650 2038 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1893 12470 1957 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1893 12388 1957 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1893 12306 1957 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1893 12224 1957 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1893 12142 1957 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1893 12060 1957 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1893 11978 1957 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1893 11896 1957 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1893 11814 1957 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1893 11732 1957 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1893 11650 1957 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1812 12470 1876 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1812 12388 1876 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1812 12306 1876 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1812 12224 1876 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1812 12142 1876 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1812 12060 1876 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1812 11978 1876 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1812 11896 1876 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1812 11814 1876 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1812 11732 1876 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1812 11650 1876 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1731 12470 1795 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1731 12388 1795 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1731 12306 1795 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1731 12224 1795 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1731 12142 1795 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1731 12060 1795 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1731 11978 1795 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1731 11896 1795 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1731 11814 1795 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1731 11732 1795 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1731 11650 1795 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1650 12470 1714 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1650 12388 1714 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1650 12306 1714 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1650 12224 1714 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1650 12142 1714 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1650 12060 1714 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1650 11978 1714 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1650 11896 1714 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1650 11814 1714 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1650 11732 1714 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1650 11650 1714 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1569 12470 1633 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1569 12388 1633 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1569 12306 1633 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1569 12224 1633 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1569 12142 1633 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1569 12060 1633 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1569 11978 1633 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1569 11896 1633 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1569 11814 1633 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1569 11732 1633 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1569 11650 1633 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1488 12470 1552 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1488 12388 1552 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1488 12306 1552 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1488 12224 1552 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1488 12142 1552 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1488 12060 1552 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1488 11978 1552 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1488 11896 1552 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1488 11814 1552 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1488 11732 1552 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1488 11650 1552 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1407 12470 1471 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1407 12388 1471 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1407 12306 1471 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1407 12224 1471 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1407 12142 1471 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1407 12060 1471 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1407 11978 1471 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1407 11896 1471 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1407 11814 1471 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1407 11732 1471 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1407 11650 1471 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1326 12470 1390 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1326 12388 1390 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1326 12306 1390 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1326 12224 1390 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1326 12142 1390 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1326 12060 1390 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1326 11978 1390 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1326 11896 1390 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1326 11814 1390 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1326 11732 1390 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1326 11650 1390 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1245 12470 1309 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1245 12388 1309 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1245 12306 1309 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1245 12224 1309 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1245 12142 1309 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1245 12060 1309 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1245 11978 1309 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1245 11896 1309 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1245 11814 1309 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1245 11732 1309 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1245 11650 1309 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1164 12470 1228 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1164 12388 1228 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1164 12306 1228 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1164 12224 1228 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1164 12142 1228 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1164 12060 1228 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1164 11978 1228 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1164 11896 1228 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1164 11814 1228 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1164 11732 1228 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1164 11650 1228 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1083 12470 1147 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1083 12388 1147 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1083 12306 1147 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1083 12224 1147 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1083 12142 1147 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1083 12060 1147 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1083 11978 1147 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1083 11896 1147 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1083 11814 1147 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1083 11732 1147 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1083 11650 1147 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1002 12470 1066 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1002 12388 1066 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1002 12306 1066 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1002 12224 1066 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1002 12142 1066 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1002 12060 1066 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1002 11978 1066 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1002 11896 1066 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1002 11814 1066 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1002 11732 1066 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1002 11650 1066 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 921 12470 985 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 921 12388 985 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 921 12306 985 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 921 12224 985 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 921 12142 985 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 921 12060 985 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 921 11978 985 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 921 11896 985 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 921 11814 985 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 921 11732 985 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 921 11650 985 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 840 12470 904 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 840 12388 904 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 840 12306 904 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 840 12224 904 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 840 12142 904 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 840 12060 904 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 840 11978 904 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 840 11896 904 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 840 11814 904 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 840 11732 904 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 840 11650 904 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 759 12470 823 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 759 12388 823 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 759 12306 823 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 759 12224 823 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 759 12142 823 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 759 12060 823 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 759 11978 823 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 759 11896 823 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 759 11814 823 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 759 11732 823 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 759 11650 823 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 678 12470 742 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 678 12388 742 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 678 12306 742 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 678 12224 742 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 678 12142 742 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 678 12060 742 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 678 11978 742 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 678 11896 742 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 678 11814 742 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 678 11732 742 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 678 11650 742 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 597 12470 661 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 597 12388 661 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 597 12306 661 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 597 12224 661 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 597 12142 661 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 597 12060 661 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 597 11978 661 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 597 11896 661 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 597 11814 661 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 597 11732 661 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 597 11650 661 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 515 12470 579 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 515 12388 579 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 515 12306 579 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 515 12224 579 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 515 12142 579 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 515 12060 579 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 515 11978 579 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 515 11896 579 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 515 11814 579 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 515 11732 579 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 515 11650 579 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 433 12470 497 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 433 12388 497 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 433 12306 497 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 433 12224 497 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 433 12142 497 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 433 12060 497 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 433 11978 497 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 433 11896 497 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 433 11814 497 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 433 11732 497 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 433 11650 497 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 351 12470 415 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 351 12388 415 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 351 12306 415 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 351 12224 415 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 351 12142 415 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 351 12060 415 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 351 11978 415 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 351 11896 415 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 351 11814 415 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 351 11732 415 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 351 11650 415 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 269 12470 333 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 269 12388 333 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 269 12306 333 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 269 12224 333 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 269 12142 333 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 269 12060 333 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 269 11978 333 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 269 11896 333 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 269 11814 333 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 269 11732 333 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 269 11650 333 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 187 12470 251 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 187 12388 251 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 187 12306 251 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 187 12224 251 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 187 12142 251 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 187 12060 251 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 187 11978 251 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 187 11896 251 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 187 11814 251 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 187 11732 251 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 187 11650 251 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 105 12470 169 12534 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 105 12388 169 12452 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 105 12306 169 12370 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 105 12224 169 12288 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 105 12142 169 12206 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 105 12060 169 12124 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 105 11978 169 12042 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 105 11896 169 11960 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 105 11814 169 11878 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 105 11732 169 11796 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 105 11650 169 11714 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10078 11648 14858 12536 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 0 11647 4874 12537 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal4 s 10083 11647 15000 12537 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal5 s 0 11667 254 12517 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal5 s 14746 11667 15000 12517 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14800 12482 14840 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14800 12400 14840 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14800 12318 14840 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14800 12236 14840 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14800 12154 14840 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14800 12072 14840 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14800 11990 14840 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14800 11908 14840 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14800 11826 14840 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14800 11744 14840 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14800 11662 14840 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14719 12482 14759 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14719 12400 14759 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14719 12318 14759 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14719 12236 14759 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14719 12154 14759 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14719 12072 14759 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14719 11990 14759 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14719 11908 14759 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14719 11826 14759 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14719 11744 14759 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14719 11662 14759 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14638 12482 14678 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14638 12400 14678 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14638 12318 14678 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14638 12236 14678 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14638 12154 14678 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14638 12072 14678 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14638 11990 14678 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14638 11908 14678 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14638 11826 14678 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14638 11744 14678 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14638 11662 14678 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14557 12482 14597 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14557 12400 14597 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14557 12318 14597 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14557 12236 14597 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14557 12154 14597 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14557 12072 14597 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14557 11990 14597 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14557 11908 14597 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14557 11826 14597 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14557 11744 14597 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14557 11662 14597 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14476 12482 14516 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14476 12400 14516 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14476 12318 14516 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14476 12236 14516 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14476 12154 14516 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14476 12072 14516 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14476 11990 14516 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14476 11908 14516 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14476 11826 14516 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14476 11744 14516 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14476 11662 14516 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14395 12482 14435 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14395 12400 14435 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14395 12318 14435 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14395 12236 14435 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14395 12154 14435 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14395 12072 14435 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14395 11990 14435 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14395 11908 14435 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14395 11826 14435 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14395 11744 14435 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14395 11662 14435 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14314 12482 14354 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14314 12400 14354 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14314 12318 14354 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14314 12236 14354 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14314 12154 14354 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14314 12072 14354 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14314 11990 14354 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14314 11908 14354 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14314 11826 14354 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14314 11744 14354 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14314 11662 14354 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14233 12482 14273 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14233 12400 14273 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14233 12318 14273 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14233 12236 14273 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14233 12154 14273 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14233 12072 14273 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14233 11990 14273 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14233 11908 14273 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14233 11826 14273 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14233 11744 14273 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14233 11662 14273 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14152 12482 14192 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14152 12400 14192 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14152 12318 14192 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14152 12236 14192 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14152 12154 14192 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14152 12072 14192 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14152 11990 14192 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14152 11908 14192 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14152 11826 14192 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14152 11744 14192 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14152 11662 14192 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14071 12482 14111 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14071 12400 14111 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14071 12318 14111 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14071 12236 14111 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14071 12154 14111 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14071 12072 14111 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14071 11990 14111 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14071 11908 14111 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14071 11826 14111 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14071 11744 14111 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 14071 11662 14111 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13990 12482 14030 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13990 12400 14030 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13990 12318 14030 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13990 12236 14030 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13990 12154 14030 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13990 12072 14030 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13990 11990 14030 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13990 11908 14030 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13990 11826 14030 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13990 11744 14030 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13990 11662 14030 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13909 12482 13949 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13909 12400 13949 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13909 12318 13949 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13909 12236 13949 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13909 12154 13949 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13909 12072 13949 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13909 11990 13949 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13909 11908 13949 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13909 11826 13949 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13909 11744 13949 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13909 11662 13949 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13828 12482 13868 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13828 12400 13868 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13828 12318 13868 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13828 12236 13868 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13828 12154 13868 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13828 12072 13868 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13828 11990 13868 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13828 11908 13868 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13828 11826 13868 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13828 11744 13868 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13828 11662 13868 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13747 12482 13787 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13747 12400 13787 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13747 12318 13787 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13747 12236 13787 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13747 12154 13787 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13747 12072 13787 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13747 11990 13787 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13747 11908 13787 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13747 11826 13787 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13747 11744 13787 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13747 11662 13787 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13666 12482 13706 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13666 12400 13706 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13666 12318 13706 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13666 12236 13706 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13666 12154 13706 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13666 12072 13706 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13666 11990 13706 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13666 11908 13706 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13666 11826 13706 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13666 11744 13706 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13666 11662 13706 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13585 12482 13625 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13585 12400 13625 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13585 12318 13625 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13585 12236 13625 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13585 12154 13625 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13585 12072 13625 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13585 11990 13625 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13585 11908 13625 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13585 11826 13625 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13585 11744 13625 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13585 11662 13625 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13504 12482 13544 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13504 12400 13544 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13504 12318 13544 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13504 12236 13544 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13504 12154 13544 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13504 12072 13544 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13504 11990 13544 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13504 11908 13544 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13504 11826 13544 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13504 11744 13544 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13504 11662 13544 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13423 12482 13463 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13423 12400 13463 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13423 12318 13463 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13423 12236 13463 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13423 12154 13463 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13423 12072 13463 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13423 11990 13463 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13423 11908 13463 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13423 11826 13463 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13423 11744 13463 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13423 11662 13463 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13342 12482 13382 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13342 12400 13382 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13342 12318 13382 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13342 12236 13382 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13342 12154 13382 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13342 12072 13382 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13342 11990 13382 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13342 11908 13382 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13342 11826 13382 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13342 11744 13382 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13342 11662 13382 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13261 12482 13301 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13261 12400 13301 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13261 12318 13301 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13261 12236 13301 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13261 12154 13301 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13261 12072 13301 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13261 11990 13301 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13261 11908 13301 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13261 11826 13301 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13261 11744 13301 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13261 11662 13301 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13180 12482 13220 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13180 12400 13220 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13180 12318 13220 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13180 12236 13220 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13180 12154 13220 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13180 12072 13220 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13180 11990 13220 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13180 11908 13220 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13180 11826 13220 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13180 11744 13220 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13180 11662 13220 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13099 12482 13139 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13099 12400 13139 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13099 12318 13139 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13099 12236 13139 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13099 12154 13139 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13099 12072 13139 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13099 11990 13139 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13099 11908 13139 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13099 11826 13139 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13099 11744 13139 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13099 11662 13139 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13018 12482 13058 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13018 12400 13058 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13018 12318 13058 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13018 12236 13058 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13018 12154 13058 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13018 12072 13058 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13018 11990 13058 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13018 11908 13058 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13018 11826 13058 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13018 11744 13058 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 13018 11662 13058 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12937 12482 12977 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12937 12400 12977 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12937 12318 12977 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12937 12236 12977 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12937 12154 12977 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12937 12072 12977 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12937 11990 12977 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12937 11908 12977 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12937 11826 12977 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12937 11744 12977 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12937 11662 12977 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12856 12482 12896 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12856 12400 12896 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12856 12318 12896 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12856 12236 12896 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12856 12154 12896 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12856 12072 12896 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12856 11990 12896 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12856 11908 12896 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12856 11826 12896 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12856 11744 12896 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12856 11662 12896 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12775 12482 12815 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12775 12400 12815 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12775 12318 12815 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12775 12236 12815 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12775 12154 12815 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12775 12072 12815 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12775 11990 12815 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12775 11908 12815 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12775 11826 12815 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12775 11744 12815 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12775 11662 12815 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12694 12482 12734 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12694 12400 12734 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12694 12318 12734 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12694 12236 12734 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12694 12154 12734 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12694 12072 12734 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12694 11990 12734 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12694 11908 12734 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12694 11826 12734 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12694 11744 12734 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12694 11662 12734 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12613 12482 12653 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12613 12400 12653 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12613 12318 12653 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12613 12236 12653 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12613 12154 12653 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12613 12072 12653 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12613 11990 12653 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12613 11908 12653 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12613 11826 12653 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12613 11744 12653 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12613 11662 12653 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12532 12482 12572 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12532 12400 12572 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12532 12318 12572 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12532 12236 12572 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12532 12154 12572 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12532 12072 12572 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12532 11990 12572 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12532 11908 12572 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12532 11826 12572 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12532 11744 12572 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12532 11662 12572 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12451 12482 12491 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12451 12400 12491 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12451 12318 12491 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12451 12236 12491 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12451 12154 12491 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12451 12072 12491 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12451 11990 12491 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12451 11908 12491 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12451 11826 12491 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12451 11744 12491 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12451 11662 12491 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12370 12482 12410 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12370 12400 12410 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12370 12318 12410 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12370 12236 12410 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12370 12154 12410 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12370 12072 12410 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12370 11990 12410 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12370 11908 12410 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12370 11826 12410 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12370 11744 12410 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12370 11662 12410 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12289 12482 12329 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12289 12400 12329 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12289 12318 12329 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12289 12236 12329 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12289 12154 12329 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12289 12072 12329 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12289 11990 12329 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12289 11908 12329 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12289 11826 12329 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12289 11744 12329 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12289 11662 12329 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12208 12482 12248 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12208 12400 12248 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12208 12318 12248 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12208 12236 12248 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12208 12154 12248 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12208 12072 12248 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12208 11990 12248 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12208 11908 12248 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12208 11826 12248 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12208 11744 12248 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12208 11662 12248 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12127 12482 12167 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12127 12400 12167 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12127 12318 12167 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12127 12236 12167 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12127 12154 12167 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12127 12072 12167 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12127 11990 12167 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12127 11908 12167 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12127 11826 12167 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12127 11744 12167 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12127 11662 12167 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12046 12482 12086 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12046 12400 12086 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12046 12318 12086 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12046 12236 12086 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12046 12154 12086 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12046 12072 12086 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12046 11990 12086 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12046 11908 12086 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12046 11826 12086 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12046 11744 12086 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 12046 11662 12086 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11965 12482 12005 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11965 12400 12005 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11965 12318 12005 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11965 12236 12005 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11965 12154 12005 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11965 12072 12005 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11965 11990 12005 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11965 11908 12005 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11965 11826 12005 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11965 11744 12005 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11965 11662 12005 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11884 12482 11924 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11884 12400 11924 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11884 12318 11924 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11884 12236 11924 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11884 12154 11924 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11884 12072 11924 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11884 11990 11924 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11884 11908 11924 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11884 11826 11924 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11884 11744 11924 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11884 11662 11924 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11803 12482 11843 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11803 12400 11843 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11803 12318 11843 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11803 12236 11843 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11803 12154 11843 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11803 12072 11843 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11803 11990 11843 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11803 11908 11843 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11803 11826 11843 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11803 11744 11843 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11803 11662 11843 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11722 12482 11762 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11722 12400 11762 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11722 12318 11762 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11722 12236 11762 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11722 12154 11762 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11722 12072 11762 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11722 11990 11762 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11722 11908 11762 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11722 11826 11762 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11722 11744 11762 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11722 11662 11762 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11641 12482 11681 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11641 12400 11681 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11641 12318 11681 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11641 12236 11681 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11641 12154 11681 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11641 12072 11681 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11641 11990 11681 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11641 11908 11681 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11641 11826 11681 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11641 11744 11681 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11641 11662 11681 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11560 12482 11600 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11560 12400 11600 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11560 12318 11600 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11560 12236 11600 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11560 12154 11600 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11560 12072 11600 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11560 11990 11600 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11560 11908 11600 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11560 11826 11600 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11560 11744 11600 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11560 11662 11600 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11479 12482 11519 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11479 12400 11519 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11479 12318 11519 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11479 12236 11519 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11479 12154 11519 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11479 12072 11519 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11479 11990 11519 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11479 11908 11519 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11479 11826 11519 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11479 11744 11519 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11479 11662 11519 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11398 12482 11438 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11398 12400 11438 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11398 12318 11438 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11398 12236 11438 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11398 12154 11438 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11398 12072 11438 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11398 11990 11438 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11398 11908 11438 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11398 11826 11438 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11398 11744 11438 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11398 11662 11438 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11317 12482 11357 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11317 12400 11357 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11317 12318 11357 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11317 12236 11357 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11317 12154 11357 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11317 12072 11357 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11317 11990 11357 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11317 11908 11357 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11317 11826 11357 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11317 11744 11357 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11317 11662 11357 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11236 12482 11276 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11236 12400 11276 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11236 12318 11276 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11236 12236 11276 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11236 12154 11276 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11236 12072 11276 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11236 11990 11276 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11236 11908 11276 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11236 11826 11276 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11236 11744 11276 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11236 11662 11276 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11155 12482 11195 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11155 12400 11195 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11155 12318 11195 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11155 12236 11195 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11155 12154 11195 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11155 12072 11195 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11155 11990 11195 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11155 11908 11195 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11155 11826 11195 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11155 11744 11195 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11155 11662 11195 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11074 12482 11114 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11074 12400 11114 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11074 12318 11114 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11074 12236 11114 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11074 12154 11114 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11074 12072 11114 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11074 11990 11114 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11074 11908 11114 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11074 11826 11114 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11074 11744 11114 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 11074 11662 11114 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10993 12482 11033 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10993 12400 11033 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10993 12318 11033 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10993 12236 11033 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10993 12154 11033 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10993 12072 11033 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10993 11990 11033 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10993 11908 11033 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10993 11826 11033 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10993 11744 11033 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10993 11662 11033 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10912 12482 10952 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10912 12400 10952 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10912 12318 10952 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10912 12236 10952 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10912 12154 10952 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10912 12072 10952 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10912 11990 10952 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10912 11908 10952 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10912 11826 10952 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10912 11744 10952 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10912 11662 10952 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10831 12482 10871 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10831 12400 10871 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10831 12318 10871 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10831 12236 10871 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10831 12154 10871 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10831 12072 10871 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10831 11990 10871 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10831 11908 10871 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10831 11826 10871 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10831 11744 10871 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10831 11662 10871 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10750 12482 10790 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10750 12400 10790 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10750 12318 10790 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10750 12236 10790 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10750 12154 10790 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10750 12072 10790 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10750 11990 10790 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10750 11908 10790 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10750 11826 10790 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10750 11744 10790 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10750 11662 10790 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10669 12482 10709 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10669 12400 10709 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10669 12318 10709 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10669 12236 10709 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10669 12154 10709 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10669 12072 10709 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10669 11990 10709 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10669 11908 10709 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10669 11826 10709 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10669 11744 10709 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10669 11662 10709 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10588 12482 10628 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10588 12400 10628 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10588 12318 10628 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10588 12236 10628 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10588 12154 10628 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10588 12072 10628 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10588 11990 10628 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10588 11908 10628 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10588 11826 10628 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10588 11744 10628 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10588 11662 10628 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10506 12482 10546 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10506 12400 10546 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10506 12318 10546 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10506 12236 10546 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10506 12154 10546 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10506 12072 10546 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10506 11990 10546 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10506 11908 10546 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10506 11826 10546 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10506 11744 10546 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10506 11662 10546 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10424 12482 10464 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10424 12400 10464 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10424 12318 10464 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10424 12236 10464 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10424 12154 10464 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10424 12072 10464 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10424 11990 10464 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10424 11908 10464 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10424 11826 10464 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10424 11744 10464 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10424 11662 10464 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10342 12482 10382 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10342 12400 10382 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10342 12318 10382 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10342 12236 10382 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10342 12154 10382 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10342 12072 10382 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10342 11990 10382 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10342 11908 10382 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10342 11826 10382 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10342 11744 10382 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10342 11662 10382 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10260 12482 10300 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10260 12400 10300 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10260 12318 10300 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10260 12236 10300 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10260 12154 10300 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10260 12072 10300 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10260 11990 10300 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10260 11908 10300 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10260 11826 10300 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10260 11744 10300 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10260 11662 10300 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10178 12482 10218 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10178 12400 10218 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10178 12318 10218 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10178 12236 10218 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10178 12154 10218 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10178 12072 10218 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10178 11990 10218 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10178 11908 10218 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10178 11826 10218 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10178 11744 10218 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10178 11662 10218 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10096 12482 10136 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10096 12400 10136 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10096 12318 10136 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10096 12236 10136 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10096 12154 10136 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10096 12072 10136 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10096 11990 10136 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10096 11908 10136 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10096 11826 10136 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10096 11744 10136 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 10096 11662 10136 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4821 12482 4861 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4821 12400 4861 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4821 12318 4861 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4821 12236 4861 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4821 12154 4861 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4821 12072 4861 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4821 11990 4861 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4821 11908 4861 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4821 11826 4861 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4821 11744 4861 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4821 11662 4861 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4740 12482 4780 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4740 12400 4780 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4740 12318 4780 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4740 12236 4780 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4740 12154 4780 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4740 12072 4780 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4740 11990 4780 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4740 11908 4780 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4740 11826 4780 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4740 11744 4780 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4740 11662 4780 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4659 12482 4699 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4659 12400 4699 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4659 12318 4699 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4659 12236 4699 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4659 12154 4699 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4659 12072 4699 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4659 11990 4699 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4659 11908 4699 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4659 11826 4699 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4659 11744 4699 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4659 11662 4699 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4578 12482 4618 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4578 12400 4618 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4578 12318 4618 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4578 12236 4618 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4578 12154 4618 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4578 12072 4618 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4578 11990 4618 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4578 11908 4618 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4578 11826 4618 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4578 11744 4618 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4578 11662 4618 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4497 12482 4537 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4497 12400 4537 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4497 12318 4537 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4497 12236 4537 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4497 12154 4537 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4497 12072 4537 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4497 11990 4537 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4497 11908 4537 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4497 11826 4537 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4497 11744 4537 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4497 11662 4537 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4416 12482 4456 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4416 12400 4456 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4416 12318 4456 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4416 12236 4456 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4416 12154 4456 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4416 12072 4456 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4416 11990 4456 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4416 11908 4456 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4416 11826 4456 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4416 11744 4456 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4416 11662 4456 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4335 12482 4375 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4335 12400 4375 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4335 12318 4375 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4335 12236 4375 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4335 12154 4375 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4335 12072 4375 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4335 11990 4375 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4335 11908 4375 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4335 11826 4375 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4335 11744 4375 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4335 11662 4375 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4254 12482 4294 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4254 12400 4294 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4254 12318 4294 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4254 12236 4294 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4254 12154 4294 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4254 12072 4294 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4254 11990 4294 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4254 11908 4294 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4254 11826 4294 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4254 11744 4294 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4254 11662 4294 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4173 12482 4213 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4173 12400 4213 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4173 12318 4213 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4173 12236 4213 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4173 12154 4213 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4173 12072 4213 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4173 11990 4213 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4173 11908 4213 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4173 11826 4213 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4173 11744 4213 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4173 11662 4213 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4092 12482 4132 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4092 12400 4132 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4092 12318 4132 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4092 12236 4132 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4092 12154 4132 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4092 12072 4132 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4092 11990 4132 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4092 11908 4132 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4092 11826 4132 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4092 11744 4132 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4092 11662 4132 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4011 12482 4051 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4011 12400 4051 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4011 12318 4051 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4011 12236 4051 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4011 12154 4051 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4011 12072 4051 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4011 11990 4051 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4011 11908 4051 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4011 11826 4051 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4011 11744 4051 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 4011 11662 4051 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3930 12482 3970 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3930 12400 3970 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3930 12318 3970 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3930 12236 3970 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3930 12154 3970 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3930 12072 3970 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3930 11990 3970 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3930 11908 3970 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3930 11826 3970 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3930 11744 3970 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3930 11662 3970 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3849 12482 3889 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3849 12400 3889 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3849 12318 3889 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3849 12236 3889 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3849 12154 3889 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3849 12072 3889 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3849 11990 3889 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3849 11908 3889 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3849 11826 3889 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3849 11744 3889 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3849 11662 3889 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3768 12482 3808 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3768 12400 3808 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3768 12318 3808 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3768 12236 3808 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3768 12154 3808 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3768 12072 3808 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3768 11990 3808 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3768 11908 3808 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3768 11826 3808 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3768 11744 3808 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3768 11662 3808 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3687 12482 3727 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3687 12400 3727 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3687 12318 3727 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3687 12236 3727 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3687 12154 3727 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3687 12072 3727 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3687 11990 3727 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3687 11908 3727 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3687 11826 3727 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3687 11744 3727 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3687 11662 3727 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3606 12482 3646 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3606 12400 3646 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3606 12318 3646 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3606 12236 3646 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3606 12154 3646 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3606 12072 3646 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3606 11990 3646 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3606 11908 3646 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3606 11826 3646 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3606 11744 3646 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3606 11662 3646 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3525 12482 3565 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3525 12400 3565 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3525 12318 3565 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3525 12236 3565 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3525 12154 3565 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3525 12072 3565 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3525 11990 3565 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3525 11908 3565 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3525 11826 3565 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3525 11744 3565 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3525 11662 3565 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3444 12482 3484 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3444 12400 3484 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3444 12318 3484 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3444 12236 3484 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3444 12154 3484 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3444 12072 3484 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3444 11990 3484 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3444 11908 3484 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3444 11826 3484 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3444 11744 3484 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3444 11662 3484 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3363 12482 3403 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3363 12400 3403 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3363 12318 3403 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3363 12236 3403 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3363 12154 3403 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3363 12072 3403 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3363 11990 3403 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3363 11908 3403 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3363 11826 3403 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3363 11744 3403 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3363 11662 3403 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3282 12482 3322 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3282 12400 3322 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3282 12318 3322 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3282 12236 3322 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3282 12154 3322 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3282 12072 3322 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3282 11990 3322 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3282 11908 3322 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3282 11826 3322 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3282 11744 3322 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3282 11662 3322 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3201 12482 3241 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3201 12400 3241 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3201 12318 3241 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3201 12236 3241 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3201 12154 3241 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3201 12072 3241 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3201 11990 3241 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3201 11908 3241 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3201 11826 3241 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3201 11744 3241 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3201 11662 3241 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3120 12482 3160 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3120 12400 3160 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3120 12318 3160 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3120 12236 3160 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3120 12154 3160 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3120 12072 3160 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3120 11990 3160 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3120 11908 3160 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3120 11826 3160 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3120 11744 3160 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3120 11662 3160 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3039 12482 3079 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3039 12400 3079 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3039 12318 3079 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3039 12236 3079 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3039 12154 3079 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3039 12072 3079 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3039 11990 3079 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3039 11908 3079 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3039 11826 3079 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3039 11744 3079 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 3039 11662 3079 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2958 12482 2998 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2958 12400 2998 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2958 12318 2998 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2958 12236 2998 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2958 12154 2998 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2958 12072 2998 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2958 11990 2998 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2958 11908 2998 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2958 11826 2998 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2958 11744 2998 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2958 11662 2998 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2877 12482 2917 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2877 12400 2917 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2877 12318 2917 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2877 12236 2917 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2877 12154 2917 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2877 12072 2917 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2877 11990 2917 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2877 11908 2917 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2877 11826 2917 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2877 11744 2917 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2877 11662 2917 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2796 12482 2836 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2796 12400 2836 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2796 12318 2836 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2796 12236 2836 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2796 12154 2836 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2796 12072 2836 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2796 11990 2836 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2796 11908 2836 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2796 11826 2836 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2796 11744 2836 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2796 11662 2836 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2715 12482 2755 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2715 12400 2755 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2715 12318 2755 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2715 12236 2755 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2715 12154 2755 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2715 12072 2755 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2715 11990 2755 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2715 11908 2755 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2715 11826 2755 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2715 11744 2755 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2715 11662 2755 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2634 12482 2674 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2634 12400 2674 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2634 12318 2674 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2634 12236 2674 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2634 12154 2674 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2634 12072 2674 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2634 11990 2674 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2634 11908 2674 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2634 11826 2674 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2634 11744 2674 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2634 11662 2674 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2553 12482 2593 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2553 12400 2593 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2553 12318 2593 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2553 12236 2593 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2553 12154 2593 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2553 12072 2593 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2553 11990 2593 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2553 11908 2593 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2553 11826 2593 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2553 11744 2593 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2553 11662 2593 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2472 12482 2512 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2472 12400 2512 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2472 12318 2512 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2472 12236 2512 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2472 12154 2512 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2472 12072 2512 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2472 11990 2512 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2472 11908 2512 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2472 11826 2512 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2472 11744 2512 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2472 11662 2512 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2391 12482 2431 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2391 12400 2431 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2391 12318 2431 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2391 12236 2431 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2391 12154 2431 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2391 12072 2431 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2391 11990 2431 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2391 11908 2431 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2391 11826 2431 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2391 11744 2431 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2391 11662 2431 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2310 12482 2350 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2310 12400 2350 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2310 12318 2350 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2310 12236 2350 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2310 12154 2350 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2310 12072 2350 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2310 11990 2350 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2310 11908 2350 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2310 11826 2350 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2310 11744 2350 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2310 11662 2350 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2229 12482 2269 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2229 12400 2269 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2229 12318 2269 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2229 12236 2269 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2229 12154 2269 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2229 12072 2269 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2229 11990 2269 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2229 11908 2269 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2229 11826 2269 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2229 11744 2269 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2229 11662 2269 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2148 12482 2188 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2148 12400 2188 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2148 12318 2188 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2148 12236 2188 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2148 12154 2188 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2148 12072 2188 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2148 11990 2188 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2148 11908 2188 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2148 11826 2188 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2148 11744 2188 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2148 11662 2188 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2067 12482 2107 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2067 12400 2107 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2067 12318 2107 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2067 12236 2107 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2067 12154 2107 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2067 12072 2107 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2067 11990 2107 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2067 11908 2107 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2067 11826 2107 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2067 11744 2107 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 2067 11662 2107 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1986 12482 2026 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1986 12400 2026 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1986 12318 2026 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1986 12236 2026 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1986 12154 2026 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1986 12072 2026 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1986 11990 2026 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1986 11908 2026 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1986 11826 2026 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1986 11744 2026 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1986 11662 2026 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1905 12482 1945 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1905 12400 1945 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1905 12318 1945 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1905 12236 1945 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1905 12154 1945 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1905 12072 1945 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1905 11990 1945 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1905 11908 1945 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1905 11826 1945 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1905 11744 1945 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1905 11662 1945 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1824 12482 1864 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1824 12400 1864 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1824 12318 1864 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1824 12236 1864 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1824 12154 1864 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1824 12072 1864 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1824 11990 1864 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1824 11908 1864 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1824 11826 1864 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1824 11744 1864 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1824 11662 1864 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1743 12482 1783 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1743 12400 1783 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1743 12318 1783 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1743 12236 1783 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1743 12154 1783 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1743 12072 1783 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1743 11990 1783 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1743 11908 1783 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1743 11826 1783 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1743 11744 1783 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1743 11662 1783 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1662 12482 1702 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1662 12400 1702 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1662 12318 1702 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1662 12236 1702 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1662 12154 1702 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1662 12072 1702 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1662 11990 1702 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1662 11908 1702 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1662 11826 1702 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1662 11744 1702 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1662 11662 1702 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1581 12482 1621 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1581 12400 1621 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1581 12318 1621 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1581 12236 1621 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1581 12154 1621 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1581 12072 1621 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1581 11990 1621 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1581 11908 1621 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1581 11826 1621 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1581 11744 1621 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1581 11662 1621 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1500 12482 1540 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1500 12400 1540 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1500 12318 1540 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1500 12236 1540 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1500 12154 1540 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1500 12072 1540 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1500 11990 1540 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1500 11908 1540 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1500 11826 1540 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1500 11744 1540 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1500 11662 1540 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1419 12482 1459 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1419 12400 1459 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1419 12318 1459 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1419 12236 1459 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1419 12154 1459 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1419 12072 1459 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1419 11990 1459 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1419 11908 1459 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1419 11826 1459 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1419 11744 1459 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1419 11662 1459 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1338 12482 1378 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1338 12400 1378 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1338 12318 1378 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1338 12236 1378 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1338 12154 1378 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1338 12072 1378 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1338 11990 1378 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1338 11908 1378 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1338 11826 1378 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1338 11744 1378 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1338 11662 1378 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1257 12482 1297 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1257 12400 1297 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1257 12318 1297 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1257 12236 1297 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1257 12154 1297 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1257 12072 1297 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1257 11990 1297 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1257 11908 1297 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1257 11826 1297 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1257 11744 1297 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1257 11662 1297 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1176 12482 1216 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1176 12400 1216 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1176 12318 1216 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1176 12236 1216 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1176 12154 1216 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1176 12072 1216 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1176 11990 1216 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1176 11908 1216 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1176 11826 1216 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1176 11744 1216 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1176 11662 1216 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1095 12482 1135 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1095 12400 1135 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1095 12318 1135 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1095 12236 1135 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1095 12154 1135 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1095 12072 1135 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1095 11990 1135 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1095 11908 1135 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1095 11826 1135 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1095 11744 1135 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1095 11662 1135 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1014 12482 1054 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1014 12400 1054 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1014 12318 1054 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1014 12236 1054 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1014 12154 1054 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1014 12072 1054 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1014 11990 1054 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1014 11908 1054 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1014 11826 1054 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1014 11744 1054 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 1014 11662 1054 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 933 12482 973 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 933 12400 973 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 933 12318 973 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 933 12236 973 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 933 12154 973 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 933 12072 973 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 933 11990 973 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 933 11908 973 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 933 11826 973 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 933 11744 973 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 933 11662 973 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 852 12482 892 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 852 12400 892 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 852 12318 892 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 852 12236 892 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 852 12154 892 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 852 12072 892 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 852 11990 892 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 852 11908 892 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 852 11826 892 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 852 11744 892 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 852 11662 892 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 771 12482 811 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 771 12400 811 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 771 12318 811 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 771 12236 811 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 771 12154 811 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 771 12072 811 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 771 11990 811 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 771 11908 811 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 771 11826 811 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 771 11744 811 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 771 11662 811 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 690 12482 730 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 690 12400 730 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 690 12318 730 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 690 12236 730 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 690 12154 730 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 690 12072 730 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 690 11990 730 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 690 11908 730 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 690 11826 730 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 690 11744 730 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 690 11662 730 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 609 12482 649 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 609 12400 649 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 609 12318 649 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 609 12236 649 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 609 12154 649 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 609 12072 649 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 609 11990 649 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 609 11908 649 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 609 11826 649 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 609 11744 649 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 609 11662 649 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 527 12482 567 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 527 12400 567 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 527 12318 567 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 527 12236 567 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 527 12154 567 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 527 12072 567 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 527 11990 567 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 527 11908 567 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 527 11826 567 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 527 11744 567 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 527 11662 567 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 445 12482 485 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 445 12400 485 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 445 12318 485 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 445 12236 485 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 445 12154 485 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 445 12072 485 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 445 11990 485 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 445 11908 485 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 445 11826 485 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 445 11744 485 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 445 11662 485 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 363 12482 403 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 363 12400 403 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 363 12318 403 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 363 12236 403 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 363 12154 403 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 363 12072 403 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 363 11990 403 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 363 11908 403 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 363 11826 403 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 363 11744 403 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 363 11662 403 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 281 12482 321 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 281 12400 321 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 281 12318 321 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 281 12236 321 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 281 12154 321 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 281 12072 321 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 281 11990 321 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 281 11908 321 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 281 11826 321 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 281 11744 321 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 281 11662 321 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 199 12482 239 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 199 12400 239 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 199 12318 239 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 199 12236 239 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 199 12154 239 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 199 12072 239 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 199 11990 239 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 199 11908 239 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 199 11826 239 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 199 11744 239 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 199 11662 239 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 117 12482 157 12522 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 117 12400 157 12440 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 117 12318 157 12358 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 117 12236 157 12276 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 117 12154 157 12194 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 117 12072 157 12112 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 117 11990 157 12030 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 117 11908 157 11948 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 117 11826 157 11866 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 117 11744 157 11784 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal3 s 117 11662 157 11702 6 VSSIO_Q
port 7 nsew ground bidirectional
rlabel metal5 s 0 3007 193 3657 6 VDDA
port 8 nsew power bidirectional
rlabel metal5 s 14807 3007 15000 3657 6 VDDA
port 8 nsew power bidirectional
rlabel metal4 s 0 2987 193 3677 6 VDDA
port 8 nsew power bidirectional
rlabel metal4 s 14807 2987 15000 3677 6 VDDA
port 8 nsew power bidirectional
rlabel metal4 s 14807 2987 15000 3677 6 VDDA
port 8 nsew power bidirectional
rlabel metal5 s 0 3007 193 3657 6 VDDA
port 8 nsew power bidirectional
rlabel metal5 s 14807 3007 15000 3657 6 VDDA
port 8 nsew power bidirectional
rlabel metal4 s 14807 2987 15000 3677 6 VDDA
port 8 nsew power bidirectional
rlabel metal5 s 0 3007 193 3657 6 VDDA
port 8 nsew power bidirectional
rlabel metal5 s 14807 3007 15000 3657 6 VDDA
port 8 nsew power bidirectional
rlabel metal5 s 0 1797 254 2687 6 VCCD
port 9 nsew power bidirectional
rlabel metal5 s 14746 1797 15000 2687 6 VCCD
port 9 nsew power bidirectional
rlabel metal4 s 0 1777 254 2707 6 VCCD
port 9 nsew power bidirectional
rlabel metal4 s 14746 1777 15000 2707 6 VCCD
port 9 nsew power bidirectional
rlabel metal4 s 14746 1777 15000 2707 6 VCCD
port 9 nsew power bidirectional
rlabel metal5 s 0 1797 254 2687 6 VCCD
port 9 nsew power bidirectional
rlabel metal5 s 14746 1797 15000 2687 6 VCCD
port 9 nsew power bidirectional
rlabel metal4 s 14746 1777 15000 2707 6 VCCD
port 9 nsew power bidirectional
rlabel metal5 s 0 1797 254 2687 6 VCCD
port 9 nsew power bidirectional
rlabel metal5 s 14746 1797 15000 2687 6 VCCD
port 9 nsew power bidirectional
rlabel metal5 s 0 427 254 1477 6 VCCHIB
port 10 nsew power bidirectional
rlabel metal5 s 14746 427 15000 1477 6 VCCHIB
port 10 nsew power bidirectional
rlabel metal4 s 0 407 254 1497 6 VCCHIB
port 10 nsew power bidirectional
rlabel metal4 s 14746 407 15000 1497 6 VCCHIB
port 10 nsew power bidirectional
rlabel metal4 s 14746 407 15000 1497 6 VCCHIB
port 10 nsew power bidirectional
rlabel metal5 s 0 427 254 1477 6 VCCHIB
port 10 nsew power bidirectional
rlabel metal5 s 14746 427 15000 1477 6 VCCHIB
port 10 nsew power bidirectional
rlabel metal4 s 14746 407 15000 1497 6 VCCHIB
port 10 nsew power bidirectional
rlabel metal5 s 0 427 254 1477 6 VCCHIB
port 10 nsew power bidirectional
rlabel metal5 s 14746 427 15000 1477 6 VCCHIB
port 10 nsew power bidirectional
rlabel metal4 s 0 9673 15000 10269 6 AMUXBUS_B
port 11 nsew signal bidirectional
rlabel metal4 s 14746 9673 15000 10269 6 AMUXBUS_B
port 11 nsew signal bidirectional
rlabel metal4 s 14746 9673 15000 10269 6 AMUXBUS_B
port 11 nsew signal bidirectional
rlabel metal4 s 14746 9673 15000 10269 6 AMUXBUS_B
port 11 nsew signal bidirectional
rlabel metal4 s 0 10625 15000 11221 6 AMUXBUS_A
port 12 nsew signal bidirectional
rlabel metal4 s 14746 10625 15000 11221 6 AMUXBUS_A
port 12 nsew signal bidirectional
rlabel metal4 s 14746 10625 15000 11221 6 AMUXBUS_A
port 12 nsew signal bidirectional
rlabel metal4 s 14746 10625 15000 11221 6 AMUXBUS_A
port 12 nsew signal bidirectional
<< properties >>
string LEFclass PAD
string FIXED_BBOX 0 0 15000 40000
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 22420376
string GDS_START 21945206
<< end >>
