magic
tech sky130A
magscale 1 2
timestamp 1624883981
<< checkpaint >>
rect -1260 -1349 1904 1563
<< nwell >>
rect 0 0 644 240
<< pmos >>
rect 95 36 125 204
rect 181 36 211 204
rect 267 36 297 204
rect 353 36 383 204
rect 439 36 469 204
rect 525 36 555 204
<< pdiff >>
rect 42 173 95 204
rect 42 139 50 173
rect 84 139 95 173
rect 42 101 95 139
rect 42 67 50 101
rect 84 67 95 101
rect 42 36 95 67
rect 125 173 181 204
rect 125 139 136 173
rect 170 139 181 173
rect 125 101 181 139
rect 125 67 136 101
rect 170 67 181 101
rect 125 36 181 67
rect 211 173 267 204
rect 211 139 222 173
rect 256 139 267 173
rect 211 101 267 139
rect 211 67 222 101
rect 256 67 267 101
rect 211 36 267 67
rect 297 173 353 204
rect 297 139 308 173
rect 342 139 353 173
rect 297 101 353 139
rect 297 67 308 101
rect 342 67 353 101
rect 297 36 353 67
rect 383 173 439 204
rect 383 139 394 173
rect 428 139 439 173
rect 383 101 439 139
rect 383 67 394 101
rect 428 67 439 101
rect 383 36 439 67
rect 469 173 525 204
rect 469 139 480 173
rect 514 139 525 173
rect 469 101 525 139
rect 469 67 480 101
rect 514 67 525 101
rect 469 36 525 67
rect 555 173 608 204
rect 555 139 566 173
rect 600 139 608 173
rect 555 101 608 139
rect 555 67 566 101
rect 600 67 608 101
rect 555 36 608 67
<< pdiffc >>
rect 50 139 84 173
rect 50 67 84 101
rect 136 139 170 173
rect 136 67 170 101
rect 222 139 256 173
rect 222 67 256 101
rect 308 139 342 173
rect 308 67 342 101
rect 394 139 428 173
rect 394 67 428 101
rect 480 139 514 173
rect 480 67 514 101
rect 566 139 600 173
rect 566 67 600 101
<< poly >>
rect 95 287 555 303
rect 95 253 138 287
rect 172 253 206 287
rect 240 253 274 287
rect 308 253 342 287
rect 376 253 410 287
rect 444 253 478 287
rect 512 253 555 287
rect 95 230 555 253
rect 95 204 125 230
rect 181 204 211 230
rect 267 204 297 230
rect 353 204 383 230
rect 439 204 469 230
rect 525 204 555 230
rect 95 10 125 36
rect 181 10 211 36
rect 267 10 297 36
rect 353 10 383 36
rect 439 10 469 36
rect 525 10 555 36
<< polycont >>
rect 138 253 172 287
rect 206 253 240 287
rect 274 253 308 287
rect 342 253 376 287
rect 410 253 444 287
rect 478 253 512 287
<< locali >>
rect 122 287 528 303
rect 122 253 128 287
rect 172 253 200 287
rect 240 253 272 287
rect 308 253 342 287
rect 378 253 410 287
rect 450 253 478 287
rect 522 253 528 287
rect 122 235 528 253
rect 50 173 84 189
rect 50 101 84 139
rect 50 51 84 67
rect 136 173 170 189
rect 136 101 170 139
rect 136 51 170 67
rect 222 173 256 189
rect 222 101 256 139
rect 222 51 256 67
rect 308 173 342 189
rect 308 101 342 139
rect 308 51 342 67
rect 394 173 428 189
rect 394 101 428 139
rect 394 51 428 67
rect 480 173 514 189
rect 480 101 514 139
rect 480 51 514 67
rect 566 173 600 189
rect 566 101 600 139
rect 566 51 600 67
<< viali >>
rect 128 253 138 287
rect 138 253 162 287
rect 200 253 206 287
rect 206 253 234 287
rect 272 253 274 287
rect 274 253 306 287
rect 344 253 376 287
rect 376 253 378 287
rect 416 253 444 287
rect 444 253 450 287
rect 488 253 512 287
rect 512 253 522 287
rect 50 139 84 173
rect 50 67 84 101
rect 136 139 170 173
rect 136 67 170 101
rect 222 139 256 173
rect 222 67 256 101
rect 308 139 342 173
rect 308 67 342 101
rect 394 139 428 173
rect 394 67 428 101
rect 480 139 514 173
rect 480 67 514 101
rect 566 139 600 173
rect 566 67 600 101
<< metal1 >>
rect 116 287 534 299
rect 116 253 128 287
rect 162 253 200 287
rect 234 253 272 287
rect 306 253 344 287
rect 378 253 416 287
rect 450 253 488 287
rect 522 253 534 287
rect 116 241 534 253
rect 44 173 90 189
rect 44 139 50 173
rect 84 139 90 173
rect 44 101 90 139
rect 44 67 50 101
rect 84 67 90 101
rect 44 -29 90 67
rect 127 178 179 189
rect 127 114 179 126
rect 127 51 179 62
rect 216 173 262 189
rect 216 139 222 173
rect 256 139 262 173
rect 216 101 262 139
rect 216 67 222 101
rect 256 67 262 101
rect 216 -29 262 67
rect 299 178 351 189
rect 299 114 351 126
rect 299 51 351 62
rect 388 173 434 189
rect 388 139 394 173
rect 428 139 434 173
rect 388 101 434 139
rect 388 67 394 101
rect 428 67 434 101
rect 388 -29 434 67
rect 471 178 523 189
rect 471 114 523 126
rect 471 51 523 62
rect 560 173 606 189
rect 560 139 566 173
rect 600 139 606 173
rect 560 101 606 139
rect 560 67 566 101
rect 600 67 606 101
rect 560 -29 606 67
rect 44 -89 606 -29
<< via1 >>
rect 127 173 179 178
rect 127 139 136 173
rect 136 139 170 173
rect 170 139 179 173
rect 127 126 179 139
rect 127 101 179 114
rect 127 67 136 101
rect 136 67 170 101
rect 170 67 179 101
rect 127 62 179 67
rect 299 173 351 178
rect 299 139 308 173
rect 308 139 342 173
rect 342 139 351 173
rect 299 126 351 139
rect 299 101 351 114
rect 299 67 308 101
rect 308 67 342 101
rect 342 67 351 101
rect 299 62 351 67
rect 471 173 523 178
rect 471 139 480 173
rect 480 139 514 173
rect 514 139 523 173
rect 471 126 523 139
rect 471 101 523 114
rect 471 67 480 101
rect 480 67 514 101
rect 514 67 523 101
rect 471 62 523 67
<< metal2 >>
rect 120 188 186 197
rect 120 132 125 188
rect 181 132 186 188
rect 120 126 127 132
rect 179 126 186 132
rect 120 114 186 126
rect 120 108 127 114
rect 179 108 186 114
rect 120 52 125 108
rect 181 52 186 108
rect 120 43 186 52
rect 292 188 358 197
rect 292 132 297 188
rect 353 132 358 188
rect 292 126 299 132
rect 351 126 358 132
rect 292 114 358 126
rect 292 108 299 114
rect 351 108 358 114
rect 292 52 297 108
rect 353 52 358 108
rect 292 43 358 52
rect 464 188 530 197
rect 464 132 469 188
rect 525 132 530 188
rect 464 126 471 132
rect 523 126 530 132
rect 464 114 530 126
rect 464 108 471 114
rect 523 108 530 114
rect 464 52 469 108
rect 525 52 530 108
rect 464 43 530 52
<< via2 >>
rect 125 178 181 188
rect 125 132 127 178
rect 127 132 179 178
rect 179 132 181 178
rect 125 62 127 108
rect 127 62 179 108
rect 179 62 181 108
rect 125 52 181 62
rect 297 178 353 188
rect 297 132 299 178
rect 299 132 351 178
rect 351 132 353 178
rect 297 62 299 108
rect 299 62 351 108
rect 351 62 353 108
rect 297 52 353 62
rect 469 178 525 188
rect 469 132 471 178
rect 471 132 523 178
rect 523 132 525 178
rect 469 62 471 108
rect 471 62 523 108
rect 523 62 525 108
rect 469 52 525 62
<< metal3 >>
rect 120 188 530 197
rect 120 132 125 188
rect 181 132 297 188
rect 353 132 469 188
rect 525 132 530 188
rect 120 131 530 132
rect 120 108 186 131
rect 120 52 125 108
rect 181 52 186 108
rect 120 43 186 52
rect 292 108 358 131
rect 292 52 297 108
rect 353 52 358 108
rect 292 43 358 52
rect 464 108 530 131
rect 464 52 469 108
rect 525 52 530 108
rect 464 43 530 52
<< labels >>
flabel metal3 s 120 131 530 197 0 FreeSans 400 0 0 0 DRAIN
port 1 nsew
flabel metal1 s 44 -89 606 -29 0 FreeSans 400 0 0 0 SOURCE
port 2 nsew
flabel metal1 s 116 241 534 299 0 FreeSans 400 0 0 0 GATE
port 3 nsew
flabel nwell s 84 232 91 238 0 FreeSans 400 0 0 0 BULK
port 4 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 9196312
string GDS_START 9186848
string path 1.675 4.725 1.675 -2.225 
<< end >>
