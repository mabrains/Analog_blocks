magic
tech sky130A
magscale 1 2
timestamp 1624883981
<< checkpaint >>
rect -1260 -1260 2136 2178
<< pwell >>
rect 467 350 491 401
<< poly >>
rect 0 902 876 918
rect 0 868 80 902
rect 114 868 148 902
rect 182 868 216 902
rect 250 868 284 902
rect 318 868 352 902
rect 386 868 420 902
rect 454 868 488 902
rect 522 868 556 902
rect 590 868 624 902
rect 658 868 692 902
rect 726 868 760 902
rect 794 868 876 902
rect 0 816 876 868
rect 0 782 16 816
rect 50 782 826 816
rect 860 782 876 816
rect 0 748 876 782
rect 0 714 16 748
rect 50 714 826 748
rect 860 714 876 748
rect 0 680 876 714
rect 0 646 16 680
rect 50 646 826 680
rect 860 646 876 680
rect 0 612 876 646
rect 0 578 16 612
rect 50 578 826 612
rect 860 578 876 612
rect 0 544 876 578
rect 0 510 16 544
rect 50 510 826 544
rect 860 510 876 544
rect 0 476 876 510
rect 0 442 16 476
rect 50 442 826 476
rect 860 442 876 476
rect 0 408 876 442
rect 0 374 16 408
rect 50 374 826 408
rect 860 374 876 408
rect 0 340 876 374
rect 0 306 16 340
rect 50 306 826 340
rect 860 306 876 340
rect 0 272 876 306
rect 0 238 16 272
rect 50 238 826 272
rect 860 238 876 272
rect 0 204 876 238
rect 0 170 16 204
rect 50 170 826 204
rect 860 170 876 204
rect 0 136 876 170
rect 0 102 16 136
rect 50 102 826 136
rect 860 102 876 136
rect 0 50 876 102
rect 0 16 80 50
rect 114 16 148 50
rect 182 16 216 50
rect 250 16 284 50
rect 318 16 352 50
rect 386 16 420 50
rect 454 16 488 50
rect 522 16 556 50
rect 590 16 624 50
rect 658 16 692 50
rect 726 16 760 50
rect 794 16 876 50
rect 0 0 876 16
<< polycont >>
rect 80 868 114 902
rect 148 868 182 902
rect 216 868 250 902
rect 284 868 318 902
rect 352 868 386 902
rect 420 868 454 902
rect 488 868 522 902
rect 556 868 590 902
rect 624 868 658 902
rect 692 868 726 902
rect 760 868 794 902
rect 16 782 50 816
rect 826 782 860 816
rect 16 714 50 748
rect 826 714 860 748
rect 16 646 50 680
rect 826 646 860 680
rect 16 578 50 612
rect 826 578 860 612
rect 16 510 50 544
rect 826 510 860 544
rect 16 442 50 476
rect 826 442 860 476
rect 16 374 50 408
rect 826 374 860 408
rect 16 306 50 340
rect 826 306 860 340
rect 16 238 50 272
rect 826 238 860 272
rect 16 170 50 204
rect 826 170 860 204
rect 16 102 50 136
rect 826 102 860 136
rect 80 16 114 50
rect 148 16 182 50
rect 216 16 250 50
rect 284 16 318 50
rect 352 16 386 50
rect 420 16 454 50
rect 488 16 522 50
rect 556 16 590 50
rect 624 16 658 50
rect 692 16 726 50
rect 760 16 794 50
<< locali >>
rect 0 902 876 918
rect 0 868 80 902
rect 131 868 148 902
rect 203 868 216 902
rect 275 868 284 902
rect 347 868 352 902
rect 419 868 420 902
rect 454 868 457 902
rect 522 868 529 902
rect 590 868 601 902
rect 658 868 673 902
rect 726 868 745 902
rect 794 868 876 902
rect 0 852 876 868
rect 0 836 66 852
rect 0 782 16 836
rect 50 782 66 836
rect 810 836 876 852
rect 100 784 776 816
rect 100 782 421 784
rect 0 764 66 782
rect 0 714 16 764
rect 50 746 66 764
rect 411 750 421 782
rect 455 782 776 784
rect 810 782 826 836
rect 860 782 876 836
rect 455 750 465 782
rect 50 714 377 746
rect 0 712 377 714
rect 411 712 465 750
rect 810 764 876 782
rect 810 746 826 764
rect 499 714 826 746
rect 860 714 876 764
rect 499 712 876 714
rect 0 692 66 712
rect 0 646 16 692
rect 50 646 66 692
rect 411 678 421 712
rect 455 678 465 712
rect 411 676 465 678
rect 810 692 876 712
rect 0 620 66 646
rect 100 642 776 676
rect 810 646 826 692
rect 860 646 876 692
rect 0 578 16 620
rect 50 606 66 620
rect 411 640 465 642
rect 411 606 421 640
rect 455 606 465 640
rect 810 620 876 646
rect 810 606 826 620
rect 50 578 377 606
rect 0 572 377 578
rect 0 548 66 572
rect 0 510 16 548
rect 50 510 66 548
rect 411 568 465 606
rect 499 578 826 606
rect 860 578 876 620
rect 499 572 876 578
rect 411 536 421 568
rect 0 476 66 510
rect 100 534 421 536
rect 455 536 465 568
rect 810 548 876 572
rect 455 534 776 536
rect 100 502 776 534
rect 810 510 826 548
rect 860 510 876 548
rect 0 442 16 476
rect 50 442 66 476
rect 0 408 66 442
rect 411 416 465 502
rect 810 476 876 510
rect 810 442 826 476
rect 860 442 876 476
rect 0 370 16 408
rect 50 370 66 408
rect 100 384 776 416
rect 100 382 421 384
rect 0 346 66 370
rect 411 350 421 382
rect 455 382 776 384
rect 810 408 876 442
rect 455 350 465 382
rect 0 340 377 346
rect 0 298 16 340
rect 50 312 377 340
rect 411 312 465 350
rect 810 370 826 408
rect 860 370 876 408
rect 810 346 876 370
rect 499 340 876 346
rect 499 312 826 340
rect 50 298 66 312
rect 0 272 66 298
rect 411 278 421 312
rect 455 278 465 312
rect 411 276 465 278
rect 810 298 826 312
rect 860 298 876 340
rect 0 226 16 272
rect 50 226 66 272
rect 100 242 776 276
rect 810 272 876 298
rect 0 206 66 226
rect 411 240 465 242
rect 411 206 421 240
rect 455 206 465 240
rect 810 226 826 272
rect 860 226 876 272
rect 810 206 876 226
rect 0 204 377 206
rect 0 154 16 204
rect 50 172 377 204
rect 50 154 66 172
rect 0 136 66 154
rect 411 168 465 206
rect 499 204 876 206
rect 499 172 826 204
rect 411 136 421 168
rect 0 82 16 136
rect 50 82 66 136
rect 100 134 421 136
rect 455 136 465 168
rect 810 154 826 172
rect 860 154 876 204
rect 810 136 876 154
rect 455 134 776 136
rect 100 102 776 134
rect 0 66 66 82
rect 810 82 826 136
rect 860 82 876 136
rect 810 66 876 82
rect 0 50 876 66
rect 0 16 80 50
rect 131 16 148 50
rect 203 16 216 50
rect 275 16 284 50
rect 347 16 352 50
rect 419 16 420 50
rect 454 16 457 50
rect 522 16 529 50
rect 590 16 601 50
rect 658 16 673 50
rect 726 16 745 50
rect 794 16 876 50
rect 0 0 876 16
<< viali >>
rect 97 868 114 902
rect 114 868 131 902
rect 169 868 182 902
rect 182 868 203 902
rect 241 868 250 902
rect 250 868 275 902
rect 313 868 318 902
rect 318 868 347 902
rect 385 868 386 902
rect 386 868 419 902
rect 457 868 488 902
rect 488 868 491 902
rect 529 868 556 902
rect 556 868 563 902
rect 601 868 624 902
rect 624 868 635 902
rect 673 868 692 902
rect 692 868 707 902
rect 745 868 760 902
rect 760 868 779 902
rect 16 816 50 836
rect 16 802 50 816
rect 16 748 50 764
rect 16 730 50 748
rect 421 750 455 784
rect 826 816 860 836
rect 826 802 860 816
rect 826 748 860 764
rect 826 730 860 748
rect 16 680 50 692
rect 16 658 50 680
rect 421 678 455 712
rect 826 680 860 692
rect 826 658 860 680
rect 16 612 50 620
rect 16 586 50 612
rect 421 606 455 640
rect 826 612 860 620
rect 16 544 50 548
rect 16 514 50 544
rect 826 586 860 612
rect 421 534 455 568
rect 826 544 860 548
rect 826 514 860 544
rect 16 442 50 476
rect 826 442 860 476
rect 16 374 50 404
rect 16 370 50 374
rect 421 350 455 384
rect 16 306 50 332
rect 826 374 860 404
rect 826 370 860 374
rect 16 298 50 306
rect 421 278 455 312
rect 826 306 860 332
rect 826 298 860 306
rect 16 238 50 260
rect 16 226 50 238
rect 421 206 455 240
rect 826 238 860 260
rect 826 226 860 238
rect 16 170 50 188
rect 16 154 50 170
rect 16 102 50 116
rect 16 82 50 102
rect 421 134 455 168
rect 826 170 860 188
rect 826 154 860 170
rect 826 102 860 116
rect 826 82 860 102
rect 97 16 114 50
rect 114 16 131 50
rect 169 16 182 50
rect 182 16 203 50
rect 241 16 250 50
rect 250 16 275 50
rect 313 16 318 50
rect 318 16 347 50
rect 385 16 386 50
rect 386 16 419 50
rect 457 16 488 50
rect 488 16 491 50
rect 529 16 556 50
rect 556 16 563 50
rect 601 16 624 50
rect 624 16 635 50
rect 673 16 692 50
rect 692 16 707 50
rect 745 16 760 50
rect 760 16 779 50
<< metal1 >>
rect 0 911 876 918
rect 0 859 52 911
rect 104 902 116 911
rect 168 902 180 911
rect 232 902 244 911
rect 168 868 169 902
rect 232 868 241 902
rect 104 859 116 868
rect 168 859 180 868
rect 232 859 244 868
rect 296 859 308 911
rect 360 902 516 911
rect 360 868 385 902
rect 419 868 457 902
rect 491 868 516 902
rect 360 859 516 868
rect 568 859 580 911
rect 632 902 644 911
rect 696 902 708 911
rect 760 902 772 911
rect 635 868 644 902
rect 707 868 708 902
rect 632 859 644 868
rect 696 859 708 868
rect 760 859 772 868
rect 824 859 876 911
rect 0 852 876 859
rect 0 842 66 852
rect 0 790 7 842
rect 59 790 66 842
rect 0 778 66 790
rect 0 726 7 778
rect 59 726 66 778
rect 0 714 66 726
rect 0 662 7 714
rect 59 662 66 714
rect 0 658 16 662
rect 50 658 66 662
rect 0 650 66 658
rect 0 598 7 650
rect 59 598 66 650
rect 0 586 16 598
rect 50 586 66 598
rect 0 534 7 586
rect 59 534 66 586
rect 0 514 16 534
rect 50 514 66 534
rect 0 476 66 514
rect 0 442 16 476
rect 50 442 66 476
rect 0 404 66 442
rect 0 384 16 404
rect 50 384 66 404
rect 0 332 7 384
rect 59 332 66 384
rect 0 320 16 332
rect 50 320 66 332
rect 0 268 7 320
rect 59 268 66 320
rect 0 260 66 268
rect 0 256 16 260
rect 50 256 66 260
rect 0 204 7 256
rect 59 204 66 256
rect 0 192 66 204
rect 0 140 7 192
rect 59 140 66 192
rect 0 128 66 140
rect 0 76 7 128
rect 59 76 66 128
rect 113 491 141 824
rect 169 519 197 852
rect 225 491 253 824
rect 281 519 309 852
rect 337 491 365 824
rect 411 818 465 824
rect 411 766 412 818
rect 464 766 465 818
rect 411 754 421 766
rect 455 754 465 766
rect 411 702 412 754
rect 464 702 465 754
rect 411 690 421 702
rect 455 690 465 702
rect 411 638 412 690
rect 464 638 465 690
rect 411 626 421 638
rect 455 626 465 638
rect 411 574 412 626
rect 464 574 465 626
rect 411 568 465 574
rect 411 562 421 568
rect 455 562 465 568
rect 411 510 412 562
rect 464 510 465 562
rect 411 491 465 510
rect 511 491 539 824
rect 567 519 595 852
rect 623 491 651 824
rect 679 519 707 852
rect 810 842 876 852
rect 735 491 763 824
rect 113 485 763 491
rect 113 433 119 485
rect 171 433 183 485
rect 235 433 247 485
rect 299 433 311 485
rect 363 433 513 485
rect 565 433 577 485
rect 629 433 641 485
rect 693 433 705 485
rect 757 433 763 485
rect 113 427 763 433
rect 113 94 141 427
rect 0 66 66 76
rect 169 66 197 399
rect 225 94 253 427
rect 281 66 309 399
rect 337 94 365 427
rect 411 408 465 427
rect 411 356 412 408
rect 464 356 465 408
rect 411 350 421 356
rect 455 350 465 356
rect 411 344 465 350
rect 411 292 412 344
rect 464 292 465 344
rect 411 280 421 292
rect 455 280 465 292
rect 411 228 412 280
rect 464 228 465 280
rect 411 216 421 228
rect 455 216 465 228
rect 411 164 412 216
rect 464 164 465 216
rect 411 152 421 164
rect 455 152 465 164
rect 411 100 412 152
rect 464 100 465 152
rect 411 94 465 100
rect 511 94 539 427
rect 567 66 595 399
rect 623 94 651 427
rect 679 66 707 399
rect 735 94 763 427
rect 810 790 817 842
rect 869 790 876 842
rect 810 778 876 790
rect 810 726 817 778
rect 869 726 876 778
rect 810 714 876 726
rect 810 662 817 714
rect 869 662 876 714
rect 810 658 826 662
rect 860 658 876 662
rect 810 650 876 658
rect 810 598 817 650
rect 869 598 876 650
rect 810 586 826 598
rect 860 586 876 598
rect 810 534 817 586
rect 869 534 876 586
rect 810 514 826 534
rect 860 514 876 534
rect 810 476 876 514
rect 810 442 826 476
rect 860 442 876 476
rect 810 404 876 442
rect 810 384 826 404
rect 860 384 876 404
rect 810 332 817 384
rect 869 332 876 384
rect 810 320 826 332
rect 860 320 876 332
rect 810 268 817 320
rect 869 268 876 320
rect 810 260 876 268
rect 810 256 826 260
rect 860 256 876 260
rect 810 204 817 256
rect 869 204 876 256
rect 810 192 876 204
rect 810 140 817 192
rect 869 140 876 192
rect 810 128 876 140
rect 810 76 817 128
rect 869 76 876 128
rect 810 66 876 76
rect 0 59 876 66
rect 0 7 52 59
rect 104 50 116 59
rect 168 50 180 59
rect 232 50 244 59
rect 168 16 169 50
rect 232 16 241 50
rect 104 7 116 16
rect 168 7 180 16
rect 232 7 244 16
rect 296 7 308 59
rect 360 50 516 59
rect 360 16 385 50
rect 419 16 457 50
rect 491 16 516 50
rect 360 7 516 16
rect 568 7 580 59
rect 632 50 644 59
rect 696 50 708 59
rect 760 50 772 59
rect 635 16 644 50
rect 707 16 708 50
rect 632 7 644 16
rect 696 7 708 16
rect 760 7 772 16
rect 824 7 876 59
rect 0 0 876 7
<< via1 >>
rect 52 902 104 911
rect 116 902 168 911
rect 180 902 232 911
rect 244 902 296 911
rect 52 868 97 902
rect 97 868 104 902
rect 116 868 131 902
rect 131 868 168 902
rect 180 868 203 902
rect 203 868 232 902
rect 244 868 275 902
rect 275 868 296 902
rect 52 859 104 868
rect 116 859 168 868
rect 180 859 232 868
rect 244 859 296 868
rect 308 902 360 911
rect 516 902 568 911
rect 308 868 313 902
rect 313 868 347 902
rect 347 868 360 902
rect 516 868 529 902
rect 529 868 563 902
rect 563 868 568 902
rect 308 859 360 868
rect 516 859 568 868
rect 580 902 632 911
rect 644 902 696 911
rect 708 902 760 911
rect 772 902 824 911
rect 580 868 601 902
rect 601 868 632 902
rect 644 868 673 902
rect 673 868 696 902
rect 708 868 745 902
rect 745 868 760 902
rect 772 868 779 902
rect 779 868 824 902
rect 580 859 632 868
rect 644 859 696 868
rect 708 859 760 868
rect 772 859 824 868
rect 7 836 59 842
rect 7 802 16 836
rect 16 802 50 836
rect 50 802 59 836
rect 7 790 59 802
rect 7 764 59 778
rect 7 730 16 764
rect 16 730 50 764
rect 50 730 59 764
rect 7 726 59 730
rect 7 692 59 714
rect 7 662 16 692
rect 16 662 50 692
rect 50 662 59 692
rect 7 620 59 650
rect 7 598 16 620
rect 16 598 50 620
rect 50 598 59 620
rect 7 548 59 586
rect 7 534 16 548
rect 16 534 50 548
rect 50 534 59 548
rect 7 370 16 384
rect 16 370 50 384
rect 50 370 59 384
rect 7 332 59 370
rect 7 298 16 320
rect 16 298 50 320
rect 50 298 59 320
rect 7 268 59 298
rect 7 226 16 256
rect 16 226 50 256
rect 50 226 59 256
rect 7 204 59 226
rect 7 188 59 192
rect 7 154 16 188
rect 16 154 50 188
rect 50 154 59 188
rect 7 140 59 154
rect 7 116 59 128
rect 7 82 16 116
rect 16 82 50 116
rect 50 82 59 116
rect 7 76 59 82
rect 412 784 464 818
rect 412 766 421 784
rect 421 766 455 784
rect 455 766 464 784
rect 412 750 421 754
rect 421 750 455 754
rect 455 750 464 754
rect 412 712 464 750
rect 412 702 421 712
rect 421 702 455 712
rect 455 702 464 712
rect 412 678 421 690
rect 421 678 455 690
rect 455 678 464 690
rect 412 640 464 678
rect 412 638 421 640
rect 421 638 455 640
rect 455 638 464 640
rect 412 606 421 626
rect 421 606 455 626
rect 455 606 464 626
rect 412 574 464 606
rect 412 534 421 562
rect 421 534 455 562
rect 455 534 464 562
rect 412 510 464 534
rect 119 433 171 485
rect 183 433 235 485
rect 247 433 299 485
rect 311 433 363 485
rect 513 433 565 485
rect 577 433 629 485
rect 641 433 693 485
rect 705 433 757 485
rect 412 384 464 408
rect 412 356 421 384
rect 421 356 455 384
rect 455 356 464 384
rect 412 312 464 344
rect 412 292 421 312
rect 421 292 455 312
rect 455 292 464 312
rect 412 278 421 280
rect 421 278 455 280
rect 455 278 464 280
rect 412 240 464 278
rect 412 228 421 240
rect 421 228 455 240
rect 455 228 464 240
rect 412 206 421 216
rect 421 206 455 216
rect 455 206 464 216
rect 412 168 464 206
rect 412 164 421 168
rect 421 164 455 168
rect 455 164 464 168
rect 412 134 421 152
rect 421 134 455 152
rect 455 134 464 152
rect 412 100 464 134
rect 817 836 869 842
rect 817 802 826 836
rect 826 802 860 836
rect 860 802 869 836
rect 817 790 869 802
rect 817 764 869 778
rect 817 730 826 764
rect 826 730 860 764
rect 860 730 869 764
rect 817 726 869 730
rect 817 692 869 714
rect 817 662 826 692
rect 826 662 860 692
rect 860 662 869 692
rect 817 620 869 650
rect 817 598 826 620
rect 826 598 860 620
rect 860 598 869 620
rect 817 548 869 586
rect 817 534 826 548
rect 826 534 860 548
rect 860 534 869 548
rect 817 370 826 384
rect 826 370 860 384
rect 860 370 869 384
rect 817 332 869 370
rect 817 298 826 320
rect 826 298 860 320
rect 860 298 869 320
rect 817 268 869 298
rect 817 226 826 256
rect 826 226 860 256
rect 860 226 869 256
rect 817 204 869 226
rect 817 188 869 192
rect 817 154 826 188
rect 826 154 860 188
rect 860 154 869 188
rect 817 140 869 154
rect 817 116 869 128
rect 817 82 826 116
rect 826 82 860 116
rect 860 82 869 116
rect 817 76 869 82
rect 52 50 104 59
rect 116 50 168 59
rect 180 50 232 59
rect 244 50 296 59
rect 52 16 97 50
rect 97 16 104 50
rect 116 16 131 50
rect 131 16 168 50
rect 180 16 203 50
rect 203 16 232 50
rect 244 16 275 50
rect 275 16 296 50
rect 52 7 104 16
rect 116 7 168 16
rect 180 7 232 16
rect 244 7 296 16
rect 308 50 360 59
rect 516 50 568 59
rect 308 16 313 50
rect 313 16 347 50
rect 347 16 360 50
rect 516 16 529 50
rect 529 16 563 50
rect 563 16 568 50
rect 308 7 360 16
rect 516 7 568 16
rect 580 50 632 59
rect 644 50 696 59
rect 708 50 760 59
rect 772 50 824 59
rect 580 16 601 50
rect 601 16 632 50
rect 644 16 673 50
rect 673 16 696 50
rect 708 16 745 50
rect 745 16 760 50
rect 772 16 779 50
rect 779 16 824 50
rect 580 7 632 16
rect 644 7 696 16
rect 708 7 760 16
rect 772 7 824 16
<< metal2 >>
rect 0 911 383 918
rect 0 859 52 911
rect 104 859 116 911
rect 168 859 180 911
rect 232 859 244 911
rect 296 859 308 911
rect 360 859 383 911
rect 0 852 383 859
rect 0 842 66 852
rect 0 790 7 842
rect 59 790 66 842
rect 411 824 465 918
rect 493 911 876 918
rect 493 859 516 911
rect 568 859 580 911
rect 632 859 644 911
rect 696 859 708 911
rect 760 859 772 911
rect 824 859 876 911
rect 493 852 876 859
rect 810 842 876 852
rect 94 818 782 824
rect 94 796 412 818
rect 0 778 66 790
rect 0 726 7 778
rect 59 768 66 778
rect 59 740 383 768
rect 411 766 412 796
rect 464 796 782 818
rect 464 766 465 796
rect 810 790 817 842
rect 869 790 876 842
rect 810 778 876 790
rect 810 768 817 778
rect 411 754 465 766
rect 59 726 66 740
rect 0 714 66 726
rect 0 662 7 714
rect 59 662 66 714
rect 411 712 412 754
rect 94 702 412 712
rect 464 712 465 754
rect 493 740 817 768
rect 810 726 817 740
rect 869 726 876 778
rect 810 714 876 726
rect 464 702 782 712
rect 94 690 782 702
rect 94 684 412 690
rect 0 656 66 662
rect 0 650 383 656
rect 0 598 7 650
rect 59 628 383 650
rect 411 638 412 684
rect 464 684 782 690
rect 464 638 465 684
rect 810 662 817 714
rect 869 662 876 714
rect 810 656 876 662
rect 59 598 66 628
rect 411 626 465 638
rect 493 650 876 656
rect 493 628 817 650
rect 411 600 412 626
rect 0 586 66 598
rect 0 534 7 586
rect 59 544 66 586
rect 94 574 412 600
rect 464 600 465 626
rect 464 574 782 600
rect 94 572 782 574
rect 810 598 817 628
rect 869 598 876 650
rect 810 586 876 598
rect 411 562 465 572
rect 59 534 383 544
rect 0 516 383 534
rect 0 514 66 516
rect 411 510 412 562
rect 464 510 465 562
rect 810 544 817 586
rect 493 534 817 544
rect 869 534 876 586
rect 493 516 876 534
rect 810 514 876 516
rect 411 486 465 510
rect 0 485 876 486
rect 0 433 119 485
rect 171 433 183 485
rect 235 433 247 485
rect 299 433 311 485
rect 363 433 513 485
rect 565 433 577 485
rect 629 433 641 485
rect 693 433 705 485
rect 757 433 876 485
rect 0 432 876 433
rect 411 408 465 432
rect 0 402 66 404
rect 0 384 383 402
rect 0 332 7 384
rect 59 374 383 384
rect 59 332 66 374
rect 411 356 412 408
rect 464 356 465 408
rect 810 402 876 404
rect 493 384 876 402
rect 493 374 817 384
rect 411 346 465 356
rect 0 320 66 332
rect 0 268 7 320
rect 59 290 66 320
rect 94 344 782 346
rect 94 318 412 344
rect 411 292 412 318
rect 464 318 782 344
rect 810 332 817 374
rect 869 332 876 384
rect 810 320 876 332
rect 464 292 465 318
rect 59 268 383 290
rect 0 262 383 268
rect 411 280 465 292
rect 810 290 817 320
rect 0 256 66 262
rect 0 204 7 256
rect 59 204 66 256
rect 411 234 412 280
rect 94 228 412 234
rect 464 234 465 280
rect 493 268 817 290
rect 869 268 876 320
rect 493 262 876 268
rect 810 256 876 262
rect 464 228 782 234
rect 94 216 782 228
rect 94 206 412 216
rect 0 192 66 204
rect 0 140 7 192
rect 59 178 66 192
rect 59 150 383 178
rect 411 164 412 206
rect 464 206 782 216
rect 464 164 465 206
rect 810 204 817 256
rect 869 204 876 256
rect 810 192 876 204
rect 810 178 817 192
rect 411 152 465 164
rect 59 140 66 150
rect 0 128 66 140
rect 0 76 7 128
rect 59 76 66 128
rect 411 122 412 152
rect 94 100 412 122
rect 464 122 465 152
rect 493 150 817 178
rect 810 140 817 150
rect 869 140 876 192
rect 810 128 876 140
rect 464 100 782 122
rect 94 94 782 100
rect 0 66 66 76
rect 0 59 383 66
rect 0 7 52 59
rect 104 7 116 59
rect 168 7 180 59
rect 232 7 244 59
rect 296 7 308 59
rect 360 7 383 59
rect 0 0 383 7
rect 411 0 465 94
rect 810 76 817 128
rect 869 76 876 128
rect 810 66 876 76
rect 493 59 876 66
rect 493 7 516 59
rect 568 7 580 59
rect 632 7 644 59
rect 696 7 708 59
rect 760 7 772 59
rect 824 7 876 59
rect 493 0 876 7
<< metal3 >>
rect 0 0 876 918
<< labels >>
flabel metal3 s 634 62 728 149 0 FreeSans 200 0 0 0 MET3
port 4 nsew
flabel metal2 s 291 884 317 914 0 FreeSans 400 0 0 0 C0
port 1 nsew
flabel metal2 s 420 868 458 905 0 FreeSans 400 0 0 0 C1
port 2 nsew
flabel pwell s 467 350 491 401 0 FreeSans 200 0 0 0 SUB
port 3 nsew
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_END 117848
string GDS_START 100312
<< end >>
