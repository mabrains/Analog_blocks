* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre = 0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__pfet_01v8_hvt__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_hvt__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_hvt__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_hvt__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt  sky130_fd_pr__pfet_01v8_hvt d g s b
+ 
.param  l = 1 w = 1 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1 
msky130_fd_pr__pfet_01v8_hvt d g s b sky130_fd_pr__pfet_01v8_hvt__model l = {l} w = {w} nf = {nf} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd} 
.model sky130_fd_pr__pfet_01v8_hvt__model.0 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.116496+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43657182
+ k2 = 0.035761468
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.16745888+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.6448576+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.010851298
+ ua = 8.105303e-11
+ ub = 1.2961173e-19
+ uc = -7.7670696e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 200000.0
+ a0 = 1.5
+ ags = 0.3831138
+ a1 = 0.0
+ a2 = 1.0
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.013169082
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.075489662
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0036275994
+ pdiblcb = -9.5744039e-5
+ drout = 0.56
+ pscbe1 = 746475130.0
+ pscbe2 = 9.5049925e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.7923891
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1154444600.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.44169
+ kt2 = -0.037961
+ at = 0.0
+ ute = -0.30066
+ ua1 = 2.2116e-9
+ ub1 = -7.9359e-19
+ uc1 = 1.1985e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.1 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.116496+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43657182
+ k2 = 0.035761468
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.16745888+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.6448576+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.010851298
+ ua = 8.105303e-11
+ ub = 1.2961173e-19
+ uc = -7.7670696e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 200000.0
+ a0 = 1.5
+ ags = 0.3831138
+ a1 = 0.0
+ a2 = 1.0
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.013169082
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.075489662
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0036275994
+ pdiblcb = -9.5744039e-5
+ drout = 0.56
+ pscbe1 = 746475130.0
+ pscbe2 = 9.5049925e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.7923891
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1154444600.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.44169
+ kt2 = -0.037961
+ at = 0.0
+ ute = -0.30066
+ ua1 = 2.2116e-9
+ ub1 = -7.9359e-19
+ uc1 = 1.1985e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.2 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.115360748e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -9.148055522e-09 wvth0 = -1.134309093e-07 pvth0 = 9.140455501e-13
+ k1 = 4.360524374e-01 lk1 = 4.185273404e-09 wk1 = 5.189511220e-08 pk1 = -4.181796363e-13
+ k2 = 3.635591942e-02 lk2 = -4.790190628e-09 wk2 = -5.939575652e-08 pk2 = 4.786211033e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.687790987e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.063854708e-08 wvoff = 1.319121934e-07 pvoff = -1.062970879e-12
+ nfactor = {1.558907272e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.926023542e-07 wnfactor = 8.587892214e-06 pnfactor = -6.920269540e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.081580931e-02 lu0 = 2.859738705e-10 wu0 = 3.545920340e-09 pu0 = -2.857362891e-14
+ ua = 7.518714660e-11 lua = 4.726828563e-17 wua = 5.861010140e-16 pua = -4.722901608e-21
+ ub = 1.300649646e-19 lub = -3.652241838e-27 wub = -4.528581091e-26 pub = 3.649207629e-31
+ uc = -7.712339508e-11 luc = -4.410243821e-18 wuc = -5.468462292e-17 puc = 4.406579878e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.943948519e+05 lvsat = 4.516723660e-02 wvsat = 5.600491497e-01 pvsat = -4.512971257e-6
+ a0 = 1.522637133e+00 la0 = -1.824138688e-07 wa0 = -2.261832687e-06 pa0 = 1.822623230e-11
+ ags = 4.026310119e-01 lags = -1.572730118e-07 wags = -1.950099744e-06 pags = 1.571423525e-11
+ a1 = 0.0
+ a2 = 9.848993323e-01 la2 = 1.216031654e-07 wa2 = 1.507813064e-06 pa2 = -1.215021400e-11
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.635425645e-02 lketa = 2.566667719e-08 wketa = 3.182528269e-07 pketa = -2.564535382e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.175436333e-01 lpclm = -3.388780502e-07 wpclm = -4.201903374e-06 ppclm = 3.385965171e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 3.389944705e-03 lpdiblc2 = 1.915061933e-09 wpdiblc2 = 2.374572561e-08 ppdiblc2 = -1.913470938e-13
+ pdiblcb = -1.467027103e-04 lpdiblcb = 4.106336362e-10 wpdiblcb = 5.091633585e-09 ppdiblcb = -4.102924900e-14
+ drout = 0.56
+ pscbe1 = 7.505139621e+08 lpscbe1 = -3.254559539e+01 wpscbe1 = -4.035476685e+02 ppscbe1 = 3.251855716e-3
+ pscbe2 = 9.463158972e-09 lpscbe2 = 3.371016809e-16 wpscbe2 = 4.179877361e-15 ppscbe2 = -3.368216235e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.831931358e+00 lbeta0 = -3.186382355e-07 wbeta0 = -3.950940688e-06 pbeta0 = 3.183735172e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.034211168e-10 lagidl = -2.756794046e-17 wagidl = -3.418274567e-16 pagidl = 2.754503756e-21
+ bgidl = 1.142790657e+09 lbgidl = 9.390945669e+01 wbgidl = 1.164426149e+03 pbgidl = -9.383143859e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.425026731e-01 lkt1 = 6.548657891e-09 wkt1 = 8.119979347e-08 pkt1 = -6.543217397e-13
+ kt2 = -3.814096521e-02 lkt2 = 1.450190257e-09 wkt2 = 1.798156986e-08 pkt2 = -1.448985468e-13
+ at = 1.980824625e+04 lat = -1.596182157e-01 wat = -1.979178996e+00 pat = 1.594856081e-5
+ ute = -3.004781484e-01 lute = -1.465391413e-09 wute = -1.817005592e-08 pute = 1.464173995e-13
+ ua1 = 2.227204531e-09 lua1 = -1.257439603e-16 wua1 = -1.559156666e-15 pua1 = 1.256394947e-20
+ ub1 = -8.067368925e-19 lub1 = 1.059398946e-25 wub1 = 1.313597030e-24 pub1 = -1.058518818e-29
+ uc1 = 1.211380529e-10 luc1 = -1.037934914e-17 wuc1 = -1.286982799e-16 puc1 = 1.037072618e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.3 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.132529876e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.052718416e-08 wvth0 = 5.508338126e-08 pvth0 = 2.301859117e-13
+ k1 = 4.496812128e-01 lk1 = -5.112261417e-08 wk1 = -6.021040076e-07 pk1 = 2.235859972e-12
+ k2 = 2.473168602e-02 lk2 = 4.238292463e-08 wk2 = 2.920218154e-07 pk2 = -9.474911443e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 5.439684414e-01 ldsub = 6.505878998e-08 wdsub = 1.601823986e-06 pdsub = -6.500474044e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.439825003e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.999026487e-08 wvoff = -5.466675025e-07 pvoff = 1.690820885e-12
+ nfactor = {3.089221135e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.517671454e-06 wnfactor = -2.719458015e-05 pnfactor = 7.600866048e-11
+ eta0 = 7.391517200e-02 leta0 = 2.469326643e-08 weta0 = 6.079772844e-07 peta0 = -2.467275176e-12
+ etab = -6.468055917e-02 letab = -2.158719519e-08 wetab = -5.315021543e-07 petab = 2.156926098e-12
+ u0 = 1.121725328e-02 lu0 = -1.343153981e-09 wu0 = 1.179417985e-08 pu0 = -6.204646819e-14
+ ua = 1.389910308e-10 lua = -2.116587233e-16 wua = 2.204266048e-15 pua = -1.128969041e-20
+ ub = 1.332488489e-19 lub = -1.657298547e-26 wub = -9.810181673e-25 pub = 4.162281739e-30
+ uc = -8.641091460e-11 luc = 3.328008923e-17 wuc = 1.275061871e-16 puc = -2.987032917e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.823927283e+05 lvsat = -3.119431056e-01 wvsat = -5.944706893e-01 pvsat = 1.722665183e-7
+ a0 = 1.148626736e+00 la0 = 1.335383906e-06 wa0 = 4.261233318e-06 pa0 = -8.245478465e-12
+ ags = 8.410057061e-02 lags = 1.135377669e-06 wags = 3.280997489e-06 pags = -5.514446606e-12
+ a1 = 0.0
+ a2 = 1.235978044e+00 la2 = -8.973169318e-07 wa2 = -3.015626127e-06 pa2 = 6.206671226e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = 3.646406548e-02 lketa = -1.886790523e-07 wketa = -6.188554003e-07 pketa = 1.238409112e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.839671156e-01 lpclm = 2.507971826e-06 wpclm = 8.585282079e-06 ppclm = -1.803292068e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 7.326120933e-03 lpdiblc2 = -1.405861035e-08 wpdiblc2 = -4.570039274e-08 ppdiblc2 = 9.047706036e-14
+ pdiblcb = 6.423123938e-04 lpdiblcb = -2.791323789e-09 wpdiblcb = -4.304566255e-09 ppdiblcb = -2.897872699e-15
+ drout = 0.56
+ pscbe1 = 6.833158250e+08 lpscbe1 = 2.401558684e+02 wpscbe1 = 8.070953369e+02 ppscbe1 = -1.661139410e-3
+ pscbe2 = 1.013790104e-08 lpscbe2 = -2.401116331e-15 wpscbe2 = -6.233054770e-15 ppscbe2 = 8.575286431e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.325229279e+00 lbeta0 = 1.737644938e-06 wbeta0 = -7.205805815e-06 pbeta0 = 4.504614774e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 4.343435213e-11 lagidl = 2.158685482e-16 wagidl = 9.900184142e-16 pagidl = -2.650353201e-21
+ bgidl = 1.336689108e+09 lbgidl = -6.929634212e+02 wbgidl = -2.328852298e+03 pbgidl = 4.793173933e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.273136297e-01 lkt1 = -5.509106218e-08 wkt1 = -3.290388955e-07 pkt1 = 1.010496601e-12
+ kt2 = -3.540295348e-02 lkt2 = -9.661126809e-09 wkt2 = -1.035926616e-08 pkt2 = -2.988661629e-14
+ at = -3.228964051e+05 lat = 1.231135519e+00 wat = 5.270747699e+00 pat = -1.347287421e-5
+ ute = -2.934284710e-01 lute = -3.007418042e-08 wute = -9.703555585e-07 pute = 4.010548040e-12
+ ua1 = 1.922938781e-09 lua1 = 1.109018176e-15 wua1 = 7.578342920e-15 pua1 = -2.451757722e-20
+ ub1 = -5.626399278e-19 lub1 = -8.846470846e-25 wub1 = -5.160968071e-24 pub1 = 1.568969768e-29
+ uc1 = 8.369283483e-11 luc1 = 1.415797114e-16 wuc1 = 1.857523945e-15 puc1 = -7.023354827e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.4 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.103201497e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.643954793e-10 wvth0 = 1.749042911e-07 pvth0 = -1.642589028e-14
+ k1 = 4.208874299e-01 lk1 = 8.139886086e-09 wk1 = 8.793928245e-07 pk1 = -8.133123631e-13
+ k2 = 4.611168922e-02 lk2 = -1.620756548e-09 wk2 = -2.470163350e-07 pk2 = 1.619410056e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 6.266919657e-01 ldsub = -1.052002859e-07 wdsub = -6.663655931e-06 pdsub = 1.051128876e-11
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.889773804e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.616847530e-09 wvoff = 4.018878820e-07 pvoff = -2.614673506e-13
+ nfactor = {3.855746458e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.689264014e-08 wnfactor = 1.201210771e-05 pnfactor = -4.685368267e-12
+ eta0 = 1.031707210e-01 leta0 = -3.551962676e-08 weta0 = -2.315147119e-06 peta0 = 3.549011777e-12
+ etab = -7.520844859e-02 letab = 8.099097412e-11 wetab = 5.204121513e-07 petab = -8.092368843e-15
+ u0 = 1.055098535e-02 lu0 = 2.813867794e-11 wu0 = -1.698621152e-08 pu0 = -2.811530089e-15
+ ua = 3.221364741e-11 lua = 8.107283979e-18 wua = -2.887458904e-15 pua = -8.100548610e-22
+ ub = 1.240130477e-19 lub = 2.435863480e-27 wub = 1.159556091e-24 pub = -2.433839813e-31
+ uc = -6.954668686e-11 luc = -1.429358354e-18 wuc = -8.701466337e-17 puc = 1.428170872e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.333293373e+05 lvsat = -5.145306209e-03 wvsat = -7.605583501e-01 pvsat = 5.141031592e-7
+ a0 = 1.794488058e+00 la0 = 6.091509343e-09 wa0 = 5.507363225e-07 pa0 = -6.086448639e-13
+ ags = 6.501711252e-01 lags = -2.969176410e-08 wags = -8.397293135e-07 pags = 2.966709677e-12
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.396872968e-02 lketa = -2.552986309e-09 wketa = -1.410899202e-07 pketa = 2.550865339e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.434649028e-01 lpclm = -1.829193137e-08 wpclm = -1.064355297e-06 ppclm = 1.827673480e-12
+ pdiblc1 = 3.864232508e-01 lpdiblc1 = 7.361557965e-09 wpdiblc1 = 3.573777739e-07 ppdiblc1 = -7.355442130e-13
+ pdiblc2 = 5.101340302e-04 lpdiblc2 = -3.015058607e-11 wpdiblc2 = -3.204142866e-09 ppdiblc2 = 3.012553756e-15
+ pdiblcb = -6.981996316e-04 lpdiblcb = -3.232215332e-11 wpdiblcb = -7.281678336e-09 ppdiblcb = 3.229530072e-15
+ drout = 5.827770016e-01 ldrout = -4.687894133e-08 wdrout = -2.275807889e-06 pdrout = 4.683999524e-12
+ pscbe1 = 800000000.0
+ pscbe2 = 9.005251489e-09 lpscbe2 = -6.993100867e-17 wpscbe2 = -5.461497857e-15 ppscbe2 = 6.987291139e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.289121979e+00 lbeta0 = -2.462100992e-07 wbeta0 = 2.728063817e-06 pbeta0 = 2.460055528e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.479026926e-10 lagidl = 8.549439624e-19 wagidl = -2.562002325e-16 pagidl = -8.542336921e-23
+ bgidl = 1.009958714e+09 lbgidl = -2.049672598e+01 wbgidl = -9.950440300e+02 pbgidl = 2.047969771e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.572450839e-01 lkt1 = 6.512958836e-09 wkt1 = 4.781108543e-07 pkt1 = -6.507548000e-13
+ kt2 = -4.037183061e-02 lkt2 = 5.656670423e-10 wkt2 = 2.580915386e-09 pkt2 = -5.651970974e-14
+ at = 2.796425669e+05 lat = -8.992116851e-03 wat = -1.711833354e+00 pat = 8.984646380e-7
+ ute = -4.059469952e-01 lute = 2.015080705e-07 wute = 1.076075227e-05 pute = -2.013406616e-11
+ ua1 = 2.266584461e-09 lua1 = 4.017369469e-16 wua1 = 1.516894135e-14 pua1 = -4.014031919e-20
+ ub1 = -8.822147098e-19 lub1 = -2.269078556e-25 wub1 = -8.553417108e-24 pub1 = 2.267193451e-29
+ uc1 = 1.581544240e-10 luc1 = -1.167489752e-17 wuc1 = -2.121678284e-15 puc1 = 1.166519825e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.5 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.130201236e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.873470962e-08 wvth0 = 3.671954291e-07 pvth0 = -2.199026038e-13
+ k1 = 3.533184844e-01 lk1 = 7.963931708e-08 wk1 = 3.626188190e-07 pk1 = -2.664776137e-13
+ k2 = 7.060629685e-02 lk2 = -2.754021550e-08 wk2 = -1.678265423e-07 pk2 = 7.814474258e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 7.784906946e-01 ldsub = -2.658291468e-07 wdsub = 1.532162588e-06 pdsub = 1.838719474e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.339405975e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.019557501e-08 wvoff = 7.691229931e-07 pvoff = -6.500645281e-13
+ nfactor = {-1.259055108e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.787190507e-06 wnfactor = 3.021132865e-05 pnfactor = -2.394323789e-11
+ eta0 = 1.478831241e-01 leta0 = -8.283295043e-08 weta0 = 2.084857089e-06 peta0 = -1.106940676e-12
+ etab = -1.584880103e-01 letab = 8.820492480e-08 wetab = 1.089332283e-06 petab = -6.101065849e-13
+ u0 = 1.338909091e-02 lu0 = -2.975059477e-09 wu0 = -2.510274429e-08 pu0 = 5.777141389e-15
+ ua = 4.819278446e-10 lua = -4.677667881e-16 wua = 1.425276021e-15 pua = -5.373661577e-21
+ ub = 5.487368492e-20 lub = 7.559706301e-26 wub = -7.561708063e-24 pub = 8.985196109e-30
+ uc = -6.397830380e-11 luc = -7.321654260e-18 wuc = -3.788576651e-16 puc = 4.516365963e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.156700469e+05 lvsat = -9.227577482e-02 wvsat = -1.321353239e+00 pvsat = 1.107519487e-6
+ a0 = 1.674995242e+00 la0 = 1.325352221e-07 wa0 = 8.662440896e-06 pa0 = -9.192207292e-12
+ ags = 5.274185762e-01 lags = 1.002013008e-07 wags = 2.394081854e-06 pags = -4.552122862e-13
+ a1 = 0.0
+ a2 = 8.166048401e-01 la2 = -1.757074360e-08 wa2 = -1.659104508e-06 pa2 = 1.755614617e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.268609813e-02 lketa = -3.910228537e-09 wketa = -1.181230786e-08 pketa = 1.182888429e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.685166376e-01 lpclm = -4.480092566e-08 wpclm = -9.205757449e-07 ppclm = 1.675530271e-12
+ pdiblc1 = 3.694046322e-01 lpdiblc1 = 2.537014953e-08 wpdiblc1 = 2.057825754e-06 ppdiblc1 = -2.534907252e-12
+ pdiblc2 = 7.913161930e-04 lpdiblc2 = -3.276891153e-10 wpdiblc2 = -5.175877274e-09 ppdiblc2 = 5.098983955e-15
+ pdiblcb = -1.771212109e-03 lpdiblcb = 1.103107460e-09 wpdiblcb = 1.856730307e-07 ppdiblcb = -2.009493544e-13
+ drout = 5.470954930e-01 ldrout = -9.121839370e-09 wdrout = 1.289378622e-06 pdrout = 9.114261128e-13
+ pscbe1 = 7.965929773e+08 lpscbe1 = 3.605209258e+00 wpscbe1 = 3.404192259e+02 ppscbe1 = -3.602214123e-4
+ pscbe2 = 9.275287906e-09 lpscbe2 = -3.556754440e-16 wpscbe2 = -1.424152772e-15 ppscbe2 = 2.715093690e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 2.708515230e+00 lbeta0 = 2.484510544e-06 wbeta0 = 4.022422636e-05 pbeta0 = -1.507675904e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.967579821e-10 lagidl = -5.084225782e-17 wagidl = -6.692674153e-16 pagidl = 3.516719316e-22
+ bgidl = 9.941236796e+08 lbgidl = -3.740567857e+00 wbgidl = 5.871438457e+02 pbgidl = 3.737460268e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.788433526e-01 lkt1 = 2.936759880e-08 wkt1 = 2.056593969e-07 pkt1 = -3.624548413e-13
+ kt2 = -3.461611266e-02 lkt2 = -5.524861026e-09 wkt2 = -1.990725791e-07 pkt2 = 1.568639686e-13
+ at = 4.681330673e+05 lat = -2.084471096e-01 wat = -1.403628914e+00 pat = 5.723319454e-7
+ ute = -2.654084824e-01 lute = 5.279443236e-08 wute = -1.796437976e-05 pute = 1.026200680e-11
+ ua1 = 3.612348718e-09 lua1 = -1.022310417e-15 wua1 = -5.424482002e-14 pua1 = 3.331124068e-20
+ ub1 = -1.730531725e-18 lub1 = 6.707557602e-25 wub1 = 3.925195874e-23 pub1 = -2.791428005e-29
+ uc1 = 3.818732144e-10 luc1 = -2.484074100e-16 wuc1 = -1.136636370e-15 puc1 = 1.241780216e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.6 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.077008961e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -9.556226842e-10 wvth0 = -1.978393828e-07 pvth0 = 9.548287719e-14
+ k1 = 5.205488237e-01 lk1 = -1.370364137e-08 wk1 = -2.567856268e-06 pk1 = 1.369225666e-12
+ k2 = 1.286083107e-02 lk2 = 4.691571130e-09 wk2 = 8.120041352e-07 pk2 = -4.687673467e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.732240609e-01 ldsub = 1.619553008e-08 wdsub = 7.725485392e-06 pdsub = -1.618207516e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.425720739e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.035938263e-10 wvoff = -5.393621454e-07 pvoff = 8.029262166e-14
+ nfactor = {2.093351763e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -8.402243660e-08 wnfactor = -2.772532351e-05 pnfactor = 8.395263244e-12
+ eta0 = 4.310549828e-02 leta0 = -2.434922301e-08 weta0 = -4.257010248e-06 peta0 = 2.432899416e-12
+ etab = -4.284317981e-04 letab = -1.919013535e-11 wetab = -7.150874450e-09 petab = 1.917419257e-15
+ u0 = 7.945281863e-03 lu0 = 6.351141609e-11 wu0 = -3.383542976e-09 pu0 = -6.345865208e-15
+ ua = -3.820568015e-10 lua = 1.448352182e-17 wua = -5.609341850e-15 pua = -1.447148920e-21
+ ub = 2.093582575e-19 lub = -1.063159085e-26 wub = 6.632749315e-24 pub = 1.062275834e-30
+ uc = -7.572867432e-11 luc = -7.629499476e-19 wuc = 2.937062239e-16 puc = 7.623161041e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.443328253e+04 lvsat = 3.303449926e-03 wvsat = 1.254188326e+00 pvsat = -3.300705486e-7
+ a0 = 1.912262443e+00 la0 = 9.978870383e-11 wa0 = -7.788168617e-06 pa0 = -9.970580137e-15
+ ags = 8.326356145e-01 lags = -7.016169353e-08 wags = -1.098097009e-05 pags = 7.010340460e-12
+ a1 = 0.0
+ a2 = 7.667903199e-01 la2 = 1.023422712e-08 wa2 = 3.318209016e-06 pa2 = -1.022572473e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = -6.489334968e-02 lketa = 2.903493065e-09 wketa = 7.198589268e-07 pketa = -2.901080901e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.729441980e-01 lpclm = 8.544742953e-09 wpclm = 3.610829896e-06 ppclm = -8.537644151e-13
+ pdiblc1 = 4.441053545e-01 lpdiblc1 = -1.632555261e-08 wpdiblc1 = -5.406040486e-06 ppdiblc1 = 1.631198967e-12
+ pdiblc2 = 9.096376623e-04 lpdiblc2 = -3.937326098e-10 wpdiblc2 = -6.652200213e-08 ppdiblc2 = 3.934055046e-14
+ pdiblcb = 2.050808841e-04 wpdiblcb = -1.743415785e-7
+ drout = 4.948982534e-01 ldrout = 2.001309381e-08 wdrout = 6.504766132e-06 pdrout = -1.999646734e-12
+ pscbe1 = 8.068140455e+08 lpscbe1 = -2.099884399e+00 wpscbe1 = -6.808384518e+02 ppscbe1 = 2.098139857e-4
+ pscbe2 = 7.892205808e-09 lpscbe2 = 4.163194907e-16 wpscbe2 = 7.796466385e-14 ppscbe2 = -4.159736208e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.537641680e-09 lalpha0 = -8.024484566e-16 walpha0 = -1.436447316e-13 palpha0 = 8.017817985e-20
+ alpha1 = 9.083188020e-11 lalpha1 = 5.117369427e-18 walpha1 = 9.160503106e-16 palpha1 = -5.113118019e-22
+ beta0 = 7.854541554e+00 lbeta0 = -3.878469692e-07 wbeta0 = -5.621455468e-05 pbeta0 = 3.875247537e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.056705754e-10 wagidl = -3.922292777e-17
+ bgidl = 9.941315072e+08 lbgidl = -3.744937003e+00 wbgidl = 5.863617334e+02 pbgidl = 3.741825784e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.268261322e-01 lkt1 = 3.331468905e-10 wkt1 = -3.840674415e-07 pkt1 = -3.328701188e-14
+ kt2 = -4.503746506e-02 lkt2 = 2.920252450e-10 wkt2 = 1.342348938e-07 pkt2 = -2.917826363e-14
+ at = 9.517042695e+04 lat = -2.705526606e-04 wat = -4.266879165e-01 pat = 2.703278908e-8
+ ute = -1.653227486e-01 lute = -3.070421656e-09 wute = -1.289179477e-07 pute = 3.067870811e-13
+ ua1 = 1.655805886e-09 lua1 = 6.977309585e-17 wua1 = 1.792450770e-14 pua1 = -6.971512975e-21
+ ub1 = -4.058556370e-19 lub1 = -6.863869172e-26 wub1 = -2.304527482e-23 pub1 = 6.858166807e-30
+ uc1 = -5.205499622e-11 luc1 = -6.201700656e-18 wuc1 = -2.024317218e-15 puc1 = 6.196548407e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.7 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.077206619e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -8.947104565e-10 wvth0 = -1.780900162e-07 pvth0 = 8.939671489e-14
+ k1 = 5.360338431e-01 lk1 = -1.847565980e-08 wk1 = -4.115071744e-06 pk1 = 1.846031059e-12
+ k2 = 2.692534619e-03 lk2 = 7.825135048e-09 wk2 = 1.827989019e-06 pk2 = -7.818634082e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.957845953e-01 ldsub = 9.243050194e-09 wdsub = 5.471306236e-06 pdsub = -9.235371252e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.541898097e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.776643818e-09 wvoff = 6.214462572e-07 pvoff = -2.774337038e-13
+ nfactor = {1.787411401e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.025920464e-08 wnfactor = 2.843295737e-06 pnfactor = -1.025068149e-12
+ eta0 = -3.590680988e-02 weta0 = 3.637656383e-6
+ etab = -4.907030694e-04 letab = 2.339540454e-18 wetab = -9.289206876e-10 petab = -2.337596809e-22
+ u0 = 7.882086830e-03 lu0 = 8.298622943e-11 wu0 = 2.930710213e-09 pu0 = -8.291728613e-15
+ ua = -4.512945434e-10 lua = 3.582051675e-17 wua = 1.308680213e-15 pua = -3.579075779e-21
+ ub = 2.781685427e-19 lub = -3.183685644e-26 wub = -2.425625849e-25 pub = 3.181040702e-30
+ uc = -8.097796026e-11 luc = 8.547224992e-19 wuc = 8.181987173e-16 puc = -8.540124129e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.123500318e+04 lvsat = -1.874336327e-03 wvsat = -4.245878856e-01 pvsat = 1.872779166e-7
+ a0 = 1.867795103e+00 la0 = 1.380328869e-08 wa0 = -3.345128934e-06 pa0 = -1.379182119e-12
+ ags = 3.376844041e-01 lags = 8.236742098e-08 wags = 3.847303139e-05 pags = -8.229899177e-12
+ a1 = 0.0
+ a2 = 7.809164901e-01 la2 = 5.880965231e-09 wa2 = 1.906765565e-06 pa2 = -5.876079443e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.565306657e-02 lketa = 5.591501689e-11 wketa = -2.034017208e-07 pketa = -5.586856381e-15
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.958722954e-01 lpclm = 1.478991189e-09 wpclm = 1.319924980e-06 ppclm = -1.477762473e-13
+ pdiblc1 = 3.994217871e-01 lpdiblc1 = -2.555417652e-09 wpdiblc1 = -9.413959688e-07 ppdiblc1 = 2.553294662e-13
+ pdiblc2 = -1.994982030e-04 lpdiblc2 = -5.193021021e-11 wpdiblc2 = 4.429943961e-08 ppdiblc2 = 5.188706763e-15
+ pdiblcb = -3.785228148e-02 lpdiblcb = 1.172813736e-08 wpdiblcb = 3.628232929e-06 ppdiblcb = -1.171839386e-12
+ drout = 5.656434769e-01 ldrout = -1.788461701e-09 wdrout = -5.638788429e-07 pdrout = 1.786975883e-13
+ pscbe1 = 7.999741224e+08 lpscbe1 = 7.974713567e-03 wpscbe1 = 2.585614542e+00 ppscbe1 = -7.968088334e-7
+ pscbe2 = 1.133901833e-08 lpscbe2 = -6.458847243e-16 wpscbe2 = -2.664302341e-13 ppscbe2 = 6.453481362e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.387406033e-09 lalpha0 = 9.896349709e-17 walpha0 = 1.486170326e-13 palpha0 = -9.888128020e-21
+ alpha1 = 1.074375505e-10 walpha1 = -7.431371569e-16
+ beta0 = 6.478528643e+00 lbeta0 = 3.619892962e-08 wbeta0 = 8.127242003e-05 pbeta0 = -3.616885628e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.056705754e-10 wagidl = -3.922292777e-17
+ bgidl = 1.021194081e+09 lbgidl = -1.208481044e+01 wbgidl = -2.117647365e+03 pbgidl = 1.207477062e-3
+ cgidl = 2.364927263e+02 lcgidl = 1.957103654e-05 wcgidl = 6.345451314e-03 pcgidl = -1.955477731e-9
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.310094553e-01 lkt1 = 1.622321575e-09 wkt1 = 3.391732802e-08 pkt1 = -1.620973783e-13
+ kt2 = -4.781343434e-02 lkt2 = 1.147495697e-09 wkt2 = 4.116011995e-07 pkt2 = -1.146542381e-13
+ at = 9.119027697e+04 lat = 9.560101597e-04 wat = -2.900358106e-02 pat = -9.552159256e-8
+ ute = -2.048786767e-01 lute = 9.119528696e-09 wute = 3.823388632e-06 pute = -9.111952374e-13
+ ua1 = 1.673334884e-09 lua1 = 6.437118449e-17 wua1 = 1.617306416e-14 pua1 = -6.431770620e-21
+ ub1 = -4.227640831e-19 lub1 = -6.342801591e-26 wub1 = -2.135583494e-23 pub1 = 6.337532118e-30
+ uc1 = -5.578544392e-11 luc1 = -5.052088585e-18 wuc1 = -1.651582365e-15 puc1 = 5.047891411e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.8 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -3.7585e-8
+ vth0 = {-1.086845933e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.501090964e-09 wvth0 = 7.850405458e-07 pvth0 = -1.499843888e-13
+ k1 = 5.132569025e-01 lk1 = -1.398241590e-08 wk1 = -1.839269952e-06 pk1 = 1.397079959e-12
+ k2 = 3.355576240e-03 lk2 = 8.214485978e-09 wk2 = 1.761739941e-06 pk2 = -8.207661548e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.918248643e-01 ldsub = 3.643020139e-08 wdsub = 1.585864257e-05 pdsub = -3.639993590e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.483561967e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.486270931e-09 wvoff = 3.856960449e-08 pvoff = -1.485036167e-13
+ nfactor = {2.035507946e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.231531347e-08 wnfactor = -2.194574740e-05 pnfactor = 5.227185096e-12
+ eta0 = -1.866310028e-01 leta0 = 3.846029230e-08 weta0 = 1.869755381e-05 peta0 = -3.842834026e-12
+ etab = -2.015693448e-02 letab = 5.018232271e-09 wetab = 1.964060389e-06 petab = -5.014063224e-13
+ u0 = 8.895933403e-03 lu0 = -1.697936438e-10 wu0 = -9.836971876e-08 pu0 = 1.696525826e-14
+ ua = -9.187340890e-11 lua = -5.333619208e-17 wua = -3.460357325e-14 pua = 5.329188143e-21
+ ub = -4.080572035e-20 lub = 4.728336825e-26 wub = 3.162836398e-23 pub = -4.724408617e-30
+ uc = -7.966082027e-11 luc = 5.796359200e-19 wuc = 6.865941445e-16 puc = -5.791543701e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.858955382e+04 lvsat = 6.322017382e-03 wvsat = 2.837244932e+00 pvsat = -6.316765176e-7
+ a0 = 1.919085359e+00 la0 = 1.700799593e-09 wa0 = -8.469893410e-06 pa0 = -1.699386603e-13
+ ags = 6.835189802e-01 wags = 3.918305029e-6
+ a1 = 0.0
+ a2 = 8.386837579e-01 la2 = -8.439739363e-09 wa2 = -3.865162018e-06 pa2 = 8.432727797e-13
+ b0 = 1.176374414e-24 lb0 = -3.001754592e-31 wb0 = -1.175397105e-28 pb0 = 2.999260794e-35
+ b1 = 0.0
+ keta = -1.828432198e-02 lketa = -9.475476460e-09 wketa = -3.937171659e-06 pketa = 9.467604423e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.600215177e-01 lpclm = 1.073260097e-08 wpclm = 4.902024344e-06 ppclm = -1.072368454e-12
+ pdiblc1 = 2.608638392e-01 lpdiblc1 = 3.261801436e-08 wpdiblc1 = 1.290288770e-05 ppdiblc1 = -3.259091597e-12
+ pdiblc2 = -3.365133103e-03 lpdiblc2 = 7.521381940e-10 wpdiblc2 = 3.605999349e-07 ppdiblc2 = -7.515133326e-14
+ pdiblcb = 1.509728261e-02 lpdiblcb = -9.458767599e-10 wpdiblcb = -1.662324537e-06 ppdiblcb = 9.450909444e-14
+ drout = 7.897555514e-01 ldrout = -5.910279583e-08 wdrout = -2.295646751e-05 pdrout = 5.905369441e-12
+ pscbe1 = 8.000646910e+08 lpscbe1 = -1.456647960e-02 wpscbe1 = -6.463728763e+00 ppscbe1 = 1.455437806e-6
+ pscbe2 = 8.757038745e-09 lpscbe2 = -3.314268682e-17 wpscbe2 = -8.446781241e-15 ppscbe2 = 3.311515254e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.927823646e-09 lalpha0 = 1.264605635e-15 walpha0 = 6.022815850e-13 palpha0 = -1.263555026e-19
+ alpha1 = 1.074375505e-10 walpha1 = -7.431371569e-16
+ beta0 = 5.325728347e+00 lbeta0 = 3.329427735e-07 wbeta0 = 1.964566773e-04 pbeta0 = -3.326661713e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.056705754e-10 wagidl = -3.922292777e-17
+ bgidl = 9.073455903e+08 lbgidl = 1.610332439e+01 wbgidl = 9.257743428e+03 pbgidl = -1.608994607e-3
+ cgidl = 4.587606293e+02 lcgidl = -3.574813089e-05 wcgidl = -1.586287341e-02 pcgidl = 3.571843206e-9
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -2.8385e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.302547231e-01 lkt1 = 1.545533969e-09 wkt1 = -4.149318701e-08 pkt1 = -1.544249970e-13
+ kt2 = -3.601302746e-02 lkt2 = -1.781708652e-09 wkt2 = -7.674591344e-07 pkt2 = 1.780228444e-13
+ at = 9.060605489e+04 lat = 1.173323806e-03 wat = 2.937009084e-02 pat = -1.172349032e-7
+ ute = -2.297030394e-01 lute = 1.610489129e-08 wute = 6.303762545e-06 pute = -1.609151167e-12
+ ua1 = 1.963303621e-09 lua1 = -5.025478195e-18 wua1 = -1.279971948e-14 pua1 = 5.021303128e-22
+ ub1 = -7.516381574e-19 lub1 = 1.596344288e-26 wub1 = 1.150425029e-23 pub1 = -1.595018077e-30
+ uc1 = -9.220523568e-11 luc1 = 3.880543782e-18 wuc1 = 1.987371127e-15 puc1 = -3.877319904e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.9 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.101588297e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.491637494e-06 wvth0 = -1.031154198e-07 pvth0 = 1.031754020e-11
+ k1 = 4.350967556e-01 lk1 = 1.475922413e-07 wk1 = 1.020290518e-08 pk1 = -1.020884021e-12
+ k2 = 3.938115510e-02 lk2 = -3.621792668e-07 wk2 = -2.503709330e-08 pk2 = 2.505165738e-12
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.662142270e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.245376994e-07 wvoff = -8.609167579e-09 pvoff = 8.614175531e-13
+ nfactor = {1.448509620e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.964621959e-05 wnfactor = 1.358123665e-06 pnfactor = -1.358913685e-10
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 9.894386806e-03 lu0 = 9.574678295e-08 wu0 = 6.618880092e-09 pu0 = -6.622730294e-13
+ ua = -3.186148866e-11 lua = 1.129802010e-14 wua = 7.810209182e-16 pua = -7.814752381e-20
+ ub = 1.225188563e-19 lub = 7.096999649e-25 wub = 4.906085430e-26 pub = -4.908939300e-30
+ uc = -7.883333226e-11 luc = 1.163312570e-16 wuc = 8.041864357e-18 puc = -8.046542310e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.755365116e+05 lvsat = 2.447771886e+00 wvsat = 1.692120414e-01 pvsat = -1.693104721e-5
+ a0 = 1.626458128e+00 la0 = -1.265316891e-05 wa0 = -8.747010106e-07 pa0 = 8.752098242e-11
+ ags = 4.281320677e-01 lags = -4.504445487e-06 wags = -3.113878465e-07 pags = 3.115689808e-11
+ a1 = 0.0
+ a2 = 8.767155923e-01 la2 = 1.233461164e-05 wa2 = 8.526794624e-07 pa2 = -8.531754660e-11
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.592827572e-02 lketa = 2.277243274e-06 wketa = 1.574235677e-07 pketa = -1.575151410e-11
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.371115655e-01 lpclm = -6.165774894e-06 wpclm = -4.262338999e-07 ppclm = 4.264818401e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 1.494098405e-03 lpdiblc2 = 2.134742053e-07 wpdiblc2 = 1.475725997e-08 ppdiblc2 = -1.476584427e-12
+ pdiblcb = -1.926174062e-03 lpdiblcb = 1.831494784e-07 wpdiblcb = 1.266094170e-08 ppdiblcb = -1.266830657e-12
+ drout = 0.56
+ pscbe1 = 7.293810089e+08 lpscbe1 = 1.710406471e+03 wpscbe1 = 1.182387020e+02 ppscbe1 = -1.183074814e-2
+ pscbe2 = 9.566587049e-09 lpscbe2 = -6.163037830e-15 wpscbe2 = -4.260446894e-16 ppscbe2 = 4.262925195e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.308721188e-10 lalpha0 = -2.310064171e-14 walpha0 = -1.596924438e-15 palpha0 = 1.597853369e-19
+ alpha1 = 3.852939096e-11 lalpha1 = 6.150636650e-15 walpha1 = 4.251874080e-16 palpha1 = -4.254347396e-20
+ beta0 = 3.819947759e+00 lbeta0 = 9.730070102e-05 wbeta0 = 6.726300906e-06 pbeta0 = -6.730213595e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.336878087e+09 lbgidl = -1.825396086e+04 wbgidl = -1.261878200e+03 pbgidl = 1.262612235e-1
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.355259714e-01 lkt1 = -6.167614200e-07 wkt1 = -4.263610493e-08 pkt1 = 4.266090635e-12
+ kt2 = -0.037961
+ at = 0.0
+ ute = -3.315232911e-01 lute = 3.088124430e-06 wute = 2.134789774e-07 pute = -2.136031581e-11
+ ua1 = 2.2116e-9
+ ub1 = -8.718546709e-19 lub1 = 7.831019750e-24 wub1 = 5.413506242e-25 pub1 = -5.416655279e-29
+ uc1 = 1.1985e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.10 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.175953879e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 4.112655133e-7
+ k1 = 4.424549663e-01 wk1 = -4.069326436e-8
+ k2 = 2.132470893e-02 wk2 = 9.985793641e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.724230536e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} wvoff = 3.433680173e-8
+ nfactor = {2.427971833e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = -5.416740070e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.466784236e-02 wu0 = -2.639873963e-8
+ ua = 5.314012668e-10 wua = -3.115023627e-15
+ ub = 1.579009457e-19 wub = -1.956742985e-25
+ uc = -7.303363782e-11 wuc = -3.207416971e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.975701709e+05 wvsat = -6.748852619e-1
+ a0 = 9.956344335e-01 wa0 = 3.488657283e-6
+ ags = 2.035629527e-01 wags = 1.241939206e-6
+ a1 = 0.0
+ a2 = 1.491657615e+00 wa2 = -3.400826546e-6
+ b0 = 0.0
+ b1 = 0.0
+ keta = 7.760368028e-02 wketa = -6.278681164e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.702831218e-01 wpclm = 1.699991175e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 1.213685421e-02 wpdiblc2 = -5.885785182e-8
+ pdiblcb = 7.204742588e-03 wpdiblcb = -5.049689656e-8
+ drout = 0.56
+ pscbe1 = 8.146533180e+08 wpscbe1 = -4.715832082e+2
+ pscbe2 = 9.259328818e-09 wpscbe2 = 1.699236528e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -8.208102985e-10 walpha0 = 6.369173011e-15
+ alpha1 = 3.451693611e-10 walpha1 = -1.695817347e-15
+ beta0 = 8.670873891e+00 wbeta0 = -2.682717678e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 4.268269277e+08 wbgidl = 5.032874685e+3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.662746100e-01 wkt1 = 1.700498298e-7
+ kt2 = -0.037961
+ at = 0.0
+ ute = -1.775648577e-01 wute = -8.514394977e-7
+ ua1 = 2.2116e-9
+ ub1 = -4.814392068e-19 wub1 = -2.159122689e-24
+ uc1 = 1.1985e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.11 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.218349223e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.416288885e-07 wvth0 = 5.989323423e-07 pvth0 = -1.512251211e-12
+ k1 = 6.137309884e-01 lk1 = -1.380171303e-06 wk1 = -1.177093566e-06 pk1 = 9.157306822e-12
+ k2 = -6.524407355e-02 lk2 = 6.975859659e-07 wk2 = 6.433634701e-07 pk2 = -4.379659986e-12
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.250103029e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -3.820600052e-07 wvoff = -1.708331533e-07 pvoff = 1.653294377e-12
+ nfactor = {5.680382139e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.620847515e-05 wnfactor = -1.992002797e-05 pnfactor = 1.168699594e-10
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.458006089e-02 lu0 = 7.073579886e-10 wu0 = -2.249111421e-08 pu0 = -3.148830999e-14
+ ua = 2.217428238e-10 lua = 2.495280376e-15 wua = -4.276131736e-16 pua = -2.165561029e-20
+ ub = 5.445028314e-19 lub = -3.115303717e-24 wub = -2.911920209e-24 pub = 2.188797131e-29
+ uc = -1.288046115e-10 luc = 4.494119866e-16 wuc = 3.027903196e-16 puc = -2.698394982e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.963722163e+05 lvsat = -7.961636780e-01 wvsat = -8.370125260e-01 pvsat = 1.306449056e-6
+ a0 = 1.702041139e-01 la0 = 6.651457839e-06 wa0 = 7.092841019e-06 pa0 = -2.904312526e-11
+ ags = -3.262537837e-01 lags = 4.269353330e-06 wags = 3.091539534e-06 pags = -1.490439388e-11
+ a1 = 0.0
+ a2 = 2.193373662e+00 la2 = -5.654547193e-06 wa2 = -6.851109611e-06 pa2 = 2.780296749e-11
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.219812607e-01 lketa = -1.163419087e-06 wketa = -1.330295355e-06 pketa = 5.660278098e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -9.850577616e-01 lpclm = 6.565592560e-06 wpclm = 3.424704472e-06 ppclm = -1.389803295e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 2.330904781e-02 lpdiblc2 = -9.002743530e-08 wpdiblc2 = -1.140331569e-07 ppdiblc2 = 4.446119881e-13
+ pdiblcb = 9.610145187e-03 lpdiblcb = -1.938314306e-08 wpdiblcb = -6.239572229e-08 ppdiblcb = 9.588276049e-14
+ drout = 0.56
+ pscbe1 = 6.399513998e+08 lpscbe1 = 1.407777756e+03 wpscbe1 = 3.612049508e+02 ppscbe1 = -6.710748559e-3
+ pscbe2 = 9.828202728e-09 lpscbe2 = -4.584082677e-15 wpscbe2 = 1.654898174e-15 ppscbe2 = 3.572859966e-22
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.755011481e-09 lalpha0 = 7.527951941e-15 walpha0 = 1.283096972e-14 palpha0 = -5.207025639e-20
+ alpha1 = 5.939040976e-10 lalpha1 = -2.004346792e-15 walpha1 = -3.416296119e-15 palpha1 = 1.386391042e-20
+ beta0 = 1.370051910e+01 lbeta0 = -4.052973615e-05 wbeta0 = -6.529427036e-05 pbeta0 = 3.099743795e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 9.280089982e-09 lagidl = -7.397472569e-14 wagidl = -6.381613022e-14 pagidl = 5.142412260e-19
+ bgidl = 2.406943004e+09 lbgidl = -1.595611196e+04 wbgidl = -7.579617032e+03 pbgidl = 1.016336024e-1
+ cgidl = 300.0
+ egidl = 6.232424737e-01 legidl = -4.216376804e-06 wegidl = -3.619227378e-06 pegidl = 2.916434948e-11
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.383374535e-01 lkt1 = -2.251223567e-07 wkt1 = 5.238929421e-08 pkt1 = 9.481285979e-13
+ kt2 = -4.602948251e-02 lkt2 = 6.501720374e-08 wkt2 = 7.254582875e-08 pkt2 = -5.845866208e-13
+ at = -4.644678458e+05 lat = 3.742760861e+00 wat = 1.370520960e+00 pat = -1.104389088e-5
+ ute = -2.284327672e+00 lute = 1.697665290e-05 wute = 1.370396236e-05 pute = -1.172899026e-10
+ ua1 = -4.872732784e-09 lua1 = 5.708675791e-14 wua1 = 4.755055594e-14 pua1 = -3.831704634e-19
+ ub1 = 4.280661081e-18 lub1 = -3.837381368e-23 wub1 = -3.387553793e-23 pub1 = 2.555762658e-28
+ uc1 = -8.772682101e-11 luc1 = 1.672689312e-15 wuc1 = 1.316003761e-15 puc1 = -1.060458203e-20
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.12 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.197008320e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.550238762e-07 wvth0 = 5.010757530e-07 pvth0 = -1.115132537e-12
+ k1 = 1.436482394e-01 lk1 = 5.275044066e-07 wk1 = 1.514702199e-06 pk1 = -1.766457998e-12
+ k2 = 1.482175958e-01 lk2 = -1.686777767e-07 wk2 = -5.621205905e-07 pk2 = 5.123992639e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.305467473e+00 ldsub = -3.025233734e-06 wdsub = -3.665405417e-06 pdsub = 1.487483830e-11
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-3.309449992e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.536580013e-07 wvoff = 7.465375197e-07 pvoff = -2.069551767e-12
+ nfactor = {-5.138644973e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.769697610e-05 wnfactor = 2.971692794e-05 pnfactor = -8.456524591e-11
+ eta0 = 3.629445019e-01 leta0 = -1.148236889e-06 weta0 = -1.391216046e-06 peta0 = 5.645791222e-12
+ etab = -3.173539985e-01 letab = 1.003804576e-06 wetab = 1.216220317e-06 petab = -4.935628804e-12
+ u0 = 1.920041310e-02 lu0 = -1.804281673e-08 wu0 = -4.342471394e-08 pu0 = 5.346379645e-14
+ ua = 1.248286660e-09 lua = -1.670609024e-15 wua = -5.468645293e-15 pua = -1.198244975e-21
+ ub = -6.704401318e-21 lub = -8.784110615e-25 wub = -1.297245174e-26 pub = 1.012354849e-29
+ uc = 7.072567646e-11 luc = -3.603158419e-16 wuc = -9.593953566e-16 puc = 2.423769064e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.935064971e+05 lvsat = -3.787171023e-01 wvsat = -6.713437615e-01 pvsat = 6.341370454e-7
+ a0 = 1.504119111e+00 la0 = 1.238204017e-06 wa0 = 1.802320290e-06 pa0 = -7.573292751e-12
+ ags = 9.053410156e-01 lags = -7.286677362e-07 wags = -2.399458612e-06 pags = 7.379010068e-12
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.718720861e-02 lketa = 9.123912012e-08 wketa = 2.364308178e-07 pketa = -6.977630530e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.711710877e-01 lpclm = 1.467602330e-06 wpclm = 2.670357827e-06 ppclm = -1.083676602e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 1.958338042e-03 lpdiblc2 = -3.382625427e-09 wpdiblc2 = -8.571857171e-09 ppdiblc2 = 1.663210538e-14
+ pdiblcb = 1.138689158e-02 lpdiblcb = -2.659348197e-08 wpdiblcb = -7.862398241e-08 ppdiblcb = 1.617397989e-13
+ drout = 0.56
+ pscbe1 = 1.177795099e+09 lpscbe1 = -7.748834100e+02 wpscbe1 = -2.613179234e+03 ppscbe1 = 5.359808106e-3
+ pscbe2 = 9.714411620e-09 lpscbe2 = -4.122299017e-15 wpscbe2 = -3.303811495e-15 ppscbe2 = 2.048057281e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.804308302e-03 lalpha0 = -1.138035941e-08 walpha0 = -1.939718109e-08 palpha0 = 7.871705840e-14
+ alpha1 = -1.529965338e-10 lalpha1 = 1.026702944e-15 walpha1 = 1.749957291e-15 palpha1 = -7.101624178e-21
+ beta0 = 6.830076436e+01 lbeta0 = -2.621068135e-04 wbeta0 = -4.497195919e-04 pbeta0 = 1.870037687e-9
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.827896470e-08 lagidl = 3.786460326e-14 wagidl = 1.277246235e-13 pagidl = -2.630637146e-19
+ bgidl = -3.277776617e+09 lbgidl = 7.113446663e+03 wbgidl = 2.958904719e+04 pbgidl = -4.920315572e-2
+ cgidl = 300.0
+ egidl = -9.464849474e-01 legidl = 2.153843924e-06 wegidl = 7.238454755e-06 pegidl = -1.489797042e-11
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.885254962e-01 lkt1 = 3.843662525e-07 wkt1 = 7.860510101e-07 pkt1 = -2.029195368e-12
+ kt2 = -2.961805949e-02 lkt2 = -1.583140850e-09 wkt2 = -5.037292669e-08 pkt2 = -8.576141508e-14
+ at = 7.396374157e+05 lat = -1.143702988e+00 wat = -2.078715862e+00 pat = 2.953698509e-6
+ ute = 4.275379492e+00 lute = -9.643753916e-06 wute = -3.257244387e-05 pute = 7.050762090e-11
+ ua1 = 1.778205058e-08 lua1 = -3.485020430e-14 wua1 = -1.021178964e-13 pua1 = 2.242095598e-19
+ ub1 = -1.142207047e-17 lub1 = 2.535054044e-23 wub1 = 6.995286598e-23 pub1 = -1.657770481e-28
+ uc1 = 1.053914531e-09 luc1 = -2.960285375e-15 wuc1 = -4.853423852e-15 puc1 = 1.443200403e-20
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.13 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.115038491e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.631603278e-08 wvth0 = 2.567798538e-07 pvth0 = -6.123300456e-13
+ k1 = 3.441237706e-01 lk1 = 1.148916827e-07 wk1 = 1.410361068e-06 pk1 = -1.551706214e-12
+ k2 = 9.070698347e-02 lk2 = -5.031115974e-08 wk2 = -5.554785069e-07 pk2 = 4.987287266e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -1.777998827e+00 ldsub = 3.321064100e-06 wdsub = 9.969402717e-06 pdsub = -1.318791475e-11
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-8.260781636e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.746213839e-08 wvoff = -3.338620956e-07 pvoff = 1.540943089e-13
+ nfactor = {5.718403781e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.648675933e-06 wnfactor = -2.487465546e-05 pnfactor = 2.779351330e-11
+ eta0 = -6.332327699e-01 leta0 = 9.020652863e-07 weta0 = 2.778498388e-06 peta0 = -2.936189936e-12
+ etab = -4.356761447e-01 letab = 1.247331668e-06 wetab = 3.013739089e-06 petab = -8.635228014e-12
+ u0 = 1.544821158e-02 lu0 = -1.032014812e-08 wu0 = -5.085994334e-08 pu0 = 6.876676253e-14
+ ua = 1.234268900e-09 lua = -1.641758092e-15 wua = -1.120198133e-14 pua = 1.060193525e-20
+ ub = -4.582033513e-19 lub = 5.085053234e-26 wub = 5.186701510e-24 pub = -5.782644695e-31
+ uc = -1.281517809e-10 luc = 4.900777452e-17 wuc = 3.183522009e-16 puc = -2.060526268e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.972796806e+04 lvsat = 4.069375282e-02 wvsat = -4.589710798e-01 pvsat = 1.970379633e-7
+ a0 = 7.652667837e-01 la0 = 2.758887710e-06 wa0 = 7.669779595e-06 pa0 = -1.964952147e-11
+ ags = -6.697612983e-01 lags = 2.513160593e-06 wags = 8.290140306e-06 pags = -1.462200174e-11
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.984863388e-02 lketa = -1.496405398e-07 wketa = -7.208480862e-07 pketa = 1.272479669e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.550356238e-01 lpclm = 6.009285795e-08 wpclm = -3.219465672e-06 ppclm = 1.285492006e-12
+ pdiblc1 = 5.400185245e-01 lpdiblc1 = -3.087636266e-07 wpdiblc1 = -7.050287543e-07 ppdiblc1 = 1.451069031e-12
+ pdiblc2 = 1.929540805e-04 lpdiblc2 = 2.508348806e-10 wpdiblc2 = -1.010233894e-09 ppdiblc2 = 1.068999200e-15
+ pdiblcb = -6.328925951e-02 lpdiblcb = 1.271027319e-07 wpdiblcb = 4.256558007e-07 ppdiblcb = -8.761537224e-13
+ drout = -1.281130262e-01 ldrout = 1.416253587e-06 wdrout = 2.641362983e-06 pdrout = -5.436374050e-12
+ pscbe1 = 8.026831294e+08 lpscbe1 = -2.839207079e+00 wpscbe1 = -1.855899705e+01 ppscbe1 = 1.963857391e-5
+ pscbe2 = 6.512077503e-09 lpscbe2 = 2.468648992e-15 wpscbe2 = 1.178359214e-14 ppscbe2 = -1.057186872e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.571816163e-03 lalpha0 = 5.859128675e-09 walpha0 = 3.853981849e-08 palpha0 = -4.052713603e-14
+ alpha1 = 3.458461000e-10 walpha1 = -1.700498298e-15
+ beta0 = -8.072685169e+01 lbeta0 = 4.461735508e-05 wbeta0 = 5.976938445e-04 pbeta0 = -2.857172257e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.375694777e-10 lagidl = -3.975489425e-17 wagidl = -1.847261916e-16 pagidl = 1.954717142e-22
+ bgidl = -1.144772259e+08 lbgidl = 6.028387549e+02 wbgidl = 6.782591659e+03 pbgidl = -2.263593130e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.528494218e-01 lkt1 = -1.006951735e-07 wkt1 = -2.439857979e-07 pkt1 = 9.079548943e-14
+ kt2 = -1.100563673e-02 lkt2 = -3.989067099e-08 wkt2 = -2.005427571e-07 pkt2 = 2.233136248e-13
+ at = 1.263896593e+05 lat = 1.184651468e-01 wat = -6.517949452e-01 pat = 1.685268663e-8
+ ute = 5.875887704e-01 lute = -2.053653686e-06 wute = 3.888542878e-06 pute = -4.535288194e-12
+ ua1 = 3.096559332e-09 lua1 = -4.624966773e-15 wua1 = 9.428069905e-15 pua1 = -5.371001639e-21
+ ub1 = -1.178299453e-19 lub1 = 2.084491709e-24 wub1 = -1.384060690e-23 pub1 = 6.684164009e-30
+ uc1 = -7.029051308e-10 luc1 = 6.555481491e-16 wuc1 = 3.834203493e-15 puc1 = -3.448609945e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.14 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-9.688930764e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -6.833066053e-08 wvth0 = -7.485605321e-07 pvth0 = 4.514909904e-13
+ k1 = 4.337756892e-01 lk1 = 2.002471196e-08 wk1 = -1.938973909e-07 pk1 = 1.458719600e-13
+ k2 = 6.790830539e-02 lk2 = -2.618628257e-08 wk2 = -1.491647458e-07 pk2 = 6.877969407e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.762938163e+00 ldsub = -4.258491944e-07 wdsub = -5.277183764e-06 pdsub = 2.945565661e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-4.726699562e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -9.485873468e-08 wvoff = -5.220837508e-07 pvoff = 3.532648178e-13
+ nfactor = {4.265986724e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.111771775e-06 wnfactor = -8.004954748e-06 pnfactor = 9.942502094e-12
+ eta0 = 5.598015732e-01 leta0 = -3.603678645e-07 weta0 = -7.643506933e-07 peta0 = 8.127466771e-13
+ etab = 1.576142245e+00 letab = -8.815141981e-07 wetab = -1.090896989e-05 petab = 6.097364950e-12
+ u0 = 1.868643654e-03 lu0 = 4.049343267e-09 wu0 = 5.458329076e-08 pu0 = -4.281010449e-14
+ ua = -1.879896993e-10 lua = -1.367667092e-16 wua = 6.059043419e-15 pua = -7.663163304e-21
+ ub = -1.369541069e-18 lub = 1.015200765e-24 wub = 2.290857686e-24 pub = 2.486030590e-30
+ uc = -1.451977056e-10 luc = 6.704526066e-17 wuc = 1.829306021e-16 puc = -6.275355356e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.406804453e+05 lvsat = -1.190396300e-01 wvsat = -1.494348214e+00 pvsat = 1.292642986e-6
+ a0 = 7.593313201e+00 la0 = -4.466346167e-06 wa0 = -3.227410280e-05 pa0 = 2.261789656e-11
+ ags = 3.019830496e+00 lags = -1.391054756e-06 wags = -1.484573699e-05 pags = 9.859689541e-12
+ a1 = 0.0
+ a2 = 1.137439019e-01 la2 = 7.261756153e-07 wa2 = 3.202529778e-06 pa2 = -3.388820935e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.058442930e-01 lketa = 9.976264457e-08 wketa = 1.047570979e-06 pketa = -5.988083339e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.401086399e-01 lpclm = 6.049731444e-07 wpclm = 6.593045595e-07 ppclm = -2.818906289e-12
+ pdiblc1 = 1.397527086e+00 lpdiblc1 = -1.216153461e-06 wpdiblc1 = -5.053617066e-06 ppdiblc1 = 6.052614725e-12
+ pdiblc2 = 2.319116742e-03 lpdiblc2 = -1.999006663e-09 wpdiblc2 = -1.574355450e-08 ppdiblc2 = 1.665935707e-14
+ pdiblcb = 1.481723724e-01 lpdiblcb = -9.665962308e-08 wpdiblcb = -8.514750475e-07 ppdiblcb = 4.752678272e-13
+ drout = 8.196335236e-01 ldrout = 4.133766205e-07 wdrout = -5.957456778e-07 pdrout = -2.010962779e-12
+ pscbe1 = 9.584265577e+08 lpscbe1 = -1.676422305e+02 wpscbe1 = -7.789710267e+02 ppscbe1 = 8.242837713e-4
+ pscbe2 = 8.952480327e-09 lpscbe2 = -1.137120634e-16 wpscbe2 = 8.086820754e-16 ppscbe2 = 1.041451860e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -7.360018060e-05 lalpha0 = 4.108146862e-11 walpha0 = 5.090874001e-10 palpha0 = -2.841573141e-16
+ alpha1 = 6.202939353e-10 lalpha1 = -2.904124659e-16 walpha1 = -3.598832567e-15 palpha1 = 2.008760374e-21
+ beta0 = -9.151594634e+01 lbeta0 = 5.603405137e-05 wbeta0 = 6.919674775e-04 pbeta0 = -3.854747561e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = -3.541088645e+08 lbgidl = 8.564097659e+02 wbgidl = 9.912763191e+03 pbgidl = -5.575846740e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.033063442e-01 lkt1 = -4.730317189e-08 wkt1 = -3.168241979e-07 pkt1 = 1.678708992e-13
+ kt2 = -7.089731804e-02 lkt2 = 2.348490942e-08 wkt2 = 5.188168858e-08 pkt2 = -4.379435087e-14
+ at = 4.889861352e+05 lat = -2.652235661e-01 wat = -1.547867957e+00 pat = 9.650502659e-7
+ ute = -2.740972355e+00 lute = 1.468529839e-06 wute = -8.410975546e-07 pute = 4.694754221e-13
+ ua1 = -5.717259703e-09 lua1 = 4.701552115e-15 wua1 = 1.028735372e-14 pua1 = -6.280269989e-21
+ ub1 = 6.683760870e-18 lub1 = -5.112747643e-24 wub1 = -1.894904682e-23 pub1 = 1.208976188e-29
+ uc1 = 7.827626433e-11 luc1 = -1.710745678e-16 wuc1 = 9.633200534e-16 puc1 = -4.107272158e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.15 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.143372894e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.905873933e-08 wvth0 = 2.611947650e-07 pvth0 = -1.121241237e-13
+ k1 = 1.674775243e-01 lk1 = 1.686643586e-07 wk1 = -1.256896303e-07 pk1 = 1.078004342e-13
+ k2 = 1.032089192e-01 lk2 = -4.589002615e-08 wk2 = 1.870734571e-07 pk2 = -1.188983836e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.506234072e+00 ldsub = -2.825646717e-07 wdsub = -8.031486762e-07 pdsub = 4.482934966e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-3.348552351e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 6.566439298e-08 wvoff = 7.906454829e-07 pvoff = -3.794612586e-13
+ nfactor = {-6.055308229e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.649265428e-06 wnfactor = 2.863832206e-05 pnfactor = -1.051067572e-11
+ eta0 = -7.956268817e-01 leta0 = 3.961916361e-07 weta0 = 1.544436202e-06 peta0 = -4.759489045e-13
+ etab = -6.265099033e-03 letab = 1.738109319e-09 wetab = 3.322089756e-08 petab = -1.023768400e-14
+ u0 = 1.354748408e-02 lu0 = -2.469435096e-09 wu0 = -4.213353876e-08 pu0 = 1.117432824e-14
+ ua = 1.381250568e-09 lua = -1.012669549e-15 wua = -1.780600139e-14 pua = 5.657588756e-21
+ ub = -1.404243242e-18 lub = 1.034570477e-24 wub = 1.779390502e-23 pub = -6.167305343e-30
+ uc = -9.715131829e-11 luc = 4.022720865e-17 wuc = 4.418849812e-16 puc = -2.072941194e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.066172986e+04 lvsat = 2.683373191e-02 wvsat = 1.704445450e+00 pvsat = -4.928276737e-7
+ a0 = -1.990211184e+00 la0 = 8.828896391e-07 wa0 = 1.920493706e-05 pa0 = -6.116159118e-12
+ ags = -2.704776614e+00 lags = 1.804249195e-06 wags = 1.348703437e-05 pags = -5.954813450e-12
+ a1 = 0.0
+ a2 = 2.172512196e+00 la2 = -4.229670835e-07 wa2 = -6.405059556e-06 pa2 = 1.973847203e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = 8.288594409e-03 lketa = -1.975990917e-08 wketa = 2.136651277e-07 pketa = -1.333471046e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.256475266e+00 lpclm = -4.088682150e-07 wpclm = -8.034023183e-06 ppclm = 2.033448457e-12
+ pdiblc1 = -2.368648635e+00 lpdiblc1 = 8.860128408e-07 wpdiblc1 = 1.404955946e-05 ppdiblc1 = -4.610205317e-12
+ pdiblc2 = -1.307842849e-02 lpdiblc2 = 6.595441158e-09 wpdiblc2 = 3.023236036e-08 ppdiblc2 = -9.003019333e-15
+ pdiblcb = -0.025
+ drout = 2.433146159e+00 ldrout = -4.872377272e-07 wdrout = -6.901943446e-06 pdrout = 1.508967630e-12
+ pscbe1 = 4.831468847e+08 lpscbe1 = 9.764462454e+01 wpscbe1 = 1.557942053e+03 ppscbe1 = -4.801110026e-4
+ pscbe2 = 1.830049552e-08 lpscbe2 = -5.331493705e-15 wpscbe2 = 5.971335735e-15 ppscbe2 = -1.840186534e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.675033813e-08 lalpha0 = 3.731385323e-14 walpha0 = 3.286978983e-13 palpha0 = -1.834693059e-19
+ alpha1 = 5.263175705e-10 lalpha1 = -2.379576784e-16 walpha1 = -2.096170242e-15 palpha1 = 1.170019344e-21
+ beta0 = -2.444356147e+01 lbeta0 = 1.859625830e-05 wbeta0 = 1.671889047e-04 pbeta0 = -9.255910005e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 9.705604771e+08 lbgidl = 1.170190795e+02 wbgidl = 7.494007101e+02 pbgidl = -4.611327038e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.181394052e-01 lkt1 = -3.902380224e-08 wkt1 = -4.441528544e-07 pkt1 = 2.389419354e-13
+ kt2 = -2.253777679e-02 lkt2 = -3.507935717e-09 wkt2 = -2.139369495e-08 pkt2 = -2.894230050e-15
+ at = -4.913403019e+04 lat = 3.513896664e-02 wat = 5.714547578e-01 pat = -2.178920940e-7
+ ute = -1.142593988e-01 lute = 2.377468614e-09 wute = -4.821191556e-07 pute = 2.691044491e-13
+ ua1 = 4.640423158e-09 lua1 = -1.079795728e-15 wua1 = -2.719857171e-15 pua1 = 9.799649116e-22
+ ub1 = -5.055876524e-18 lub1 = 1.439965761e-24 wub1 = 9.118556950e-24 pub1 = -3.576732520e-30
+ uc1 = -3.525897731e-10 luc1 = 6.942192829e-17 wuc1 = 5.445839179e-17 puc1 = 9.657209791e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.16 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.077690806e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.817490334e-09 wvth0 = -1.747409305e-07 pvth0 = 2.221817957e-14
+ k1 = -9.500866665e-01 lk1 = 5.130641153e-07 wk1 = 6.164307903e-06 pk1 = -1.830588106e-12
+ k2 = 6.438783750e-01 lk2 = -2.125081323e-07 wk2 = -2.607043427e-06 pk2 = 7.421646164e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 4.310802976e+00 ldsub = -1.146848671e-06 wdsub = -2.230026273e-05 pdsub = 7.073059134e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {1.361095612e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.947282830e-08 wvoff = -1.386531848e-06 pvoff = 2.914794794e-13
+ nfactor = {5.094977826e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.869182251e-07 wnfactor = -2.003488323e-05 pnfactor = 4.488945953e-12
+ eta0 = 0.49
+ etab = -6.249996470e-04 letab = -1.087886309e-16 wetab = -1.735747192e-15 petab = 5.349052139e-22
+ u0 = 2.580052328e-02 lu0 = -6.245454184e-09 wu0 = -1.210097171e-07 pu0 = 3.548160011e-14
+ ua = 3.927119329e-09 lua = -1.797229925e-15 wua = -2.897646703e-14 pua = 9.099991152e-21
+ ub = -1.850042596e-18 lub = 1.171952464e-24 wub = 1.447810786e-23 pub = -5.145476131e-30
+ uc = 7.550696401e-11 luc = -1.298089421e-17 wuc = -2.641952981e-16 puc = 1.029864029e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.785003596e+05 lvsat = -3.454204920e-02 wvsat = -1.235703209e+00 pvsat = 4.132379385e-7
+ a0 = 4.250541984e+00 la0 = -1.040323265e-06 wa0 = -1.982640326e-05 pa0 = 5.912129029e-12
+ ags = 9.614366936e+00 lags = -1.992141273e-06 wags = -2.569305810e-05 pags = 6.119315649e-12
+ a1 = 0.0
+ a2 = -2.386238860e-01 la2 = 3.200727230e-07 wa2 = 8.958846823e-06 pa2 = -2.760847826e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = 4.524069517e-01 lketa = -1.566238633e-07 wketa = -3.717613238e-06 pketa = 1.078154949e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.278602960e+00 lpclm = -1.075173065e-07 wpclm = -3.402469773e-06 ppclm = 6.061426423e-13
+ pdiblc1 = 9.884037730e-01 lpdiblc1 = -1.485299997e-07 wpdiblc1 = -5.015338425e-06 ppdiblc1 = 1.265024264e-12
+ pdiblc2 = 4.534238807e-03 lpdiblc2 = 1.167745478e-09 wpdiblc2 = 1.155654995e-08 ppdiblc2 = -3.247694837e-15
+ pdiblcb = 1.077981675e+00 lpdiblcb = -3.399058629e-07 wpdiblcb = -4.089903515e-06 ppdiblcb = 1.260385566e-12
+ drout = 3.803635885e-01 ldrout = 1.453682775e-07 wdrout = 7.176876934e-07 pdrout = -8.391740988e-13
+ pscbe1 = 7.982595082e+08 lpscbe1 = 5.363673512e-01 wpscbe1 = 1.444546677e+01 ppscbe1 = -4.451659493e-6
+ pscbe2 = -7.632256620e-08 lpscbe2 = 2.382849523e-14 wpscbe2 = 3.399181085e-13 ppscbe2 = -1.047525635e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 6.926438053e-08 lalpha0 = -4.601802615e-15 walpha0 = -3.400758642e-13 palpha0 = 2.262670452e-20
+ alpha1 = -2.458461000e-10 walpha1 = 1.700498298e-15
+ beta0 = 4.392732246e+01 lbeta0 = -2.473596996e-06 wbeta0 = -1.777579658e-04 pbeta0 = 1.374317702e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = -1.672767534e+09 lbgidl = 9.316134726e+02 wbgidl = 1.651627500e+04 pbgidl = -5.320010353e-3
+ cgidl = 3.253088227e+03 lcgidl = -9.100531990e-04 wcgidl = -1.452010447e-02 pcgidl = 4.474660596e-9
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.859663678e-01 lkt1 = -4.893856716e-08 wkt1 = -2.776421945e-07 pkt1 = 1.876283453e-13
+ kt2 = 3.128700326e-02 lkt2 = -2.009511819e-08 wkt2 = -1.355303575e-07 pkt2 = 3.227926524e-14
+ at = 1.314770788e+05 lat = -2.051995882e-02 wat = -3.076642469e-01 pat = 5.302600972e-8
+ ute = -1.881907172e+00 lute = 5.471134829e-07 wute = 1.542326393e-05 pute = -4.632457455e-12
+ ua1 = 3.718687187e-09 lua1 = -7.957443536e-16 wua1 = 2.025521818e-15 pua1 = -4.824185314e-22
+ ub1 = -1.926822064e-18 lub1 = 4.756850477e-25 wub1 = -1.095238321e-23 pub1 = 2.608529108e-30
+ uc1 = -5.286739547e-10 luc1 = 1.236857906e-16 wuc1 = 1.619350579e-15 puc1 = -3.856807273e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.17 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -3.7585e-8
+ vth0 = {-6.578848420e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -9.767502642e-08 wvth0 = -2.182049861e-06 pvth0 = 5.360090794e-13
+ k1 = 2.390136955e+00 lk1 = -3.026394673e-07 wk1 = -1.482150288e-05 pk1 = 3.393698268e-12
+ k2 = -2.124915784e-01 lk2 = -9.156529137e-09 wk2 = 3.254737873e-06 pk2 = -7.006121981e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -6.836326058e+00 ldsub = 1.615704953e-06 wdsub = 6.447181430e-05 pdsub = -1.456371387e-11
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {2.376177567e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.110472533e-07 wvoff = -2.631182126e-06 pvoff = 6.298819929e-13
+ nfactor = {-8.245015718e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.560879603e-06 wnfactor = 4.916383291e-05 pnfactor = -1.284808031e-11
+ eta0 = 2.515182791e+00 leta0 = -5.167658928e-07 weta0 = 9.318538912e-09 peta0 = -2.377811574e-15
+ etab = 4.371577051e-01 letab = -1.117090129e-07 wetab = -1.199149302e-06 petab = 3.059869276e-13
+ u0 = -5.592273068e-02 lu0 = 1.416208308e-08 wu0 = 3.499759249e-07 pu0 = -8.216721513e-14
+ ua = -2.015289989e-08 lua = 4.218986642e-15 wua = 1.041569821e-13 pua = -2.422213566e-20
+ ub = 1.556585862e-17 lub = -3.188411909e-24 wub = -7.632171593e-23 pub = 1.765664323e-29
+ uc = 3.786695771e-10 luc = -9.126544310e-17 wuc = -2.483641464e-15 puc = 5.773698106e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.222364404e+05 lvsat = 3.973143193e-02 wvsat = 3.880496570e+00 pvsat = -8.627668321e-7
+ a0 = -9.471245292e-01 la0 = 2.117095346e-07 wa0 = 1.135545682e-05 pa0 = -1.622552700e-12
+ ags = 1.25
+ a1 = 0.0
+ a2 = 3.640749875e+00 la2 = -6.469810608e-07 wa2 = -2.324683479e-05 pa2 = 5.260013294e-12
+ b0 = -5.470141024e-23 lb0 = 1.395815885e-29 wb0 = 2.689625674e-28 pb0 = -6.863117833e-35
+ b1 = 0.0
+ keta = -1.332667628e+00 lketa = 2.876941836e-07 wketa = 5.154315145e-06 pketa = -1.108738917e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.301832019e+00 lpclm = -3.762889915e-07 wpclm = -7.145943031e-06 ppclm = 1.604629713e-12
+ pdiblc1 = 1.258907372e+00 lpdiblc1 = -2.281561160e-07 wpdiblc1 = 5.999498438e-06 ppdiblc1 = -1.455337278e-12
+ pdiblc2 = 4.246648917e-02 lpdiblc2 = -8.428075992e-09 wpdiblc2 = 4.358617857e-08 ppdiblc2 = -1.165250780e-14
+ pdiblcb = -3.260303694e+00 lpdiblcb = 7.428327545e-07 wpdiblcb = 2.099336854e-05 ppdiblcb = -5.050149683e-12
+ drout = 9.210563789e-01 ldrout = 1.777573517e-08 wdrout = -2.386466509e-05 pdrout = 5.373606638e-12
+ pscbe1 = 8.043510224e+08 lpscbe1 = -9.797197118e-01 wpscbe1 = -3.611194844e+01 ppscbe1 = 8.131327431e-6
+ pscbe2 = 1.281686588e-07 lpscbe2 = -2.665071015e-14 wpscbe2 = -8.344076430e-13 ppscbe2 = 1.874231533e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.803937995e-07 lalpha0 = -5.880416203e-14 walpha0 = -1.378182749e-12 palpha0 = 2.891354780e-19
+ alpha1 = -2.458461000e-10 walpha1 = 1.700498298e-15
+ beta0 = 7.529090556e+01 lbeta0 = -1.065320188e-05 wbeta0 = -2.874869962e-04 pbeta0 = 4.272368852e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 5.584260650e+09 lbgidl = -8.536660869e+02 wbgidl = -2.309211324e+04 pbgidl = 4.407132569e-3
+ cgidl = -7.082369261e+03 lcgidl = 1.662288087e-03 wcgidl = 3.629853383e-02 pcgidl = -8.173340863e-9
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -2.8385e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -9.133765654e-01 lkt1 = 8.214757609e-08 wkt1 = 3.300222912e-06 pkt1 = -7.119430353e-13
+ kt2 = -1.055525597e+00 lkt2 = 2.557925121e-07 wkt2 = 6.284429790e-06 pkt2 = -1.603597949e-12
+ at = 5.631030081e+05 lat = -1.321226123e-01 wat = -3.238854480e+00 pat = 8.047626900e-7
+ ute = 6.892186448e+00 lute = -1.652720346e-06 wute = -4.295779153e-05 pute = 9.933982829e-12
+ ua1 = -4.036209537e-09 lua1 = 1.126274331e-15 wua1 = 2.869844507e-14 pua1 = -7.322982228e-21
+ ub1 = 6.586948311e-18 lub1 = -1.662820488e-24 wub1 = -3.925617990e-23 pub1 = 1.001699943e-29
+ uc1 = 6.855978692e-10 luc1 = -1.773315574e-16 wuc1 = -3.392632281e-15 puc1 = 8.656979791e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.18 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.119541292e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.047063488e-07 wvth0 = -1.484194283e-08 pvth0 = 1.485057639e-12
+ k1 = 4.560777990e-01 lk1 = -1.951732559e-06 wk1 = -9.295924833e-08 pk1 = 9.301332273e-12
+ k2 = 2.635887808e-02 lk2 = 9.408059408e-07 wk2 = 3.899242705e-08 pk2 = -3.901510895e-12
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.686964901e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.238329983e-07 wvoff = 3.595926197e-09 pvoff = -3.598017948e-13
+ nfactor = {1.738809537e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -9.400658863e-06 wnfactor = -6.925838434e-08 pnfactor = 6.929867194e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.092315493e-02 lu0 = -7.189872763e-09 wu0 = 1.560507476e-09 pu0 = -1.561415223e-13
+ ua = 5.981384025e-11 lua = 2.125154458e-15 wua = 3.302604766e-16 pua = -3.304525892e-20
+ ub = 1.775228247e-19 lub = -4.793896459e-24 wub = -2.213893682e-25 pub = 2.215181504e-29
+ uc = -8.803843507e-11 luc = 1.037376998e-15 wuc = 5.330263683e-17 puc = -5.333364298e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.099507328e+05 lvsat = -9.956521115e-1
+ a0 = 1.421551000e+00 la0 = 7.849463398e-06 wa0 = 1.328113581e-07 pa0 = -1.328886144e-11
+ ags = 3.638561992e-01 lags = 1.926880291e-06 wags = 4.651585385e-09 pags = -4.654291212e-13
+ a1 = 0.0
+ a2 = 1.050132918e+00 la2 = -5.017208586e-6
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.983487367e-03 lketa = -1.616196532e-06 wketa = -3.390253624e-08 pketa = 3.392225735e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 8.257014001e-03 lpclm = 6.727175723e-06 wpclm = 2.073338791e-07 ppclm = -2.074544852e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 4.539520438e-03 lpdiblc2 = -9.124515026e-08 wpdiblc2 = -2.168426241e-10 ppdiblc2 = 2.169687615e-14
+ pdiblcb = 1.210095417e-03 lpdiblcb = -1.306599062e-07 wpdiblcb = -2.759850702e-09 ppdiblcb = 2.761456107e-13
+ drout = 0.56
+ pscbe1 = 7.795801692e+08 lpscbe1 = -3.312429644e+03 wpscbe1 = -1.285866536e+02 ppscbe1 = 1.286614525e-2
+ pscbe2 = 9.390573532e-09 lpscbe2 = 1.144855257e-14 wpscbe2 = 4.394000444e-16 ppscbe2 = -4.396556434e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.308721188e-10 lalpha0 = 2.310064171e-14 walpha0 = 6.734359625e-16 palpha0 = -6.738277002e-20
+ alpha1 = 1.614706090e-10 lalpha1 = -6.150636650e-15 walpha1 = -1.793049719e-16 palpha1 = 1.794092736e-20
+ beta0 = 5.109397242e+00 lbeta0 = -3.171925459e-05 wbeta0 = 3.861783732e-07 pbeta0 = -3.864030132e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.167961556e-10 lagidl = -1.680592595e-15 wagidl = -8.258538710e-17 pagidl = 8.263342702e-21
+ bgidl = 9.155344705e+08 lbgidl = 2.390491035e+04 wbgidl = 8.098354974e+02 pbgidl = -8.103065787e-2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.529186375e-01 lkt1 = 1.123516919e-06 wkt1 = 4.288227755e-08 pkt1 = -4.290722217e-12
+ kt2 = -0.037961
+ at = 0.0
+ ute = -2.804122754e-01 lute = -2.025950268e-06 wute = -3.782990019e-08 pute = 3.785190585e-12
+ ua1 = 2.316731773e-09 lua1 = -1.051929285e-14 wua1 = -5.169247294e-16 pua1 = 5.172254245e-20
+ ub1 = -1.039756497e-18 lub1 = 2.463096916e-23 wub1 = 1.366910804e-24 pub1 = -1.367705936e-28
+ uc1 = 2.317577447e-10 luc1 = -1.119728414e-14 wuc1 = -5.502416519e-16 puc1 = 5.505617275e-20
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.19 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.104350158e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} wvth0 = 5.919560091e-8
+ k1 = 3.587741786e-01 wk1 = 3.707586418e-7
+ k2 = 7.326275519e-02 wk2 = -1.555173859e-7
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.625227963e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} wvoff = -1.434199111e-8
+ nfactor = {1.270139720e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 2.762301221e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.056470385e-02 wu0 = -6.223927611e-9
+ ua = 1.657634088e-10 wua = -1.317210799e-15
+ ub = -6.147686764e-20 wub = 8.829892982e-25
+ uc = -3.632000821e-11 wuc = -2.125922228e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 160312.5
+ a0 = 1.812885972e+00 wa0 = -5.297047859e-7
+ ags = 4.599208099e-01 wags = -1.855238194e-8
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -7.759198545e-02 wketa = 1.352168667e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 3.436403378e-01 wpclm = -8.269303894e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -9.506230630e-06 wpdiblc2 = 8.648550654e-10
+ pdiblcb = -5.303953784e-03 wpdiblcb = 1.100738782e-8
+ drout = 0.56
+ pscbe1 = 6.144390001e+08 wpscbe1 = 5.128549758e+2
+ pscbe2 = 9.961341083e-09 wpscbe2 = -1.752503022e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.020810298e-09 walpha0 = -2.685931817e-15
+ alpha1 = -1.451693611e-10 walpha1 = 7.151399031e-16
+ beta0 = 3.528033908e+00 wbeta0 = -1.540233723e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 3.301021729e-11 wagidl = 3.293835364e-16
+ bgidl = 2.107313698e+09 wbgidl = -3.229947687e+3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.969057052e-01 wkt1 = -1.710316646e-7
+ kt2 = -0.037961
+ at = 0.0
+ ute = -3.814160194e-01 wute = 1.508807641e-7
+ ua1 = 1.792292463e-09 wua1 = 2.061702456e-15
+ ub1 = 1.882203906e-19 wub1 = -5.451786696e-24
+ uc1 = -3.264828198e-10 wuc1 = 2.194583661e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.20 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.092313567e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -9.699289264e-08 wvth0 = -2.077514606e-08 pvth0 = 6.444178742e-13
+ k1 = 2.614799177e-01 lk1 = 7.840136943e-07 wk1 = 5.548974727e-07 pk1 = -1.483822003e-12
+ k2 = 1.190354553e-01 lk2 = -3.688441992e-07 wk2 = -2.627245997e-07 pk2 = 8.638939540e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.209489699e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -3.350089607e-07 wvoff = -1.908024109e-07 pvoff = 1.421948061e-12
+ nfactor = {3.126484355e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.495874065e-05 wnfactor = -7.362711767e-06 pnfactor = 6.155589236e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 8.967616489e-03 lu0 = 1.286960142e-08 wu0 = 5.104837144e-09 pu0 = -9.128911229e-14
+ ua = -2.042102782e-10 lua = 2.981310866e-15 wua = 1.666765004e-15 pua = -2.404538430e-20
+ ub = 1.392375116e-19 lub = -1.617390589e-24 wub = -9.192622423e-25 pub = 1.452284930e-29
+ uc = 4.315731916e-11 luc = -6.404418151e-16 wuc = -5.427330802e-16 puc = 2.660331153e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.317190305e+05 lvsat = -5.754059615e-01 wvsat = -2.742565407e-02 pvsat = 2.210005828e-7
+ a0 = 1.539751735e+00 la0 = 2.200962112e-06 wa0 = 3.588821891e-07 pa0 = -7.160384904e-12
+ ags = 7.318554019e-02 lags = 3.116378548e-06 wags = 1.127527535e-06 pags = -9.235306807e-12
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -6.465987841e-02 lketa = -1.042091170e-07 wketa = 7.909676807e-08 pketa = 4.522252953e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.026288934e-02 lpclm = 2.364085353e-06 wpclm = -1.665886414e-06 ppclm = 6.760450268e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -2.372773431e-04 lpdiblc2 = 1.835418346e-09 wpdiblc2 = 1.742287286e-09 ppdiblc2 = -7.070497994e-15
+ pdiblcb = -6.948780339e-03 lpdiblcb = 1.325429200e-08 wpdiblcb = 1.902322293e-08 ppdiblcb = -6.459296200e-14
+ drout = 0.56
+ pscbe1 = 6.157478114e+08 lpscbe1 = -1.054662383e+01 wpscbe1 = 4.802121070e+02 ppscbe1 = 2.630417861e-4
+ pscbe2 = 1.164565576e-08 lpscbe2 = -1.357249397e-14 wpscbe2 = -7.281376603e-15 ppscbe2 = 4.455260322e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.955011481e-09 lalpha0 = -7.527951941e-15 walpha0 = -5.410923798e-15 palpha0 = 2.195844863e-20
+ alpha1 = -3.939040976e-10 lalpha1 = 2.004346792e-15 walpha1 = 1.440679728e-15 palpha1 = -5.846523253e-21
+ beta0 = 2.122958736e+00 lbeta0 = 1.132233460e-05 wbeta0 = -8.368309095e-06 pbeta0 = 5.502179212e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -9.374125676e-09 lagidl = 7.580430024e-14 wagidl = 2.790519314e-14 pagidl = -2.222105617e-19
+ bgidl = 9.625160994e+08 lbgidl = 9.224973666e+03 wbgidl = -4.774826088e+02 pbgidl = -2.217983152e-2
+ cgidl = 300.0
+ egidl = -4.232424737e-01 legidl = 4.216376804e-06 wegidl = 1.526257483e-06 pegidl = -1.229884226e-11
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.060415940e-01 lkt1 = -7.321984546e-07 wkt1 = -5.980991277e-07 pkt1 = 3.441382219e-12
+ kt2 = -3.127516492e-02 lkt2 = -5.387559563e-8
+ at = -1.911478901e+05 lat = 1.540302194e+00 wat = 2.662805647e-02 pat = -2.145734058e-7
+ ute = 9.877237843e-01 lute = -1.103276129e-05 wute = -2.384459432e-06 pute = 2.043020231e-11
+ ua1 = 3.953351649e-09 lua1 = -1.741418231e-14 wua1 = 4.153387220e-15 pua1 = -1.685515141e-20
+ ub1 = -1.881906574e-19 lub1 = 3.033184215e-24 wub1 = -1.190254251e-23 pub1 = 5.198128696e-29
+ uc1 = -7.192353733e-10 luc1 = 3.164866844e-15 wuc1 = 4.421082055e-15 puc1 = -1.794150256e-20
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.21 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.176653586e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.452732404e-07 wvth0 = 4.009931128e-07 pvth0 = -1.067189421e-12
+ k1 = 2.347271415e-01 lk1 = 8.925810081e-07 wk1 = 1.066874341e-06 pk1 = -3.561511172e-12
+ k2 = 9.215186372e-02 lk2 = -2.597460141e-07 wk2 = -2.864497591e-07 pk2 = 9.601746841e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.641395646e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.460828147e-07 wvoff = 4.180604082e-07 pvoff = -1.048920766e-12
+ nfactor = {-2.144943869e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.433611228e-06 wnfactor = 1.499713312e-05 pnfactor = -2.918415937e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.952108394e-02 lu0 = -2.995816359e-08 wu0 = -4.500142747e-08 pu0 = 1.120506276e-13
+ ua = 2.491382712e-09 lua = -7.957863738e-15 wua = -1.158085162e-14 pua = 2.971569605e-20
+ ub = -1.522062949e-18 lub = 5.124449102e-24 wub = 7.437927331e-24 pub = -1.939204671e-29
+ uc = -2.086368653e-10 luc = 3.813817906e-16 wuc = 4.142084711e-16 puc = -1.223100343e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.725486565e+05 lvsat = -3.352825250e-01 wvsat = -7.660349378e-02 pvsat = 4.205726166e-7
+ a0 = 1.633986383e+00 la0 = 1.818541891e-06 wa0 = 1.163773041e-06 pa0 = -1.042676881e-11
+ ags = 2.059386023e-01 lags = 2.577644054e-06 wags = 1.039448501e-06 pags = -8.877867111e-12
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.524594813e-02 lketa = -2.235758465e-07 wketa = -1.896030858e-08 pketa = 8.501575821e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.249047297e-01 lpclm = 3.209107602e-08 wpclm = 9.310771008e-07 ppclm = -3.778469158e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000215
+ pdiblcb = -4.109301952e-02 lpdiblcb = 1.518174191e-07 wpdiblcb = 1.794156471e-07 ppdiblcb = -7.154926858e-13
+ drout = 0.56
+ pscbe1 = 4.222049007e+08 lpscbe1 = 7.748834100e+02 wpscbe1 = 1.101998837e+03 ppscbe1 = -2.260274466e-3
+ pscbe2 = -2.516689863e-09 lpscbe2 = 4.390071215e-14 wpscbe2 = 5.683556047e-14 ppscbe2 = -2.156448273e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -2.804308102e-03 lalpha0 = 1.138035941e-08 walpha0 = 8.179948288e-09 palpha0 = -3.319562074e-14
+ alpha1 = 3.529965338e-10 lalpha1 = -1.026702944e-15 walpha1 = -7.379711554e-16 palpha1 = 2.994812404e-21
+ beta0 = -6.500551177e+01 lbeta0 = 2.837410798e-04 wbeta0 = 2.057369700e-04 pbeta0 = -8.138538282e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.877834382e-08 lagidl = -3.844320691e-14 wagidl = -5.448327202e-14 pagidl = 1.121358360e-19
+ bgidl = 5.072005898e+09 lbgidl = -7.452034549e+03 wbgidl = -1.146618215e+04 pbgidl = 2.241417929e-2
+ cgidl = 300.0
+ egidl = 1.146484947e+00 legidl = -2.153843924e-06 wegidl = -3.052514966e-06 pegidl = 6.282594727e-12
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.557957466e-01 lkt1 = 2.813463550e-07 wkt1 = 6.251213845e-07 pkt1 = -1.522654567e-12
+ kt2 = -3.963212913e-02 lkt2 = -1.996161419e-08 wkt2 = -1.134527335e-09 pkt2 = 4.604104797e-15
+ at = 3.736849569e+05 lat = -7.518855210e-01 wat = -2.793561657e-01 pat = 1.027162585e-6
+ ute = -3.341369131e+00 lute = 6.535433703e-06 wute = 4.878515000e-06 pute = -9.044182641e-12
+ ua1 = -2.417438447e-09 lua1 = 8.439566937e-15 wua1 = -2.798584398e-15 pua1 = 1.135713124e-20
+ ub1 = 2.155285152e-18 lub1 = -6.477039009e-24 wub1 = 3.194067404e-24 pub1 = -9.283322484e-30
+ uc1 = 2.827554383e-11 luc1 = 1.313404651e-16 wuc1 = 1.895630492e-16 puc1 = -7.692790794e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.22 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.002943848e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.122509318e-07 wvth0 = -2.943807638e-07 pvth0 = 3.640082307e-13
+ k1 = 9.215888962e-01 lk1 = -5.210972496e-07 wk1 = -1.428989912e-06 pk1 = 1.575401759e-12
+ k2 = -9.950755690e-02 lk2 = 1.347216556e-07 wk2 = 3.797915514e-07 pk2 = -4.110631938e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 5.953642950e-02 ldsub = 1.030039107e-06 wdsub = 9.343851877e-07 pdsub = -1.923123562e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.028685574e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -8.584033410e-08 wvoff = -2.342416122e-07 pvoff = 2.936276837e-13
+ nfactor = {3.627615214e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.272327224e-06 wnfactor = 1.458619788e-06 pnfactor = -1.319597384e-12
+ eta0 = -6.969401366e-02 leta0 = 3.080957281e-07 weta0 = 7.622279644e-09 peta0 = -1.568794730e-14
+ etab = -6.393318239e-01 letab = 1.171781680e-06 wetab = 4.015098178e-06 petab = -8.263754618e-12
+ u0 = -2.027177630e-04 lu0 = 1.063677336e-08 wu0 = 2.609445545e-08 pu0 = -3.427678577e-14
+ ua = -2.515243708e-09 lua = 2.346624561e-15 wua = 7.234079707e-15 pua = -9.008631156e-21
+ ub = 1.624146126e-18 lub = -1.350984031e-24 wub = -5.052048447e-24 pub = 6.314446734e-30
+ uc = 2.495928184e-11 luc = -9.939879166e-17 wuc = -4.344829519e-16 puc = 5.236508833e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -6.645388311e+04 lvsat = 1.566253319e-01 wvsat = 3.089629002e-01 pvsat = -3.729885685e-7
+ a0 = 4.026097252e+00 la0 = -3.104828936e-06 wa0 = -8.363469472e-06 pa0 = 9.181915910e-12
+ ags = 2.384380940e+00 lags = -1.905960613e-06 wags = -6.726838859e-06 pags = 7.106472544e-12
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.838344618e-01 lketa = 2.880615748e-07 wketa = 8.215072282e-07 pketa = -8.796674881e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 7.078303251e-01 lpclm = -1.385838967e-07 wpclm = -2.003976500e-06 ppclm = 2.262370112e-12
+ pdiblc1 = 3.769525731e-01 lpdiblc1 = 2.685382261e-08 wpdiblc1 = 9.675380975e-08 ppdiblc1 = -1.991357886e-13
+ pdiblc2 = -1.250655000e-05 lpdiblc2 = 4.682471560e-10
+ pdiblcb = 9.369524914e-02 lpdiblcb = -1.255997518e-07 wpdiblcb = -3.462247835e-07 ppdiblcb = 3.663646792e-13
+ drout = 8.531929070e-01 ldrout = -6.034408453e-07 wdrout = -2.183641748e-06 pdrout = 4.494305937e-12
+ pscbe1 = 7.973168706e+08 lpscbe1 = 2.839207079e+00 wpscbe1 = 7.826479292e+00 ppscbe1 = -8.281745592e-6
+ pscbe2 = 2.909603293e-08 lpscbe2 = -2.116364552e-14 wpscbe2 = -9.925995514e-14 ppscbe2 = 1.056262801e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 5.571816363e-03 lalpha0 = -5.859128675e-09 walpha0 = -1.625255344e-08 palpha0 = 1.709062133e-14
+ alpha1 = -1.458461000e-10 walpha1 = 7.171138977e-16
+ beta0 = 9.057912482e+01 lbeta0 = -3.647855174e-05 wbeta0 = -2.446042802e-04 pbeta0 = 1.130250226e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.257387809e+09 lbgidl = 3.990979631e+02 wbgidl = 3.723828851e+01 pbgidl = -1.261815548e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.426574637e-01 lkt1 = -1.573284647e-07 wkt1 = -2.940988605e-07 pkt1 = 3.692569649e-13
+ kt2 = -3.805808425e-02 lkt2 = -2.320126614e-08 wkt2 = -6.752798277e-08 pkt2 = 1.412531230e-13
+ at = -1.079554326e+05 lat = 2.394122795e-01 wat = 5.004615926e-01 pat = -5.778349305e-7
+ ute = 3.388835515e+00 lute = -7.316471593e-06 wute = -9.884968868e-06 pute = 2.134157695e-11
+ ua1 = 8.186260091e-09 lua1 = -1.338464728e-14 wua1 = -1.559759173e-14 pua1 = 3.769966416e-20
+ ub1 = -4.974231773e-18 lub1 = 8.196718841e-24 wub1 = 1.003794209e-23 pub1 = -2.336918004e-29
+ uc1 = -4.655148979e-11 luc1 = 2.853472209e-16 wuc1 = 6.069638362e-16 puc1 = -1.628360857e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.23 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.104122894e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -5.186300669e-09 wvth0 = -8.364606856e-08 pvth0 = 1.410150983e-13
+ k1 = 5.081631949e-01 lk1 = -8.362257518e-08 wk1 = -5.596549539e-07 pk1 = 6.554975863e-13
+ k2 = -1.248490584e-02 lk2 = 4.263689692e-08 wk2 = 2.461224032e-07 pk2 = -2.696185112e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.069737541e+00 ldsub = -3.892540326e-08 wdsub = -1.868770375e-06 pdsub = 1.043091560e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.221553679e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.543160987e-08 wvoff = -1.538634658e-07 pvoff = 2.085739404e-13
+ nfactor = {3.511880018e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.059975496e-06 wnfactor = -4.297070899e-06 pnfactor = 4.770901830e-12
+ eta0 = 4.427862143e-01 leta0 = -2.341954748e-07 weta0 = -1.889953011e-07 peta0 = 1.923668781e-13
+ etab = 9.900491778e-01 letab = -5.523804145e-07 wetab = -8.027195996e-06 petab = 4.479039809e-12
+ u0 = 1.651954114e-02 lu0 = -7.058219339e-09 wu0 = -1.745402941e-08 pu0 = 1.180491445e-14
+ ua = 2.932745469e-09 lua = -3.418274147e-15 wua = -9.285367985e-15 pua = 8.471752808e-21
+ ub = -3.053990933e-18 lub = 3.599280261e-24 wub = 1.057316628e-23 pub = -1.021968673e-29
+ uc = -1.685344948e-10 luc = 1.053505179e-16 wuc = 2.976757741e-16 puc = -2.510975158e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.587197791e+05 lvsat = 3.600753351e-01 wvsat = 9.611637356e-01 pvsat = -1.063127927e-6
+ a0 = 7.504815302e-01 la0 = 3.613293525e-07 wa0 = 1.371566786e-06 pa0 = -1.119407408e-12
+ ags = 2.527378569e-01 lags = 3.496801486e-07 wags = -1.240158315e-06 pags = 1.300631792e-12
+ a1 = 0.0
+ a2 = 1.039742425e+00 la2 = -2.536882418e-07 wa2 = -1.350532732e-06 pa2 = 1.429093221e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.253200420e-02 lketa = 9.774532041e-10 wketa = 9.706953398e-08 pketa = -1.130892532e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.447195361e-01 lpclm = -7.180195304e-08 wpclm = -3.467512575e-07 ppclm = 5.087440768e-13
+ pdiblc1 = 1.392017393e+00 lpdiblc1 = -1.047257318e-06 wpdiblc1 = -5.026526335e-06 ppdiblc1 = 5.222165562e-12
+ pdiblc2 = -1.840832191e-03 lpdiblc2 = 2.402926499e-09 wpdiblc2 = 4.710589924e-09 ppdiblc2 = -4.984604940e-15
+ pdiblcb = 1.516004117e-02 lpdiblcb = -4.249615076e-08 wpdiblcb = -1.974637899e-07 ppdiblcb = 2.089502586e-13
+ drout = 2.415371047e-01 ldrout = 4.379497494e-08 wdrout = 2.246709322e-06 pdrout = -1.937586553e-13
+ pscbe1 = 7.857608230e+08 lpscbe1 = 1.506746996e+01 wpscbe1 = 7.001292279e+01 ppscbe1 = -7.408557451e-5
+ pscbe2 = 8.786192871e-09 lpscbe2 = 3.276179372e-16 wpscbe2 = 1.626304525e-15 ppscbe2 = -1.128533329e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.360038060e-05 lalpha0 = -4.108146862e-11 walpha0 = -2.146862777e-10 palpha0 = 1.198314396e-16
+ alpha1 = -4.202939353e-10 lalpha1 = 2.904124659e-16 walpha1 = 1.517656826e-15 palpha1 = -8.471105107e-22
+ beta0 = 1.087390033e+02 lbeta0 = -5.569479036e-05 wbeta0 = -2.926704900e-04 pbeta0 = 1.638872439e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 2.209724606e+09 lbgidl = -6.086362661e+02 wbgidl = -2.693406007e+03 pbgidl = 1.627670325e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.915139744e-01 lkt1 = 1.870292095e-10 wkt1 = 1.168858397e-07 pkt1 = -6.563471535e-14
+ kt2 = -1.105091564e-01 lkt2 = 5.346428492e-08 wkt2 = 2.466500083e-07 pkt2 = -1.912006018e-13
+ at = 1.683339169e+05 lat = -5.294882155e-02 wat = 2.875398874e-02 pat = -7.868809534e-8
+ ute = -7.191685180e+00 lute = 3.879517991e-06 wute = 2.104271025e-05 pute = -1.138516526e-11
+ ua1 = -1.282986261e-08 lua1 = 8.853983281e-15 wua1 = 4.525946745e-14 pua1 = -2.669745014e-20
+ ub1 = 8.423991597e-18 lub1 = -5.980879183e-24 wub1 = -2.750562556e-23 pub1 = 1.635829694e-29
+ uc1 = 8.571919036e-10 luc1 = -6.709669257e-16 wuc1 = -2.866547390e-15 puc1 = 2.047204517e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.24 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.179016593e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.661711554e-08 wvth0 = 4.364520526e-07 pvth0 = -1.492880700e-13
+ k1 = -2.900360589e-01 lk1 = 3.619083023e-07 wk1 = 2.123868972e-06 pk1 = -8.423649635e-13
+ k2 = 3.102580745e-01 lk2 = -1.375085524e-07 wk2 = -8.309710901e-07 pk2 = 3.315827639e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.098762963e+00 ldsub = -5.512652301e-08 wdsub = 1.200354982e-06 pdsub = -6.700021404e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.601838373e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.161174089e-08 wvoff = 4.234920439e-07 pvoff = -1.136885844e-13
+ nfactor = {-1.607109764e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.972910306e-07 wnfactor = 6.766877167e-06 pnfactor = -1.404662062e-12
+ eta0 = -5.521951740e-01 leta0 = 3.211732868e-07 weta0 = 3.475014837e-07 peta0 = -1.070895322e-13
+ etab = 1.711765137e-03 letab = -7.201209122e-10 wetab = -6.000721372e-09 petab = 1.849242305e-15
+ u0 = 5.182048296e-03 lu0 = -7.299709582e-10 wu0 = -1.001343503e-09 pu0 = 2.621518758e-15
+ ua = -4.391920263e-09 lua = 6.701345249e-16 wua = 1.058022928e-14 pua = -2.616627618e-21
+ ub = 5.515942687e-18 lub = -1.184199588e-24 wub = -1.623210941e-23 pub = 4.742214000e-30
+ uc = 5.107680032e-11 luc = -1.722991864e-17 wuc = -2.869411162e-16 puc = 7.521809387e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.934587985e+05 lvsat = -2.272191816e-01 wvsat = -2.298521687e+00 pvsat = 7.563306858e-7
+ a0 = 2.260502510e+00 la0 = -4.815190576e-07 wa0 = -1.695490612e-06 pa0 = 5.925320203e-13
+ ags = 8.133875342e-02 lags = 4.453499862e-07 wags = -2.120775717e-07 pags = 7.267879639e-13
+ a1 = 0.0
+ a2 = 3.205151502e-01 la2 = 1.477628462e-07 wa2 = 2.701065464e-06 pa2 = -8.323873440e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.591793694e-01 lketa = -9.486668418e-08 wketa = -5.282530433e-07 pketa = 2.359470498e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 3.676047941e-01 lpclm = 8.287518249e-08 wpclm = 1.253405593e-06 ppclm = -3.844154727e-13
+ pdiblc1 = -1.376418124e+00 lpdiblc1 = 4.980003344e-07 wpdiblc1 = 9.170839433e-06 ppdiblc1 = -2.702378089e-12
+ pdiblc2 = -5.938061315e-03 lpdiblc2 = 4.689876880e-09 wpdiblc2 = -4.876268074e-09 ppdiblc2 = 3.664915888e-16
+ pdiblcb = -1.053200823e-01 lpdiblcb = 2.475223977e-08 wpdiblcb = 3.949275799e-07 ppdiblcb = -1.217048323e-13
+ drout = 1.564118531e-01 ldrout = 9.130933664e-08 wdrout = 4.292581550e-06 pdrout = -1.335703157e-12
+ pscbe1 = 8.282134639e+08 lpscbe1 = -8.628320626e+00 wpscbe1 = -1.387234013e+02 ppscbe1 = 4.242477951e-5
+ pscbe2 = 3.433023715e-08 lpscbe2 = -1.393030126e-14 wpscbe2 = -7.284565351e-14 ppscbe2 = 4.043947949e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.947973579e+00 lbeta0 = 5.568707007e-09 wbeta0 = 3.005331394e-06 pbeta0 = -1.150129371e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 7.368785305e+08 lbgidl = 2.134622282e+02 wbgidl = 1.898396615e+03 pbgidl = -9.353361436e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.288821038e-01 lkt1 = 2.104479796e-08 wkt1 = 1.003603565e-07 pkt1 = -5.641068644e-14
+ kt2 = -8.220387129e-04 lkt2 = -7.759773584e-09 wkt2 = -1.281682853e-07 pkt2 = 1.801172510e-14
+ at = 1.298390884e+05 lat = -3.146216308e-02 wat = -3.085421062e-01 pat = 1.095804660e-7
+ ute = -4.568363194e-01 lute = 1.203274026e-07 wute = 1.202304842e-06 pute = -3.108461760e-13
+ ua1 = 6.243779074e-09 lua1 = -1.792351300e-15 wua1 = -1.060343315e-14 pua1 = 4.483545081e-21
+ ub1 = -5.016661917e-18 lub1 = 1.521290389e-24 wub1 = 8.925741787e-24 pub1 = -3.976599375e-30
+ uc1 = -8.219168702e-10 luc1 = 2.662612186e-16 wuc1 = 2.362103121e-15 puc1 = -8.712713388e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.25 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.035492250e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.612781185e-09 wvth0 = -3.822279392e-07 pvth0 = 1.030045431e-13
+ k1 = 1.180947716e+00 lk1 = -9.140476753e-08 wk1 = -4.313821933e-06 pk1 = 1.141538243e-12
+ k2 = -2.184074520e-01 lk2 = 2.541030289e-08 wk2 = 1.632748727e-06 pk2 = -4.276617720e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -1.524710760e+00 ldsub = 7.533493743e-07 wdsub = 6.392503140e-06 pdsub = -2.270066438e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-9.576087721e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -3.905848271e-08 wvoff = -2.464429882e-07 pvoff = 9.276529447e-14
+ nfactor = {2.420542498e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.439105671e-07 wnfactor = -6.884893331e-06 pnfactor = 2.802404053e-12
+ eta0 = 0.49
+ etab = -0.000625
+ u0 = -1.068275278e-02 lu0 = 4.159084789e-09 wu0 = 5.837570561e-08 pu0 = -1.567670647e-14
+ ua = -4.905045786e-09 lua = 8.282644174e-16 wua = 1.445059994e-14 pua = -3.809359743e-21
+ ub = 2.480390315e-18 lub = -2.487334129e-25 wub = -6.814292988e-24 pub = 1.839925512e-30
+ uc = 1.376067059e-10 luc = -4.389583965e-17 wuc = -5.695348853e-16 puc = 1.623050157e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.699839290e+05 lvsat = 1.005019637e-01 wvsat = 9.694590559e-01 pvsat = -2.507629397e-7
+ a0 = -6.833589280e-01 la0 = 4.256907216e-07 wa0 = 4.433202685e-06 pa0 = -1.296147393e-12
+ ags = 2.467194998e+00 lags = -2.898993326e-07 wags = 9.449028838e-06 pags = -2.250475198e-12
+ a1 = 0.0
+ a2 = 2.045548089e+00 la2 = -3.838405545e-07 wa2 = -2.272248611e-06 pa2 = 7.002388543e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -6.771182283e-01 lketa = 1.628551465e-07 wketa = 1.836173969e-06 pketa = -4.926984225e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.877088690e-01 lpclm = -1.082222903e-07 wpclm = -1.972166218e-06 ppclm = 6.096089924e-13
+ pdiblc1 = -2.099629808e-01 lpdiblc1 = 1.385338530e-07 wpdiblc1 = 8.769374312e-07 ppdiblc1 = -1.464463087e-13
+ pdiblc2 = 1.447875873e-02 lpdiblc2 = -1.601974554e-09 wpdiblc2 = -3.733987885e-08 ppdiblc2 = 1.037080252e-14
+ pdiblcb = -3.488722121e-01 lpdiblcb = 9.980769960e-08 wpdiblcb = 2.925825754e-06 ppdiblcb = -9.016517227e-13
+ drout = 1.875340505e+00 ldrout = -4.384129060e-07 wdrout = -6.632997197e-06 pdrout = 2.031232446e-12
+ pscbe1 = 8.038898385e+08 lpscbe1 = -1.132508999e+00 wpscbe1 = -1.323842821e+01 ppscbe1 = 3.754075350e-6
+ pscbe2 = -3.011945132e-08 lpscbe2 = 5.931159238e-15 wpscbe2 = 1.127409965e-13 ppscbe2 = -1.675275844e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.540327341e+00 lbeta0 = 4.393630482e-07 wbeta0 = 1.154051031e-06 pbeta0 = -5.796203013e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.194437432e-09 lagidl = -3.372727835e-16 wagidl = -5.381263488e-15 pagidl = 1.658343969e-21
+ bgidl = 2.431360930e+09 lbgidl = -3.087264128e+02 wbgidl = -3.663404536e+03 pbgidl = 7.786441170e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.082828250e-01 lkt1 = 1.469671823e-08 wkt1 = 3.237782848e-07 pkt1 = -1.252613894e-13
+ kt2 = 8.745660455e-02 lkt2 = -3.496460308e-08 wkt2 = -4.117119058e-07 pkt2 = 1.053913626e-13
+ at = -6.331905703e+04 lat = 2.806338258e-02 wat = 6.501331588e-01 pat = -1.858544904e-7
+ ute = 2.985790387e+00 lute = -9.405868697e-07 wute = -8.510825293e-06 pute = 2.682449138e-12
+ ua1 = 2.958899696e-09 lua1 = -7.800500222e-16 wua1 = 5.761337647e-15 pua1 = -5.595863350e-22
+ ub1 = -3.269955120e-18 lub1 = 9.830077554e-25 wub1 = -4.348302735e-24 pub1 = 1.140629255e-31
+ uc1 = 1.332525179e-10 luc1 = -2.809333177e-17 wuc1 = -1.635290257e-15 puc1 = 3.606053784e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.26 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -3.7585e-8
+ vth0 = {-1.172008839e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.667877485e-08 wvth0 = 3.458577318e-07 pvth0 = -7.542886182e-14
+ k1 = -1.577849075e+00 lk1 = 6.060331578e-07 wk1 = 4.688774931e-06 pk1 = -1.074174153e-12
+ k2 = 8.477523809e-01 lk2 = -2.448279756e-07 wk2 = -1.958398976e-06 pk2 = 4.581659216e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.164796988e+01 ldsub = -2.554151285e-06 wdsub = -2.641402707e-05 pdsub = 5.939144010e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.980482579e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 9.771287970e-09 wvoff = 2.645886504e-09 pvoff = 3.582664922e-14
+ nfactor = {-4.706534052e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.343020291e-06 wnfactor = 3.176539456e-05 pnfactor = -6.859961068e-12
+ eta0 = 2.517672943e+00 leta0 = -5.174013049e-07 weta0 = -2.925344117e-09 peta0 = 7.464600583e-16
+ etab = 4.780589970e-01 letab = -1.221457955e-07 wetab = -1.400257765e-06 petab = 3.573037738e-13
+ u0 = 2.560563108e-02 lu0 = -4.803756682e-09 wu0 = -5.089267071e-08 pu0 = 1.108633963e-14
+ ua = 3.582245044e-09 lua = -1.278318068e-15 wua = -1.254687415e-14 pua = 2.807682810e-21
+ ub = -1.374896395e-18 lub = 7.172661058e-25 wub = 6.974655086e-24 pub = -1.547270924e-30
+ uc = -3.149583487e-10 luc = 6.845200621e-17 wuc = 9.268729439e-16 puc = -2.079484296e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.932548990e+05 lvsat = -1.636311003e-01 wvsat = -6.209029379e-01 pvsat = 1.371508766e-7
+ a0 = 3.800881097e+00 la0 = -6.881680288e-07 wa0 = -1.199011650e-05 pa0 = 2.802075089e-12
+ ags = 1.25
+ a1 = 0.0
+ a2 = -2.564809090e+00 la2 = 7.651866741e-07 wa2 = 7.265414611e-06 pa2 = -1.683505310e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = 9.062933746e-02 lketa = -2.142679241e-08 wketa = -1.843925016e-06 pketa = 4.111848106e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.464425356e-01 lpclm = 1.734544777e-07 wpclm = 4.892031987e-06 ppclm = -1.098416044e-12
+ pdiblc1 = 2.123594041e+00 lpdiblc1 = -4.470316801e-07 wpdiblc1 = 1.747901528e-06 ppdiblc1 = -3.791432014e-13
+ pdiblc2 = 4.198282536e-02 lpdiblc2 = -8.734532314e-09 wpdiblc2 = 4.596431581e-08 ppdiblc2 = -1.014568596e-14
+ pdiblcb = -7.201239412e+00 lpdiblcb = 1.855450271e-06 wpdiblcb = 4.037064207e-05 ppdiblcb = -1.052080323e-11
+ drout = -7.211504163e+00 ldrout = 1.848984392e-06 wdrout = 1.612250075e-05 pdrout = -3.630303495e-12
+ pscbe1 = 7.926408446e+08 lpscbe1 = 1.657061013e+00 wpscbe1 = 2.146608218e+01 ppscbe1 = -4.833517724e-6
+ pscbe2 = -1.159166231e-07 lpscbe2 = 2.824737540e-14 wpscbe2 = 3.657406494e-13 ppscbe2 = -8.250645136e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.838035327e+01 lbeta0 = -2.295325694e-06 wbeta0 = -7.662249576e-06 pbeta0 = 1.628663226e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.296476741e-09 lagidl = 5.294300685e-16 wagidl = 1.178328921e-14 pagidl = -2.603166351e-21
+ bgidl = 7.241694018e+08 lbgidl = 1.048615029e+02 wbgidl = 8.045763402e+02 pbgidl = -3.058728247e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -2.8385e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -8.929959498e-02 lkt1 = -9.116621629e-08 wkt1 = -7.516992731e-07 pkt1 = 1.402273633e-13
+ kt2 = 5.708003139e-01 lkt2 = -1.607951064e-07 wkt2 = -1.712087862e-06 pkt2 = 4.447308767e-13
+ at = -1.267914596e+05 lat = 4.626273209e-02 wat = 1.533028062e-01 pat = -7.234413452e-8
+ ute = -7.340755986e+00 lute = 1.627301147e-06 wute = 2.702447625e-05 pute = -6.193627008e-12
+ ua1 = -1.584574924e-09 lua1 = 3.236303080e-16 wua1 = 1.664394890e-14 pua1 = -3.376444172e-21
+ ub1 = 8.338593780e-19 lub1 = 6.002132087e-27 wub1 = -1.096869036e-23 pub1 = 1.811528772e-30
+ uc1 = 2.826639753e-11 luc1 = -3.309257690e-18 wuc1 = -1.605847066e-16 puc1 = 1.004390507e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.27 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.182614171e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.976890531e-06 wvth0 = 1.691367254e-07 pvth0 = -3.392573191e-12
+ k1 = 4.299462229e-01 lk1 = 1.121935227e-06 wk1 = -1.673547929e-08 pk1 = 3.356830886e-13
+ k2 = 2.564748852e-02 lk2 = -1.143378376e-07 wk2 = 4.106749490e-08 pk2 = -8.237387942e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.723048825e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 9.758826290e-08 wvoff = 1.412132556e-08 pvoff = -2.832479487e-13
+ nfactor = {2.478776459e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.234354893e-05 wnfactor = -2.227684180e-06 pnfactor = 4.468326799e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.518011894e-02 lu0 = -1.353755247e-07 wu0 = -1.085672450e-08 pu0 = 2.177660258e-13
+ ua = 6.122257994e-10 lua = -1.801299866e-14 wua = -1.281082120e-15 pua = 2.569616295e-20
+ ub = 1.292128209e-19 lub = 2.246976360e-24 wub = -8.047285519e-26 pub = 1.614138210e-30
+ uc = -6.524268182e-11 luc = -8.817512999e-16 wuc = -1.319079733e-17 puc = 2.645832552e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.051033532e+05 lvsat = -2.904239548e+00 wvsat = -2.775527719e-01 pvsat = 5.567200683e-6
+ a0 = 9.752137169e-01 la0 = 1.315966555e-05 wa0 = 1.434742398e-06 pa0 = -2.877830693e-11
+ ags = 1.903488730e-01 lags = 5.279544564e-06 wags = 5.107589225e-07 pags = -1.024488930e-11
+ a1 = 0.0
+ a2 = 1.529618211e+00 la2 = -1.463480610e-05 wa2 = -1.398621200e-06 pa2 = 2.805378179e-11
+ b0 = 0.0
+ b1 = 0.0
+ keta = 7.988441311e-02 lketa = -2.228871635e-06 wketa = -2.582165384e-07 pketa = 5.179351224e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.603464417e-01 lpclm = 4.422678188e-06 wpclm = 6.991370082e-07 ppclm = -1.402340896e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 1.276359717e-02 lpdiblc2 = -2.502579166e-07 wpdiblc2 = -2.420583297e-08 ppdiblc2 = 4.855247127e-13
+ pdiblcb = 7.383542121e-03 lpdiblcb = -1.787958139e-07 wpdiblcb = -2.076731321e-08 ppdiblcb = 4.165542988e-13
+ drout = 0.56
+ pscbe1 = 8.019860747e+08 lpscbe1 = -2.352116235e+02 wpscbe1 = -1.939429323e+02 ppscbe1 = 3.890140306e-3
+ pscbe2 = 9.301635052e-09 lpscbe2 = 1.181435198e-15 wpscbe2 = 6.988266527e-16 ppscbe2 = -1.401718380e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -7.979948686e-10 lalpha0 = 1.801213373e-14 walpha0 = 2.619380988e-15 palpha0 = -5.253998916e-20
+ alpha1 = 3.390946632e-10 lalpha1 = -4.795801401e-15 walpha1 = -6.974204832e-16 palpha1 = 1.398897861e-20
+ beta0 = 9.024175078e+00 lbeta0 = -1.208339278e-04 wbeta0 = -1.103292322e-05 pbeta0 = 2.213002496e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 8.848364432e-11 lagidl = 1.152305475e-15
+ bgidl = 4.835789667e+08 lbgidl = 1.035846088e+04 wbgidl = 2.069816010e+03 pbgidl = -4.151672139e-2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.621928927e-01 lkt1 = 1.334448535e-07 wkt1 = 6.993455671e-08 pkt1 = -1.402759227e-12
+ kt2 = -0.037961
+ at = 0.0
+ ute = -1.733362462e-01 lute = -3.136170173e-06 wute = -3.501623254e-07 pute = 7.023615451e-12
+ ua1 = 2.139515952e-09 lua1 = 7.212597973e-15
+ ub1 = -2.667259284e-19 lub1 = -2.836373812e-23 wub1 = -8.879590665e-25 pub1 = 1.781083391e-29
+ uc1 = 4.311997794e-11 luc1 = 7.677465592e-15 puc1 = -3.308722450e-36
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.28 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.0840563+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.4858803
+ k2 = 0.019947176
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.16743962+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.3648389+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0084309726
+ ua = -2.8581219e-10
+ ub = 2.4123582e-19
+ uc = -1.0920239e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 160312.5
+ a0 = 1.6312888
+ ags = 0.45356055
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.031235975
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.060146165
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00028698955
+ pdiblcb = -0.0015303226
+ drout = 0.56
+ pscbe1 = 790259600.0
+ pscbe2 = 9.3605355e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.4593183e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.45554
+ kt2 = -0.037961
+ at = 0.0
+ ute = -0.32969
+ ua1 = 2.4991e-9
+ ub1 = -1.6808e-18
+ uc1 = 4.2588e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.29 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.099435851e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.239310382e-7
+ k1 = 4.517138262e-01 lk1 = 2.753192546e-7
+ k2 = 2.896633464e-02 lk2 = -7.267791362e-08 wk2 = 2.775557562e-23
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.863612130e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.524734131e-7
+ nfactor = {6.023470053e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.144289311e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.071769316e-02 lu0 = -1.842678302e-8
+ ua = 3.672019860e-10 lua = -5.262099242e-15 pua = 1.654361225e-36
+ ub = -1.759105254e-19 lub = 3.361436166e-24
+ uc = -1.429063055e-10 luc = 2.715918809e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.223167722e+05 lvsat = -4.996409658e-1
+ a0 = 1.662786286e+00 la0 = -2.538121004e-7
+ ags = 4.597325700e-01 lags = -4.973518661e-8
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.754336036e-02 lketa = 5.082598348e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.208481702e-01 lpclm = 4.681751122e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 3.600260080e-04 lpdiblc2 = -5.885401950e-10 wpdiblc2 = -4.336808690e-25
+ pdiblcb = -4.271034041e-04 lpdiblcb = -8.889927828e-9
+ drout = 0.56
+ pscbe1 = 7.803775502e+08 lpscbe1 = 7.963123697e+1
+ pscbe2 = 9.149402307e-09 lpscbe2 = 1.701347163e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -7.459246606e-01 lbeta0 = 3.018529772e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.925316236e-10 lagidl = -3.755090591e-16
+ bgidl = 7.988221066e+08 lbgidl = 1.621125665e+3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.110862019e-01 lkt1 = 4.476007376e-7
+ kt2 = -3.127516493e-02 lkt2 = -5.387559563e-8
+ at = -1.820190699e+05 lat = 1.466740609e+0
+ ute = 1.702663986e-01 lute = -4.028733652e-6
+ ua1 = 5.377245473e-09 lua1 = -2.319258550e-14
+ ub1 = -4.268705154e-18 lub1 = 2.085377968e-23
+ uc1 = 7.964315027e-10 luc1 = -2.985967003e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.30 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.039182268e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.205882467e-7
+ k1 = 6.004806109e-01 lk1 = -3.284016481e-7
+ k2 = -6.050885308e-03 lk2 = 6.942791788e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.208171143e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.135156818e-7
+ nfactor = {2.996480249e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.571510395e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 4.093373681e-03 lu0 = 8.455831565e-9
+ ua = -1.478847421e-09 lua = 2.229483078e-15
+ ub = 1.027860336e-18 lub = -1.523670633e-24
+ uc = -6.663496362e-11 luc = -3.793019065e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.462869005e+05 lvsat = -1.910988216e-1
+ a0 = 2.032959356e+00 la0 = -1.756037345e-6
+ ags = 5.622897495e-01 lags = -4.659296555e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -4.174605632e-02 lketa = 6.788123813e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.441032208e-01 lpclm = -1.263270664e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000215
+ pdiblcb = 2.041553198e-02 lpdiblcb = -9.347288545e-08 ppdiblcb = 2.081668171e-29
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.696808226e-08 lpscbe2 = -3.002818526e-14 ppscbe2 = -2.646977960e-35
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.526703342e+00 lbeta0 = 4.729906941e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.141087571e+09 lbgidl = 2.321542270e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.414871760e-01 lkt1 = -2.406609414e-7
+ kt2 = -4.002107588e-02 lkt2 = -1.838320215e-8
+ at = 2.779140841e+05 lat = -3.997463191e-01 pat = 4.656612873e-22
+ ute = -1.668881831e+00 lute = 3.434842518e-6
+ ua1 = -3.376869106e-09 lua1 = 1.233309966e-14 wua1 = 8.271806126e-31 pua1 = -4.963083675e-36
+ ub1 = 3.250298115e-18 lub1 = -9.659613820e-24 wub1 = -1.540743956e-39
+ uc1 = 9.326290009e-11 luc1 = -1.323892745e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.31 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.103865560e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.254096557e-8
+ k1 = 4.316923847e-01 lk1 = 1.899321537e-8
+ k2 = 3.069529095e-02 lk2 = -6.201959716e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 3.798690224e-01 ldsub = 3.707401741e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.831729372e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.482320221e-8
+ nfactor = {8.628159584e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.199334386e-7
+ eta0 = -6.708088940e-02 leta0 = 3.027174741e-7
+ etab = 7.371527644e-01 letab = -1.661257605e-06 wetab = -2.220446049e-22 petab = 5.551115123e-28
+ u0 = 8.743169528e-03 lu0 = -1.114238755e-9
+ ua = -3.520491852e-11 lua = -7.417786107e-16
+ ub = -1.078331476e-19 lub = 8.137796256e-25
+ uc = -1.239932619e-10 luc = 8.012293822e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.946698149e+04 lvsat = 2.875473117e-2
+ a0 = 1.158873009e+00 la0 = 4.298095092e-8
+ ags = 7.823807504e-02 lags = 5.303309793e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.199495869e-03 lketa = -1.351230619e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.081281139e-02 lpclm = 6.370179576e-7
+ pdiblc1 = 4.101224041e-01 lpdiblc1 = -4.141532844e-8
+ pdiblc2 = -1.250655000e-05 lpdiblc2 = 4.682471560e-10
+ pdiblcb = -0.025
+ drout = 1.045812717e-01 ldrout = 9.373291640e-7
+ pscbe1 = 800000000.0
+ pscbe2 = -4.932972695e-09 lpscbe2 = 1.504790901e-14 ppscbe2 = 3.308722450e-36
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.722141263e+00 lbeta0 = 2.269492475e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.270154104e+09 lbgidl = -3.348664091e+1
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.434825322e-01 lkt1 = -3.073715895e-8
+ kt2 = -6.120850883e-02 lkt2 = 2.522413672e-8
+ at = 6.361637926e+04 lat = 4.131478816e-2
+ ute = 0.0
+ ua1 = 2.838982471e-09 lua1 = -4.601795842e-16
+ ub1 = -1.532952888e-18 lub1 = 1.851298980e-25
+ uc1 = 1.615321807e-10 luc1 = -2.728990597e-16 wuc1 = 5.169878828e-32 puc1 = 5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.32 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.132799035e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.315750087e-8
+ k1 = 3.162982928e-01 lk1 = 1.410997816e-7
+ k2 = 7.189253146e-02 lk2 = -4.979564370e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 4.290723551e-01 ldsub = 3.186746836e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.749039384e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 6.073195684e-9
+ nfactor = {2.038727531e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.243809106e-7
+ eta0 = 3.779934975e-01 leta0 = -1.682468899e-7
+ etab = -1.761891394e+00 letab = 9.831559518e-7
+ u0 = 1.053582632e-02 lu0 = -3.011174388e-9
+ ua = -2.505305958e-10 lua = -5.139274387e-16
+ ub = 5.707773262e-19 lub = 9.569438051e-26
+ uc = -6.648316323e-11 luc = 1.926747706e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.079322663e+04 lvsat = -4.393761653e-3
+ a0 = 1.220691836e+00 la0 = -2.243387722e-8
+ ags = -1.724220597e-01 lags = 7.955720141e-7
+ a1 = 0.0
+ a2 = 5.767431634e-01 la2 = 2.362436868e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.074606562e-02 lketa = -3.779261099e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.258437974e-01 lpclm = 1.026093191e-7
+ pdiblc1 = -3.312122082e-01 lpdiblc1 = 7.430427182e-07 ppdiblc1 = -4.440892099e-28
+ pdiblc2 = -2.259141628e-04 lpdiblc2 = 6.940686897e-10
+ pdiblcb = -5.253590337e-02 lpdiblcb = 2.913766687e-8
+ drout = 1.011770015e+00 ldrout = -2.263074892e-8
+ pscbe1 = 8.097631524e+08 lpscbe1 = -1.033107499e+1
+ pscbe2 = 9.343734185e-09 lpscbe2 = -5.927390603e-17
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.403618953e+00 lbeta0 = 4.902032285e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.286351953e+09 lbgidl = -5.062671849e+1
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.514423374e-01 lkt1 = -2.231433193e-8
+ kt2 = -2.595084180e-02 lkt2 = -1.208446880e-8
+ at = 1.781915644e+05 lat = -7.992523550e-2
+ ute = 2.232680000e-02 lute = -2.362554996e-8
+ ua1 = 2.686310752e-09 lua1 = -2.986269514e-16
+ ub1 = -1.005683096e-18 lub1 = -3.728111783e-25
+ uc1 = -1.255383132e-10 luc1 = 3.087032485e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.33 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.029388988e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.456288516e-8
+ k1 = 4.380838471e-01 lk1 = 7.312273876e-8
+ k2 = 2.537863995e-02 lk2 = -2.383298488e-08 pk2 = 1.387778781e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.510277217e+00 ldsub = -2.848214344e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.149992750e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.736379029e-8
+ nfactor = {7.127593194e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.157347663e-7
+ eta0 = -4.330622374e-01 leta0 = 2.844600897e-07 weta0 = 1.110223025e-22 peta0 = -1.110223025e-28
+ etab = -3.454449539e-04 letab = -8.615047856e-11
+ u0 = 4.838760576e-03 lu0 = 1.687567961e-10
+ ua = -7.647306152e-10 lua = -2.269164139e-16
+ ub = -4.886480987e-20 lub = 4.415600316e-25
+ uc = -4.729439924e-11 luc = 8.556884661e-18 wuc = 5.169878828e-32
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.463203500e+03 lvsat = 3.207149736e-2
+ a0 = 1.679242328e+00 la0 = -2.783830052e-7
+ ags = 8.632808000e-03 lags = 6.945126186e-7
+ a1 = 0.0
+ a2 = 1.246513673e+00 la2 = -1.376021187e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.192010580e-02 lketa = -1.397763409e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 7.973062374e-01 lpclm = -4.891287104e-8
+ pdiblc1 = 1.767594446e+00 lpdiblc1 = -4.284481920e-7
+ pdiblc2 = -7.609778308e-03 lpdiblc2 = 4.815520140e-09 wpdiblc2 = -1.734723476e-24 ppdiblc2 = 8.673617380e-31
+ pdiblcb = 3.007180675e-02 lpdiblcb = -1.697147869e-08 wpdiblcb = 1.127570259e-23 ppdiblcb = -1.951563910e-30
+ drout = 1.628025270e+00 ldrout = -3.666059441e-7
+ pscbe1 = 7.806553182e+08 lpscbe1 = 5.916044807e+0
+ pscbe2 = 9.356770764e-09 lpscbe2 = -6.655053296e-17
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.978282718e+00 lbeta0 = -3.887268453e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.387700395e+09 lbgidl = -1.071963782e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.944758507e-01 lkt1 = 1.705684185e-9
+ kt2 = -4.476160421e-02 lkt2 = -1.584865548e-9
+ at = 2.406248337e+04 lat = 6.104993660e-3
+ ute = -4.465360000e-02 lute = 1.376089991e-8
+ ua1 = 2.608634511e-09 lua1 = -2.552704041e-16
+ ub1 = -1.956675470e-18 lub1 = 1.580042353e-25
+ uc1 = -1.212383460e-11 luc1 = -3.243423468e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.34 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.166530656e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.770006249e-08 wvth0 = 8.680776169e-13 pvth0 = -2.675154791e-19
+ k1 = -2.979473149e-01 lk1 = 2.999454619e-07 wk1 = -4.830962759e-13 pk1 = 1.488757793e-19
+ k2 = 3.413432603e-01 lk2 = -1.212038019e-07 wk2 = -4.407692606e-13 pk2 = 1.358318629e-19
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 6.668127176e-01 ldsub = -2.489097951e-08 wdsub = 9.437577653e-14 pdsub = -2.908378294e-20
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.802482028e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.256028214e-09 wvoff = -4.965571776e-14 pvoff = 1.530240268e-20
+ nfactor = {6.021415600e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.168296093e-07 wnfactor = 3.380179052e-13 pnfactor = -1.041669790e-19
+ eta0 = 0.49
+ etab = -0.000625
+ u0 = 9.330025161e-03 lu0 = -1.215316211e-09 wu0 = -6.640704098e-15 pu0 = 2.046465782e-21
+ ua = 4.901202858e-11 lua = -4.776874844e-16 wua = -2.931482960e-22 pua = 9.033951151e-29
+ ub = 1.442659296e-19 lub = 3.820429316e-25 wub = -3.741528940e-31 pub = 1.153026971e-37
+ uc = -5.764530464e-11 luc = 1.174672318e-17 wuc = -8.973958388e-26 puc = 2.765506480e-32
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.237295108e+04 lvsat = 1.453362044e-02 wvsat = -3.941697534e-08 pvsat = 1.214712916e-14
+ a0 = 8.364632238e-01 la0 = -1.866376866e-08 wa0 = 1.405915384e-14 pa0 = -4.332609826e-21
+ ags = 5.706578265e+00 lags = -1.061423233e-06 wags = 5.189918895e-13 pags = -1.599377306e-19
+ a1 = 0.0
+ a2 = 1.266559229e+00 la2 = -1.437795575e-07 wa2 = 1.133107531e-12 pa2 = -3.491897465e-19
+ b0 = 0.0
+ b1 = 0.0
+ keta = -4.762797474e-02 lketa = -6.055240113e-09 wketa = -7.478275776e-16 pketa = 2.304580415e-22
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 3.115967848e-01 lpclm = 1.007682110e-07 wpclm = -4.935660769e-15 ppclm = 1.521022419e-21
+ pdiblc1 = 9.067498340e-02 lpdiblc1 = 8.832807881e-08 wpdiblc1 = -6.057398672e-14 ppdiblc1 = 1.866708566e-20
+ pdiblc2 = 1.677635450e-03 lpdiblc2 = 1.953417842e-09 wpdiblc2 = -7.268879387e-16 ppdiblc2 = 2.240050576e-22
+ pdiblcb = 6.541801203e-01 lpdiblcb = -2.093029377e-07 wpdiblcb = 3.389152086e-13 ppdiblcb = -1.044434999e-19
+ drout = -3.986309342e-01 ldrout = 2.579486982e-07 wdrout = 1.217462398e-13 pdrout = -3.751853939e-20
+ pscbe1 = 7.993513496e+08 lpscbe1 = 1.544888388e-01 wpscbe1 = -9.871315002e-06 ppscbe1 = 3.042043686e-12
+ pscbe2 = 8.531220678e-09 lpscbe2 = 1.878592369e-16 wpscbe2 = 1.012557796e-21 ppscbe2 = -3.120399299e-28
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.935967157e+00 lbeta0 = 2.406535410e-07 wbeta0 = 5.459137640e-13 pbeta0 = -1.682342443e-19
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -6.504056172e-10 lagidl = 2.312524990e-16 wagidl = -2.108872347e-22 pagidl = 6.498911873e-29
+ bgidl = 1.175446303e+09 lbgidl = -4.178603485e+01 wbgidl = 4.681397247e-04 pbgidl = -1.442666187e-10
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.00081386752815302
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207367379934e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.972827986e-01 lkt1 = -2.824629868e-08 wkt1 = -1.343097296e-13 pkt1 = 4.139022947e-20
+ kt2 = -5.368940352e-02 lkt2 = 1.166414366e-09 wkt2 = -9.624533615e-15 pkt2 = 2.965992507e-21
+ at = 1.595642032e+05 lat = -3.565257133e-02 wat = 7.373574679e-08 pat = -2.272314514e-14
+ ute = 6.804857687e-02 lute = -2.097052994e-08 wute = -1.588384718e-14 pute = 4.894925187e-21
+ ua1 = 4.934042916e-09 lua1 = -9.718915122e-16 wua1 = -1.063410055e-21 pua1 = 3.277110750e-28
+ ub1 = -4.760671593e-18 lub1 = 1.022111720e-24 wub1 = 9.422620943e-31 pub1 = -2.903769120e-37
+ uc1 = -4.273693199e-10 luc1 = 9.553196652e-17 wuc1 = -8.450445622e-23 puc1 = 2.604173824e-29
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.35 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -3.7585e-8
+ vth0 = {-1.053438633e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.195347515e-10 wvth0 = -2.310718486e-12 pvth0 = 5.245233119e-19
+ k1 = 2.959003898e-02 lk1 = 2.377771388e-07 wk1 = 4.146701045e-13 pk1 = -6.958087262e-20
+ k2 = 1.763597441e-01 lk2 = -8.775619308e-08 wk2 = 9.772795266e-13 pk2 = -2.163162951e-19
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.592524967e+00 ldsub = -5.180516323e-07 wdsub = -5.689937588e-13 pdsub = 1.381122914e-19
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.971411873e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.205363687e-08 wvoff = 3.223197531e-14 pvoff = -4.500630979e-21
+ nfactor = {6.183503667e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.008760125e-06 wnfactor = 3.956690620e-12 pnfactor = -1.034978883e-18
+ eta0 = 2.516669947e+00 leta0 = -5.171453704e-07 weta0 = 3.173815486e-13 peta0 = -8.098624971e-20
+ etab = -1.987355131e-03 letab = 3.476321587e-10 wetab = 1.088014248e-15 petab = -2.776285955e-22
+ u0 = 8.158236193e-03 lu0 = -1.003057159e-09 wu0 = 1.928223645e-14 pu0 = -4.422219160e-21
+ ua = -7.191628324e-10 lua = -3.157684853e-16 wua = -2.879780082e-21 pua = 7.568185617e-28
+ ub = 1.016204300e-18 lub = 1.868197203e-25 wub = 8.648478087e-31 pub = -1.926230821e-37
+ uc = 2.798840580e-12 luc = -2.838356597e-18 wuc = 7.787041477e-24 puc = -1.980289244e-30
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.803922899e+05 lvsat = -1.166119995e-01 wvsat = 6.895976840e-07 pvsat = -1.730085083e-13
+ a0 = -3.096564702e-01 la0 = 2.724594189e-07 wa0 = 9.631694056e-13 pa0 = -2.468263194e-19
+ ags = 1.250000445e+00 lags = -1.001533834e-13 wags = -1.297417981e-12 pags = 2.921396067e-19
+ a1 = 0.0
+ a2 = -7.402697799e-02 la2 = 1.880351869e-07 wa2 = -2.529967301e-12 pa2 = 5.605927367e-19
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.415183716e-01 lketa = 1.195385640e-07 wketa = 5.443786768e-13 pketa = -1.388530224e-19
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.530678399e+00 lpclm = -2.031122527e-07 wpclm = 1.037176027e-12 ppclm = -2.642860517e-19
+ pdiblc1 = 2.722822646e+00 lpdiblc1 = -5.770123950e-07 wpdiblc1 = -1.571613858e-12 ppdiblc1 = 4.055715426e-19
+ pdiblc2 = 5.774061431e-02 lpdiblc2 = -1.221274222e-08 wpdiblc2 = 7.454702389e-14 ppdiblc2 = -1.896765008e-20
+ pdiblcb = 6.638917389e+00 lpdiblcb = -1.751367885e-06 wpdiblcb = -1.578673689e-11 ppdiblcb = 4.002884220e-18
+ drout = -1.684274215e+00 ldrout = 6.044180500e-07 wdrout = 2.120507261e-12 pdrout = -5.502203733e-19
+ pscbe1 = 7.999999915e+08 lpscbe1 = 1.904934883e-06 wpscbe1 = 2.467712402e-05 ppscbe1 = -5.556547165e-12
+ pscbe2 = 9.469195193e-09 lpscbe2 = -3.807478098e-17 wpscbe2 = -2.449329333e-21 ppscbe2 = 5.490571458e-28
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.575352607e+01 lbeta0 = -1.736975698e-06 wbeta0 = 4.706656114e-13 pbeta0 = -1.610413278e-19
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.743154854e-09 lagidl = -3.630060808e-16 wagidl = -1.059802806e-21 pagidl = 2.862456731e-28
+ bgidl = 1.000000401e+09 lbgidl = -9.034009647e-05 wbgidl = -1.170293617e-03 pbgidl = 2.635150146e-10
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -2.8385e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.00081386752815302
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207367379934e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.470026340e-01 lkt1 = -4.309244094e-08 wkt1 = 3.908287027e-13 pkt1 = -8.965501053e-20
+ kt2 = -1.614990125e-02 lkt2 = -8.329284585e-09 wkt2 = 1.329673434e-13 pkt2 = -3.320747144e-20
+ at = -7.423509248e+04 lat = 2.146120041e-02 wat = -1.726912934e-08 pat = -1.123354145e-15
+ ute = 1.923967872e+00 lute = -4.960422823e-07 wute = -5.991085649e-13 pute = 1.540657640e-19
+ ua1 = 4.121420959e-09 lua1 = -8.339060390e-16 wua1 = 3.978325149e-21 pua1 = -9.353972706e-28
+ ub1 = -2.926504077e-18 lub1 = 6.270430641e-25 wub1 = -3.470167355e-30 pub1 = 8.148163087e-37
+ uc1 = -2.678646886e-11 luc1 = 1.340817170e-19 wuc1 = 2.105902421e-22 puc1 = -4.739877946e-29
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.36 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.094380677e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.070881130e-7
+ k1 = 4.212158315e-01 lk1 = 1.297050901e-6
+ k2 = 4.707115360e-02 lk2 = -5.440573537e-7
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.649382158e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.017359110e-8
+ nfactor = {1.316661266e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 9.663551657e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 9.516495432e-03 lu0 = -2.177360149e-8
+ ua = -5.607584256e-11 lua = -4.608090712e-15 pua = 3.308722450e-36
+ ub = 8.723257589e-20 lub = 3.089023251e-24
+ uc = -7.212392024e-11 luc = -7.437262497e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 160312.5
+ a0 = 1.723675260e+00 la0 = -1.853103320e-6
+ ags = 4.567962936e-01 lags = -6.490309596e-8
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.481931420e-02 lketa = 4.730386269e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.043721062e-01 lpclm = -2.892908447e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 1.361491196e-04 lpdiblc2 = 3.025582995e-9
+ pdiblcb = -3.450134580e-03 lpdiblcb = 3.850791507e-8
+ drout = 0.56
+ pscbe1 = 7.008119360e+08 lpscbe1 = 1.794156450e+3
+ pscbe2 = 9.666191697e-09 lpscbe2 = -6.130903958e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 5.684566553e-10 lalpha0 = -9.396383230e-15
+ alpha1 = -2.472842568e-11 lalpha1 = 2.501823966e-15 walpha1 = -1.817535526e-32 palpha1 = 7.108583389e-37
+ beta0 = 3.268634049e+00 lbeta0 = -5.388307414e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 8.848364432e-11 lagidl = 1.152305475e-15
+ bgidl = 1.563339129e+09 lbgidl = -1.129955201e+4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.257101581e-01 lkt1 = -5.983320405e-7
+ kt2 = -0.037961
+ at = 0.0
+ ute = -3.560052987e-01 lute = 5.278367351e-7
+ ua1 = 2.139515952e-09 lua1 = 7.212597973e-15
+ ub1 = -7.299472105e-19 lub1 = -1.907236690e-23 wub1 = 1.540743956e-39
+ uc1 = 4.311997794e-11 luc1 = 7.677465592e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.37 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.0840563+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.4858803
+ k2 = 0.019947176
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.16743962+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.3648389+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0084309726
+ ua = -2.8581219e-10
+ ub = 2.4123582e-19
+ uc = -1.0920239e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 160312.5
+ a0 = 1.6312888
+ ags = 0.45356055
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.031235975
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.060146165
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00028698955
+ pdiblcb = -0.0015303226
+ drout = 0.56
+ pscbe1 = 790259600.0
+ pscbe2 = 9.3605355e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.4593183e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.45554
+ kt2 = -0.037961
+ at = 0.0
+ ute = -0.32969
+ ua1 = 2.4991e-9
+ ub1 = -1.6808e-18
+ uc1 = 4.2588e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.38 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.099435851e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.239310382e-7
+ k1 = 4.517138262e-01 lk1 = 2.753192546e-7
+ k2 = 2.896633464e-02 lk2 = -7.267791362e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.863612130e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.524734131e-7
+ nfactor = {6.023470053e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.144289311e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.071769316e-02 lu0 = -1.842678302e-8
+ ua = 3.672019860e-10 lua = -5.262099242e-15
+ ub = -1.759105254e-19 lub = 3.361436166e-24
+ uc = -1.429063055e-10 luc = 2.715918809e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.223167722e+05 lvsat = -4.996409658e-1
+ a0 = 1.662786286e+00 la0 = -2.538121004e-7
+ ags = 4.597325700e-01 lags = -4.973518661e-8
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.754336036e-02 lketa = 5.082598348e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.208481702e-01 lpclm = 4.681751122e-06 wpclm = -2.220446049e-22 ppclm = -2.664535259e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 3.600260080e-04 lpdiblc2 = -5.885401950e-10
+ pdiblcb = -4.271034041e-04 lpdiblcb = -8.889927828e-9
+ drout = 0.56
+ pscbe1 = 7.803775502e+08 lpscbe1 = 7.963123697e+1
+ pscbe2 = 9.149402307e-09 lpscbe2 = 1.701347163e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -7.459246606e-01 lbeta0 = 3.018529772e-05 pbeta0 = 2.842170943e-26
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.925316236e-10 lagidl = -3.755090591e-16
+ bgidl = 7.988221066e+08 lbgidl = 1.621125665e+3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.110862019e-01 lkt1 = 4.476007376e-7
+ kt2 = -3.127516492e-02 lkt2 = -5.387559563e-8
+ at = -1.820190699e+05 lat = 1.466740609e+0
+ ute = 1.702663986e-01 lute = -4.028733652e-6
+ ua1 = 5.377245473e-09 lua1 = -2.319258550e-14
+ ub1 = -4.268705154e-18 lub1 = 2.085377968e-23 pub1 = -2.465190329e-44
+ uc1 = 7.964315027e-10 luc1 = -2.985967003e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.39 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.039182268e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.205882467e-7
+ k1 = 6.004806109e-01 lk1 = -3.284016481e-7
+ k2 = -6.050885308e-03 lk2 = 6.942791788e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.208171143e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.135156818e-7
+ nfactor = {2.996480249e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.571510395e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 4.093373681e-03 lu0 = 8.455831565e-9
+ ua = -1.478847421e-09 lua = 2.229483078e-15
+ ub = 1.027860336e-18 lub = -1.523670633e-24 pub = -3.081487911e-45
+ uc = -6.663496362e-11 luc = -3.793019065e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.462869005e+05 lvsat = -1.910988216e-1
+ a0 = 2.032959356e+00 la0 = -1.756037345e-06 wa0 = -3.552713679e-21
+ ags = 5.622897495e-01 lags = -4.659296555e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -4.174605632e-02 lketa = 6.788123813e-08 wketa = -5.551115123e-23
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.441032208e-01 lpclm = -1.263270664e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000215
+ pdiblcb = 2.041553198e-02 lpdiblcb = -9.347288545e-08 wpdiblcb = -6.938893904e-24 ppdiblcb = -2.775557562e-29
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.696808226e-08 lpscbe2 = -3.002818526e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.526703342e+00 lbeta0 = 4.729906941e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.141087571e+09 lbgidl = 2.321542270e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.414871760e-01 lkt1 = -2.406609414e-7
+ kt2 = -4.002107588e-02 lkt2 = -1.838320215e-8
+ at = 2.779140841e+05 lat = -3.997463191e-1
+ ute = -1.668881831e+00 lute = 3.434842518e-6
+ ua1 = -3.376869106e-09 lua1 = 1.233309966e-14 wua1 = 3.308722450e-30
+ ub1 = 3.250298115e-18 lub1 = -9.659613820e-24 wub1 = 3.081487911e-39
+ uc1 = 9.326290009e-11 luc1 = -1.323892745e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.40 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.103865560e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.254096557e-8
+ k1 = 4.316923847e-01 lk1 = 1.899321537e-8
+ k2 = 3.069529095e-02 lk2 = -6.201959716e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 3.798690224e-01 ldsub = 3.707401741e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.831729372e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.482320221e-8
+ nfactor = {8.628159584e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.199334386e-7
+ eta0 = -6.708088940e-02 leta0 = 3.027174741e-07 peta0 = 2.220446049e-28
+ etab = 7.371527644e-01 letab = -1.661257605e-06 wetab = -2.220446049e-22
+ u0 = 8.743169528e-03 lu0 = -1.114238755e-9
+ ua = -3.520491852e-11 lua = -7.417786107e-16
+ ub = -1.078331476e-19 lub = 8.137796256e-25 pub = -7.703719778e-46
+ uc = -1.239932619e-10 luc = 8.012293822e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.946698149e+04 lvsat = 2.875473117e-2
+ a0 = 1.158873009e+00 la0 = 4.298095092e-8
+ ags = 7.823807504e-02 lags = 5.303309793e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.199495869e-03 lketa = -1.351230619e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.081281139e-02 lpclm = 6.370179576e-7
+ pdiblc1 = 4.101224041e-01 lpdiblc1 = -4.141532844e-8
+ pdiblc2 = -1.250655000e-05 lpdiblc2 = 4.682471560e-10
+ pdiblcb = -0.025
+ drout = 1.045812717e-01 ldrout = 9.373291640e-7
+ pscbe1 = 800000000.0
+ pscbe2 = -4.932972695e-09 lpscbe2 = 1.504790901e-14 ppscbe2 = -1.323488980e-35
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.722141263e+00 lbeta0 = 2.269492475e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.270154104e+09 lbgidl = -3.348664091e+1
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.434825322e-01 lkt1 = -3.073715895e-8
+ kt2 = -6.120850883e-02 lkt2 = 2.522413672e-8
+ at = 6.361637926e+04 lat = 4.131478816e-2
+ ute = 0.0
+ ua1 = 2.838982471e-09 lua1 = -4.601795842e-16
+ ub1 = -1.532952888e-18 lub1 = 1.851298980e-25
+ uc1 = 1.615321807e-10 luc1 = -2.728990597e-16 puc1 = 2.067951531e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.41 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.132799035e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.315750087e-8
+ k1 = 3.162982928e-01 lk1 = 1.410997816e-7
+ k2 = 7.189253146e-02 lk2 = -4.979564370e-08 pk2 = 5.551115123e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 4.290723551e-01 ldsub = 3.186746836e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.749039384e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 6.073195684e-9
+ nfactor = {2.038727531e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.243809106e-7
+ eta0 = 3.779934975e-01 leta0 = -1.682468899e-7
+ etab = -1.761891394e+00 letab = 9.831559518e-7
+ u0 = 1.053582632e-02 lu0 = -3.011174388e-9
+ ua = -2.505305958e-10 lua = -5.139274387e-16
+ ub = 5.707773262e-19 lub = 9.569438051e-26
+ uc = -6.648316323e-11 luc = 1.926747706e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.079322663e+04 lvsat = -4.393761653e-3
+ a0 = 1.220691836e+00 la0 = -2.243387722e-8
+ ags = -1.724220597e-01 lags = 7.955720141e-7
+ a1 = 0.0
+ a2 = 5.767431634e-01 la2 = 2.362436868e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.074606562e-02 lketa = -3.779261099e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.258437974e-01 lpclm = 1.026093191e-7
+ pdiblc1 = -3.312122082e-01 lpdiblc1 = 7.430427182e-7
+ pdiblc2 = -2.259141628e-04 lpdiblc2 = 6.940686897e-10
+ pdiblcb = -5.253590337e-02 lpdiblcb = 2.913766687e-8
+ drout = 1.011770015e+00 ldrout = -2.263074892e-8
+ pscbe1 = 8.097631524e+08 lpscbe1 = -1.033107499e+1
+ pscbe2 = 9.343734185e-09 lpscbe2 = -5.927390603e-17
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.403618953e+00 lbeta0 = 4.902032285e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.286351953e+09 lbgidl = -5.062671849e+1
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.514423374e-01 lkt1 = -2.231433193e-8
+ kt2 = -2.595084180e-02 lkt2 = -1.208446880e-8
+ at = 1.781915644e+05 lat = -7.992523550e-2
+ ute = 2.232680000e-02 lute = -2.362554996e-8
+ ua1 = 2.686310752e-09 lua1 = -2.986269514e-16
+ ub1 = -1.005683096e-18 lub1 = -3.728111783e-25
+ uc1 = -1.255383132e-10 luc1 = 3.087032485e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.42 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-8.668778017e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.052717541e-07 wvth0 = -3.115212686e-07 pvth0 = 1.738818265e-13
+ k1 = 2.197818184e+00 lk1 = -9.091081763e-07 wk1 = -3.373273465e-06 pk1 = 1.882860050e-12
+ k2 = -6.857050043e-01 lk2 = 3.730725728e-07 wk2 = 1.363091882e-06 pk2 = -7.608369955e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.364245581e+00 ldsub = -2.033109558e-07 wdsub = 2.799312569e-07 pdsub = -1.562492297e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.575692294e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -3.602518826e-09 wvoff = 8.160328219e-08 pvoff = -4.554850402e-14
+ nfactor = {3.744918809e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.376725696e-06 wnfactor = -5.812413234e-06 pnfactor = 3.244314695e-12
+ eta0 = -4.330622374e-01 leta0 = 2.844600897e-07 peta0 = 1.110223025e-28
+ etab = -3.454449539e-04 letab = -8.615047856e-11
+ u0 = -2.291306406e-03 lu0 = 4.148546284e-09 wu0 = 1.366778226e-08 pu0 = -7.628946024e-15
+ ua = -3.567249323e-09 lua = 1.337365453e-15 wua = 5.372209766e-15 pua = -2.998606325e-21
+ ub = 2.192522649e-18 lub = -8.095152065e-25 wub = -4.296564931e-24 pub = 2.398213648e-30
+ uc = 2.162181862e-11 luc = -2.991008066e-17 wuc = -1.321070142e-16 puc = 7.373817210e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.072975598e+04 lvsat = -1.552173424e-02 wvsat = -1.634493303e-01 pvsat = 9.123251270e-8
+ a0 = 1.569744855e+00 la0 = -2.172648008e-07 wa0 = 2.098981145e-07 pa0 = -1.171588306e-13
+ ags = -6.218574500e+00 lags = 4.170352922e-06 wags = 1.193707069e-05 pags = -6.662914745e-12
+ a1 = 0.0
+ a2 = 4.029800599e-01 la2 = 3.332330383e-07 wa2 = 1.616988141e-06 pa2 = -9.025542707e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.744526730e-02 lketa = 5.851445310e-09 wketa = 6.809896364e-08 pketa = -3.801079853e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.388497834e+00 lpclm = -3.788982843e-07 wpclm = -1.133268177e-06 ppclm = 6.325562984e-13
+ pdiblc1 = 2.285801753e+00 lpdiblc1 = -7.176959647e-07 wpdiblc1 = -9.933629876e-07 ppdiblc1 = 5.544654188e-13
+ pdiblc2 = 3.850624342e-03 lpdiblc2 = -1.581332808e-09 wpdiblc2 = -2.196869797e-08 ppdiblc2 = 1.226226815e-14
+ pdiblcb = -1.197876649e+00 lpdiblcb = 6.684325109e-07 wpdiblcb = 2.353881410e-06 ppdiblcb = -1.313865987e-12
+ drout = 3.141370484e+00 ldrout = -1.211309843e-06 wdrout = -2.900964736e-06 pdrout = 1.619231487e-12
+ pscbe1 = 7.815616898e+08 lpscbe1 = 5.410135393e+00 wpscbe1 = -1.737443585e+00 ppscbe1 = 9.697888860e-7
+ pscbe2 = 1.045891105e-08 lpscbe2 = -6.817321773e-16 wpscbe2 = -2.112716964e-15 ppscbe2 = 1.179255228e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.139015951e+01 lbeta0 = -1.176794112e-06 wbeta0 = -2.706457676e-06 pbeta0 = 1.510663481e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.456723035e-09 lagidl = -7.572820964e-16 wagidl = -2.600732234e-15 pagidl = 1.451650711e-21
+ bgidl = 1.142547715e+09 lbgidl = 2.964049296e+01 wbgidl = 4.699385650e+02 pbgidl = -2.623056088e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.00081386752815302
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207367379934e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -6.601924130e-01 lkt1 = 9.420369776e-08 wkt1 = 3.176657240e-07 pkt1 = -1.773114772e-13
+ kt2 = -3.791842149e-02 lkt2 = -5.404524849e-09 wkt2 = -1.311784751e-08 pkt2 = 7.321988946e-15
+ at = -1.851057374e+05 lat = 1.228564194e-01 wat = 4.009591641e-01 pat = -2.238033766e-7
+ ute = -1.676844580e-01 lute = 8.243303395e-08 wute = 2.358405585e-07 pute = -1.316391245e-13
+ ua1 = -3.093302472e-09 lua1 = 2.927379762e-15 wua1 = 1.093016845e-14 pua1 = -6.100892122e-21
+ ub1 = 4.039895863e-18 lub1 = -3.189101986e-24 wub1 = -1.149495951e-23 pub1 = 6.416141552e-30
+ uc1 = 5.483475960e-10 luc1 = -3.452725731e-16 wuc1 = -1.074380016e-15 puc1 = 5.996866934e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.43 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.746927297e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.659330990e-07 wvth0 = 1.112575959e-06 pvth0 = -2.649822163e-13
+ k1 = -6.582713057e+00 lk1 = 1.796788136e-06 wk1 = 1.204740523e-05 pk1 = -2.869330504e-12
+ k2 = 2.880927474e+00 lk2 = -7.260565580e-07 wk2 = -4.868185291e-06 pk2 = 1.159455691e-12
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.188354326e+00 ldsub = -1.491065479e-07 wdsub = -9.997544889e-07 pdsub = 2.381115266e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.821267712e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.346632754e-08 wvoff = -2.914402935e-07 pvoff = 6.941233471e-14
+ nfactor = {-1.076892670e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.096006075e-06 wnfactor = 2.075861869e-05 pnfactor = -4.944080214e-12
+ eta0 = 0.49
+ etab = -0.000625
+ u0 = 3.479454663e-02 lu0 = -7.280201048e-09 wu0 = -4.881350807e-08 pu0 = 1.162591322e-14
+ ua = 1.005800726e-08 lua = -2.861529868e-15 wua = -1.918646345e-14 pua = 4.569640000e-21
+ ub = -7.860689477e-18 lub = 2.288583175e-24 wub = 1.534487475e-23 pub = -3.654688820e-30
+ uc = -3.037746542e-10 luc = 7.036735037e-17 wuc = 4.718107649e-16 puc = -1.123711699e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.421504712e+05 lvsat = 8.706196536e-02 wvsat = 5.837476082e-01 pvsat = -1.390311679e-7
+ a0 = 1.227525634e+00 la0 = -1.118031034e-07 wa0 = -7.496361233e-07 pa0 = 1.785408355e-13
+ ags = 2.794660464e+01 lags = -6.358330333e-06 wags = -4.263239531e-05 pags = 1.015375759e-11
+ a1 = 0.0
+ a2 = 4.279179867e+00 la2 = -8.612954564e-07 wa2 = -5.774957647e-06 pa2 = 1.375421663e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = 7.924760166e-02 lketa = -3.627319612e-08 wketa = -2.432105844e-07 pketa = 5.792546489e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.799801776e+00 lpclm = 6.036400064e-07 wpclm = 4.047386347e-06 ppclm = -9.639660063e-13
+ pdiblc1 = -1.760065431e+00 lpdiblc1 = 5.291189255e-07 wpdiblc1 = 3.547724956e-06 ppdiblc1 = -8.449616527e-13
+ pdiblc2 = -3.925237439e-02 lpdiblc2 = 1.170171831e-08 wpdiblc2 = 7.845963560e-08 ppdiblc2 = -1.868673141e-14
+ pdiblcb = 5.039710497e+00 lpdiblcb = -1.253804720e-06 wpdiblcb = -8.406719321e-06 ppdiblcb = 2.002228341e-12
+ drout = -5.803435209e+00 ldrout = 1.545210928e-06 wdrout = 1.036058834e-05 pdrout = -2.467581325e-12
+ pscbe1 = 7.961143031e+08 lpscbe1 = 9.254565495e-01 wpscbe1 = 6.205155662e+00 ppscbe1 = -1.477881924e-6
+ pscbe2 = 4.595005894e-09 lpscbe2 = 1.125347475e-15 wpscbe2 = 7.545417730e-15 ppscbe2 = -1.797092141e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 2.893550342e+00 lbeta0 = 1.441605934e-06 wbeta0 = 9.665920273e-06 pbeta0 = -2.302132231e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -5.495845138e-09 lagidl = 1.385290837e-15 wagidl = 9.288329406e-15 pagidl = -2.212201415e-21
+ bgidl = 2.050991832e+09 lbgidl = -2.503147305e+02 wbgidl = -1.678352018e+03 pbgidl = 3.997331001e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.00081386752815302
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207367379934e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 1.945619966e-01 lkt1 = -1.692059687e-07 wkt1 = -1.134520443e-06 pkt1 = 2.702087339e-13
+ kt2 = -7.812934684e-02 lkt2 = 6.987276018e-09 wkt2 = 4.684945540e-08 pkt2 = -1.115813479e-14
+ at = 9.065936015e+05 lat = -2.135725658e-01 wat = -1.431997015e+00 pat = 3.410587289e-7
+ ute = 5.074444902e-01 lute = -1.256214540e-07 wute = -8.422877088e-07 pute = 2.006076636e-13
+ ua1 = 2.529810302e-08 lua1 = -5.821999668e-15 wua1 = -3.903631588e-14 pua1 = 9.297279353e-21
+ ub1 = -2.617699729e-17 lub1 = 6.122837978e-24 wub1 = 4.105342684e-23 pub1 = -9.777694670e-30
+ uc1 = -2.429053045e-09 luc1 = 5.722729824e-16 wuc1 = 3.837071485e-15 puc1 = -9.138753156e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.44 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -3.7585e-8
+ vth0 = {-1.104829786e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.393298119e-08 wvth0 = 9.851052022e-08 pvth0 = -2.513692944e-14
+ k1 = 1.509024879e-01 lk1 = 2.068218601e-07 wk1 = -2.325460876e-07 pk1 = 5.933878518e-14
+ k2 = 1.660529626e-01 lk2 = -8.512619440e-08 wk2 = 1.975827347e-08 pk2 = -5.041718641e-15
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.744671206e+00 ldsub = -5.568747918e-07 wdsub = -2.916530423e-07 pdsub = 7.442110681e-14
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-4.877784046e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.132123641e-08 wvoff = -4.760931314e-07 pvoff = 1.214846843e-13
+ nfactor = {6.916152080e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.195710033e-06 wnfactor = -1.404425904e-06 pnfactor = 3.583673579e-13
+ eta0 = -2.106274900e-02 leta0 = 1.304078817e-07 weta0 = 4.864635952e-06 peta0 = -1.241309156e-12
+ etab = -1.686473160e+00 letab = 4.301778749e-07 wetab = 3.229027898e-06 petab = -8.239510488e-13
+ u0 = 2.355796531e-02 lu0 = -4.932605777e-09 wu0 = -2.952006025e-08 pu0 = 7.532633773e-15
+ ua = 9.801920811e-09 lua = -3.000433387e-15 wua = -2.016809958e-14 pua = 5.146293970e-21
+ ub = -1.130914586e-17 lub = 3.331879335e-24 wub = 2.362673574e-23 pub = -6.028834159e-30
+ uc = -7.305766055e-11 luc = 1.651794680e-17 wuc = 1.454110036e-16 puc = -3.710452580e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.754943121e+05 lvsat = -1.408791809e-01 wvsat = -1.823024689e-01 pvsat = 4.651812099e-8
+ a0 = -9.557950160e+00 la0 = 2.632346519e-06 wa0 = 1.772825860e-05 pa0 = -4.523719747e-12
+ ags = 1.249999768e+00 lags = 5.224698008e-14
+ a1 = 0.0
+ a2 = -2.410682015e+00 la2 = 7.842794083e-07 wa2 = 4.479182916e-06 pa2 = -1.142953105e-12
+ b0 = 7.893132003e-23 lb0 = -2.014090493e-29 wb0 = -1.513051839e-28 pb0 = 3.860854377e-35
+ b1 = 0.0
+ keta = -8.078682022e-01 lketa = 1.875030503e-07 wketa = 5.105723943e-07 pketa = -1.302827579e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.952226074e+00 lpclm = -5.658485727e-07 wpclm = -2.724994975e-06 ppclm = 6.953369678e-13
+ pdiblc1 = 2.940665188e+00 lpdiblc1 = -6.325992741e-07 wpdiblc1 = -4.175887331e-07 ppdiblc1 = 1.065561170e-13
+ pdiblc2 = 7.670937173e-02 lpdiblc2 = -1.705300002e-08 wpdiblc2 = -3.636155387e-08 ppdiblc2 = 9.278377701e-15
+ pdiblcb = 4.649456788e+01 lpdiblcb = -1.192133423e-05 wpdiblcb = -7.640018903e-05 ppdiblcb = 1.949503623e-11
+ drout = -1.684270945e+00 ldrout = 6.044172108e-07 wdrout = -4.148540071e-12 pdrout = 1.058582971e-18
+ pscbe1 = 7.860086385e+08 lpscbe1 = 3.570175834e+00 wpscbe1 = 2.682035703e+01 ppscbe1 = -6.843750505e-6
+ pscbe2 = -4.803328210e-08 lpscbe2 = 1.463483231e-14 wpscbe2 = 1.102277613e-13 ppscbe2 = -2.812681786e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 2.382792894e+01 lbeta0 = -3.797321099e-06 wbeta0 = -1.547800002e-05 pbeta0 = 3.949521266e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.195082110e-08 lagidl = -5.519396268e-15 wagidl = -3.873652105e-14 pagidl = 9.884398077e-21
+ bgidl = 9.999997907e+08 lbgidl = 4.712768364e-5
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -2.8385e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.717392102e-01 lkt1 = 1.425359646e-08 wkt1 = 4.308028779e-07 pkt1 = -1.099279704e-13
+ kt2 = -1.614973469e-02 lkt2 = -8.329326711e-09 wkt2 = -1.863225081e-13 pkt2 = 4.754391436e-20
+ at = 2.325308195e+05 lat = -5.681626023e-02 wat = -5.880463428e-01 pat = 1.500517853e-7
+ ute = 1.923966989e+00 lute = -4.960420565e-07 wute = 1.092911242e-12 pute = -2.788781609e-19
+ ua1 = 6.368792505e-09 lua1 = -1.407367795e-15 wua1 = -4.308031979e-15 pua1 = 1.099280520e-21
+ ub1 = -2.926506882e-18 lub1 = 6.270437430e-25 wub1 = 1.906941532e-30 pub1 = -4.865942709e-37
+ uc1 = -1.008137180e-09 luc1 = 2.505453461e-16 wuc1 = 1.881172979e-15 puc1 = -4.800189092e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.45 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.094380677e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.070881130e-07 wvth0 = -1.421085472e-20
+ k1 = 4.212158315e-01 lk1 = 1.297050901e-6
+ k2 = 4.707115360e-02 lk2 = -5.440573537e-7
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.649382158e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.017359110e-8
+ nfactor = {1.316661266e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 9.663551657e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 9.516495432e-03 lu0 = -2.177360149e-8
+ ua = -5.607584256e-11 lua = -4.608090712e-15
+ ub = 8.723257589e-20 lub = 3.089023251e-24 wub = -1.540743956e-39
+ uc = -7.212392024e-11 luc = -7.437262497e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 160312.5
+ a0 = 1.723675260e+00 la0 = -1.853103320e-6
+ ags = 4.567962936e-01 lags = -6.490309596e-8
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.481931420e-02 lketa = 4.730386269e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.043721062e-01 lpclm = -2.892908447e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 1.361491196e-04 lpdiblc2 = 3.025582995e-9
+ pdiblcb = -3.450134580e-03 lpdiblcb = 3.850791507e-8
+ drout = 0.56
+ pscbe1 = 7.008119360e+08 lpscbe1 = 1.794156450e+3
+ pscbe2 = 9.666191697e-09 lpscbe2 = -6.130903958e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 5.684566553e-10 lalpha0 = -9.396383230e-15
+ alpha1 = -2.472842568e-11 lalpha1 = 2.501823966e-15 walpha1 = -1.033975766e-31 palpha1 = 1.292469707e-35
+ beta0 = 3.268634049e+00 lbeta0 = -5.388307414e-06 wbeta0 = 5.684341886e-20
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 8.848364432e-11 lagidl = 1.152305475e-15
+ bgidl = 1.563339129e+09 lbgidl = -1.129955201e+4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.257101581e-01 lkt1 = -5.983320405e-07 wkt1 = -7.105427358e-21
+ kt2 = -0.037961
+ at = 0.0
+ ute = -3.560052987e-01 lute = 5.278367351e-7
+ ua1 = 2.139515952e-09 lua1 = 7.212597973e-15
+ ub1 = -7.299472105e-19 lub1 = -1.907236690e-23
+ uc1 = 4.311997794e-11 luc1 = 7.677465592e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.46 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.0840563+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.4858803
+ k2 = 0.019947176
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.16743962+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.3648389+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0084309726
+ ua = -2.8581219e-10
+ ub = 2.4123582e-19
+ uc = -1.0920239e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 160312.5
+ a0 = 1.6312888
+ ags = 0.45356055
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.031235975
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.060146165
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00028698955
+ pdiblcb = -0.0015303226
+ drout = 0.56
+ pscbe1 = 790259600.0
+ pscbe2 = 9.3605355e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.4593183e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.45554
+ kt2 = -0.037961
+ at = 0.0
+ ute = -0.32969
+ ua1 = 2.4991e-9
+ ub1 = -1.6808e-18
+ uc1 = 4.2588e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.47 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.099435851e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.239310382e-7
+ k1 = 4.517138262e-01 lk1 = 2.753192546e-7
+ k2 = 2.896633464e-02 lk2 = -7.267791362e-08 wk2 = -4.440892099e-22
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.863612130e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.524734131e-7
+ nfactor = {6.023470053e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.144289311e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.071769316e-02 lu0 = -1.842678302e-8
+ ua = 3.672019860e-10 lua = -5.262099242e-15 pua = 2.646977960e-35
+ ub = -1.759105254e-19 lub = 3.361436166e-24
+ uc = -1.429063055e-10 luc = 2.715918809e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.223167722e+05 lvsat = -4.996409658e-1
+ a0 = 1.662786286e+00 la0 = -2.538121004e-7
+ ags = 4.597325700e-01 lags = -4.973518661e-8
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.754336036e-02 lketa = 5.082598348e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.208481702e-01 lpclm = 4.681751122e-06 wpclm = 1.776356839e-21 ppclm = -7.105427358e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 3.600260080e-04 lpdiblc2 = -5.885401950e-10
+ pdiblcb = -4.271034041e-04 lpdiblcb = -8.889927828e-9
+ drout = 0.56
+ pscbe1 = 7.803775502e+08 lpscbe1 = 7.963123697e+1
+ pscbe2 = 9.149402307e-09 lpscbe2 = 1.701347163e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -7.459246606e-01 lbeta0 = 3.018529772e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.925316236e-10 lagidl = -3.755090591e-16 wagidl = 3.308722450e-30
+ bgidl = 7.988221066e+08 lbgidl = 1.621125665e+3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.110862019e-01 lkt1 = 4.476007376e-7
+ kt2 = -3.127516492e-02 lkt2 = -5.387559563e-8
+ at = -1.820190699e+05 lat = 1.466740609e+0
+ ute = 1.702663986e-01 lute = -4.028733652e-6
+ ua1 = 5.377245473e-09 lua1 = -2.319258550e-14 pua1 = 2.117582368e-34
+ ub1 = -4.268705154e-18 lub1 = 2.085377968e-23 wub1 = -4.930380658e-38
+ uc1 = 7.964315027e-10 luc1 = -2.985967003e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.48 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.039182268e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.205882467e-7
+ k1 = 6.004806109e-01 lk1 = -3.284016481e-7
+ k2 = -6.050885308e-03 lk2 = 6.942791788e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.208171143e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.135156818e-7
+ nfactor = {2.996480249e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.571510395e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 4.093373681e-03 lu0 = 8.455831565e-9
+ ua = -1.478847421e-09 lua = 2.229483078e-15
+ ub = 1.027860336e-18 lub = -1.523670633e-24
+ uc = -6.663496362e-11 luc = -3.793019065e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.462869005e+05 lvsat = -1.910988216e-1
+ a0 = 2.032959356e+00 la0 = -1.756037345e-6
+ ags = 5.622897495e-01 lags = -4.659296555e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -4.174605632e-02 lketa = 6.788123813e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.441032208e-01 lpclm = -1.263270664e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 0.000215
+ pdiblcb = 2.041553198e-02 lpdiblcb = -9.347288545e-08 wpdiblcb = 1.110223025e-22 ppdiblcb = -2.220446049e-28
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.696808226e-08 lpscbe2 = -3.002818526e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.526703342e+00 lbeta0 = 4.729906941e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.141087571e+09 lbgidl = 2.321542270e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.414871760e-01 lkt1 = -2.406609414e-7
+ kt2 = -4.002107588e-02 lkt2 = -1.838320215e-8
+ at = 2.779140841e+05 lat = -3.997463191e-1
+ ute = -1.668881831e+00 lute = 3.434842518e-6
+ ua1 = -3.376869106e-09 lua1 = 1.233309966e-14 wua1 = 1.323488980e-29 pua1 = -1.323488980e-35
+ ub1 = 3.250298115e-18 lub1 = -9.659613820e-24 pub1 = 4.930380658e-44
+ uc1 = 9.326290009e-11 luc1 = -1.323892745e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.49 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.103865560e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.254096557e-8
+ k1 = 4.316923847e-01 lk1 = 1.899321537e-8
+ k2 = 3.069529095e-02 lk2 = -6.201959716e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 3.798690224e-01 ldsub = 3.707401741e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.831729372e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.482320221e-8
+ nfactor = {8.628159584e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.199334386e-7
+ eta0 = -6.708088940e-02 leta0 = 3.027174741e-7
+ etab = 7.371527644e-01 letab = -1.661257605e-06 wetab = -1.776356839e-21 petab = 3.552713679e-27
+ u0 = 8.743169528e-03 lu0 = -1.114238755e-9
+ ua = -3.520491852e-11 lua = -7.417786107e-16
+ ub = -1.078331476e-19 lub = 8.137796256e-25 pub = -6.162975822e-45
+ uc = -1.239932619e-10 luc = 8.012293822e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.946698149e+04 lvsat = 2.875473117e-2
+ a0 = 1.158873009e+00 la0 = 4.298095092e-8
+ ags = 7.823807504e-02 lags = 5.303309793e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.199495869e-03 lketa = -1.351230619e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.081281139e-02 lpclm = 6.370179576e-7
+ pdiblc1 = 4.101224041e-01 lpdiblc1 = -4.141532844e-8
+ pdiblc2 = -1.250655000e-05 lpdiblc2 = 4.682471560e-10
+ pdiblcb = -0.025
+ drout = 1.045812717e-01 ldrout = 9.373291640e-7
+ pscbe1 = 800000000.0
+ pscbe2 = -4.932972695e-09 lpscbe2 = 1.504790901e-14 ppscbe2 = -5.293955920e-35
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.722141263e+00 lbeta0 = 2.269492475e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.270154104e+09 lbgidl = -3.348664091e+1
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.434825322e-01 lkt1 = -3.073715895e-8
+ kt2 = -6.120850883e-02 lkt2 = 2.522413672e-8
+ at = 6.361637926e+04 lat = 4.131478816e-2
+ ute = 0.0
+ ua1 = 2.838982471e-09 lua1 = -4.601795842e-16
+ ub1 = -1.532952888e-18 lub1 = 1.851298980e-25
+ uc1 = 1.615321807e-10 luc1 = -2.728990597e-16 puc1 = -1.654361225e-36
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.50 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.132799035e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.315750087e-8
+ k1 = 3.162982928e-01 lk1 = 1.410997816e-7
+ k2 = 7.189253146e-02 lk2 = -4.979564370e-08 pk2 = -4.440892099e-28
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 4.290723551e-01 ldsub = 3.186746836e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.749039384e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 6.073195684e-9
+ nfactor = {2.038727531e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.243809106e-7
+ eta0 = 3.779934975e-01 leta0 = -1.682468899e-7
+ etab = -1.761891394e+00 letab = 9.831559518e-7
+ u0 = 1.053582632e-02 lu0 = -3.011174388e-9
+ ua = -2.505305958e-10 lua = -5.139274387e-16
+ ub = 5.707773262e-19 lub = 9.569438051e-26
+ uc = -6.648316323e-11 luc = 1.926747706e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.079322663e+04 lvsat = -4.393761653e-3
+ a0 = 1.220691836e+00 la0 = -2.243387722e-8
+ ags = -1.724220597e-01 lags = 7.955720141e-7
+ a1 = 0.0
+ a2 = 5.767431634e-01 la2 = 2.362436868e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.074606562e-02 lketa = -3.779261099e-08 pketa = 2.220446049e-28
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.258437974e-01 lpclm = 1.026093191e-7
+ pdiblc1 = -3.312122082e-01 lpdiblc1 = 7.430427182e-7
+ pdiblc2 = -2.259141628e-04 lpdiblc2 = 6.940686897e-10
+ pdiblcb = -5.253590337e-02 lpdiblcb = 2.913766687e-8
+ drout = 1.011770015e+00 ldrout = -2.263074892e-8
+ pscbe1 = 8.097631524e+08 lpscbe1 = -1.033107499e+1
+ pscbe2 = 9.343734185e-09 lpscbe2 = -5.927390603e-17
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.403618953e+00 lbeta0 = 4.902032285e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.0e-10
+ bgidl = 1.286351953e+09 lbgidl = -5.062671849e+1
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.514423374e-01 lkt1 = -2.231433193e-8
+ kt2 = -2.595084180e-02 lkt2 = -1.208446880e-8
+ at = 1.781915644e+05 lat = -7.992523550e-2
+ ute = 2.232680000e-02 lute = -2.362554996e-8
+ ua1 = 2.686310752e-09 lua1 = -2.986269514e-16
+ ub1 = -1.005683096e-18 lub1 = -3.728111783e-25
+ uc1 = -1.255383132e-10 luc1 = 3.087032485e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.51 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.061953872e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.613856140e-9
+ k1 = 8.545861681e-02 lk1 = 2.699475635e-7
+ k2 = 1.678694856e-01 lk2 = -1.033671002e-7
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.539539839e+00 ldsub = -3.011549518e-07 wdsub = -2.842170943e-20
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.064688737e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -3.212520435e-8
+ nfactor = {1.051585494e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.548792881e-7
+ eta0 = -4.330622374e-01 leta0 = 2.844600897e-07 weta0 = -1.776356839e-21 peta0 = -1.776356839e-27
+ etab = -3.454449539e-04 letab = -8.615047856e-11
+ u0 = 6.267522554e-03 lu0 = -6.287352768e-10
+ ua = -2.031465263e-10 lua = -5.403758048e-16
+ ub = -4.980063377e-19 lub = 6.922573582e-25 pub = -6.162975822e-45
+ uc = -6.110420944e-11 luc = 1.626510642e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.162297653e+04 lvsat = 4.160849047e-2
+ a0 = 1.701184033e+00 la0 = -2.906302066e-7
+ ags = 1.256474806e+00 lags = -1.995349257e-9
+ a1 = 0.0
+ a2 = 1.415545571e+00 la2 = -2.319506531e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.480137885e-02 lketa = -1.795109391e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.788400188e-01 lpclm = 1.721141822e-8
+ pdiblc1 = 1.663753220e+00 lpdiblc1 = -3.704871349e-07 wpdiblc1 = 2.842170943e-20
+ pdiblc2 = -9.906276727e-03 lpdiblc2 = 6.097356662e-09 wpdiblc2 = -2.775557562e-23 ppdiblc2 = 4.857225733e-29
+ pdiblcb = 2.761348617e-01 lpdiblcb = -1.543164941e-07 wpdiblcb = -4.787836794e-22 ppdiblcb = -1.734723476e-29
+ drout = 1.324772845e+00 ldrout = -1.973395382e-7
+ pscbe1 = 7.804736945e+08 lpscbe1 = 6.017421714e+0
+ pscbe2 = 9.135917840e-09 lpscbe2 = 5.672294325e-17
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.695363093e+00 lbeta0 = -2.308095986e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.718676123e-10 lagidl = 1.517483452e-16 pagidl = -8.271806126e-37
+ bgidl = 1.436825435e+09 lbgidl = -1.346165020e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.00081386752815302
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207367379934e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.612686559e-01 lkt1 = -1.682957573e-8
+ kt2 = -4.613287874e-02 lkt2 = -8.194612417e-10
+ at = 6.597676011e+04 lat = -1.729029819e-2
+ ute = -2.000000103e-02 lute = 5.744525966e-16
+ ua1 = 3.751219957e-09 lua1 = -8.930273222e-16
+ ub1 = -3.158301365e-18 lub1 = 8.287157609e-25
+ uc1 = -1.244341778e-10 luc1 = 3.025402956e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.52 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.05022704562893+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.961428255393082
+ k2 = -0.167552846831761
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.562303405039308
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.210713947389937+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.2302170822327+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.49
+ etab = -0.000625
+ u0 = 0.0042273003490566
+ ua = -1.95664558459119e-9
+ ub = 1.74834261966667e-18
+ uc = -8.324553995283e-12
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 123395.002071882
+ a0 = 0.758099999261006
+ ags = 1.24999997272013
+ a1 = 0.0
+ a2 = 0.662874470440252
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.0730519999606918
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.734690420259434
+ pdiblc1 = 0.461536473183962
+ pdiblc2 = 0.00987941513820755
+ pdiblcb = -0.224616327814465
+ drout = 0.684413503600629
+ pscbe1 = 800000000.518868
+ pscbe2 = 9.31998164677673e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.94639467130503
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 3.20550031084906e-10
+ bgidl = 999999975.393082
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.00081386752815302
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207367379934e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.515879992940252
+ kt2 = -0.0487919994941038
+ at = 9870.39612421382
+ ute = -0.0199999991650943
+ ua1 = 8.53380055896226e-10
+ ub1 = -4.69150049528303e-19
+ uc1 = -2.62609955581761e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.53 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.65e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -3.7585e-8
+ vth0 = {-1.043132251e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.810378780e-09 wvth0 = -1.563052137e-11 pvth0 = 3.988440142e-18
+ k1 = 5.284632489e-03 lk1 = 2.439791683e-07 wk1 = -5.730661996e-12 pk1 = 1.462293028e-18
+ k2 = 1.784277218e-01 lk2 = -8.828386171e-08 wk2 = -3.251757761e-12 pk2 = 8.297510306e-19
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.562013534e+00 ldsub = -5.102660337e-07 wdsub = 3.701273437e-11 pdsub = -9.444539430e-18
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-3.469089678e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.475288335e-08 wvoff = -9.752647259e-13 pvoff = 2.488582993e-19
+ nfactor = {6.036669578e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -9.712924834e-07 wnfactor = 3.905132462e-11 pnfactor = -9.964726473e-18
+ eta0 = 3.025184562e+00 leta0 = -6.469030446e-07 weta0 = 1.660446952e-11 peta0 = -4.236962482e-18
+ etab = 3.355614817e-01 letab = -8.578470453e-08 wetab = -3.705085124e-12 petab = 9.454265712e-19
+ u0 = 5.072378819e-03 lu0 = -2.156386731e-10 wu0 = -2.050421521e-14 pu0 = 5.232060674e-21
+ ua = -2.827442228e-09 lua = 2.222011795e-16 wua = 8.103105750e-21 pua = -2.067669469e-27
+ ub = 3.486046144e-18 lub = -4.434098082e-25 wub = -3.186039670e-29 pub = 8.129817424e-36
+ uc = 1.799934937e-11 luc = -6.717070422e-18 wuc = 6.124976884e-23 puc = -1.562910329e-29
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.613323153e+05 lvsat = -1.117484642e-01 wvsat = 5.335359782e-06 pvsat = -1.361423753e-12
+ a0 = 1.543564847e+00 la0 = -2.004270651e-07 wa0 = 5.052448728e-12 pa0 = -1.289233339e-18
+ ags = 1.249999768e+00 lags = 5.224698896e-14
+ a1 = 0.0
+ a2 = 3.941906188e-01 la2 = 6.856005843e-08 wa2 = 2.010070102e-11 pa2 = -5.129095896e-18
+ b0 = -1.581659877e-23 lb0 = 4.035921509e-30 wb0 = -1.478669219e-34 pb0 = 3.773120241e-41
+ b1 = 0.0
+ keta = -4.881434186e-01 lketa = 1.059188773e-07 wketa = -3.146608186e-12 pketa = 8.029200114e-19
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.245823844e+00 lpclm = -1.304259157e-07 wpclm = -3.713497335e-12 ppclm = 9.475730991e-19
+ pdiblc1 = 2.679180663e+00 lpdiblc1 = -5.658762678e-07 wpdiblc1 = -1.834207040e-11 ppdiblc1 = 4.680346095e-18
+ pdiblc2 = 5.393945724e-02 lpdiblc2 = -1.124280094e-08 wpdiblc2 = 2.235090690e-13 ppdiblc2 = -5.703280914e-20
+ pdiblcb = -1.347587131e+00 lpdiblcb = 2.865484598e-07 wpdiblcb = 8.280548514e-13 ppdiblcb = -2.112947541e-19
+ drout = -1.684296194e+00 ldrout = 6.044236534e-07 wdrout = 3.617153584e-11 pdrout = -9.229890821e-18
+ pscbe1 = 8.028026777e+08 lpscbe1 = -7.151591360e-01 wpscbe1 = 1.586447754e-03 ppscbe1 = -4.048138580e-10
+ pscbe2 = 2.099176548e-08 lpscbe2 = -2.978289081e-15 wpscbe2 = 1.442918262e-19 ppscbe2 = -3.681894547e-26
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.413555115e+01 lbeta0 = -1.324117059e-06 wbeta0 = -2.870326716e-11 pbeta0 = 7.324212675e-18
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.306161918e-09 lagidl = 6.702580881e-16 wagidl = -1.122079977e-20 pagidl = 2.863211469e-27
+ bgidl = 9.999997907e+08 lbgidl = 4.712767029e-5
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -2.8385e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.00081386752815302
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207367379934e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.019677198e-01 lkt1 = -5.458399475e-08 wkt1 = -1.150076400e-12 pkt1 = 2.934649785e-19
+ kt2 = -1.615086867e-02 lkt2 = -8.329037351e-09 wkt2 = 1.624564582e-12 pkt2 = -4.145401444e-19
+ at = -1.357048845e+05 lat = 3.714644437e-02 wat = -2.645832148e-06 pat = 6.751369890e-13
+ ute = 1.923973641e+00 lute = -4.960437538e-07 wute = -9.529202440e-12 pute = 2.431566577e-18
+ ua1 = 3.671078700e-09 lua1 = -7.189921630e-16 wua1 = 6.545575743e-21 pua1 = -1.670234570e-27
+ ub1 = -2.926495276e-18 lub1 = 6.270407815e-25 wub1 = -1.662681395e-29 pub1 = 4.242664120e-36
+ uc1 = 1.698601538e-10 luc1 = -5.004423369e-17 wuc1 = 3.120320697e-21 puc1 = -7.962122327e-28
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.54 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.152338226e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.513704283e-06 wvth0 = 9.081495803e-08 pvth0 = -5.181209623e-12
+ k1 = 1.970483572e-01 lk1 = 8.115548820e-06 wk1 = 3.512529473e-07 pk1 = -1.068405440e-11
+ k2 = 1.286906531e-01 lk2 = -2.162487226e-06 wk2 = -1.278913895e-07 pk2 = 2.535953373e-12
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.769994509e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.760540277e-06 wvoff = 1.889901472e-08 pvoff = -2.837247396e-12
+ nfactor = {1.373005597e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.630239487e-05 wnfactor = -8.828717197e-08 pnfactor = 2.705878434e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.347566517e-02 lu0 = -1.558540694e-07 wu0 = -6.203710162e-09 pu0 = 2.100936349e-13
+ ua = 3.049974204e-10 lua = 1.472650480e-14 wua = -5.657736393e-16 pua = -3.029580307e-20
+ ub = 2.490599981e-19 lub = -5.028257986e-23 wub = -2.535709480e-25 pub = 8.362913910e-29
+ uc = 6.808688066e-11 luc = -5.821482037e-15 wuc = -2.196993886e-16 puc = 7.956447253e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.603106084e+05 lvsat = 1.892678981e-04 wvsat = 2.963956202e-06 pvsat = -2.965680335e-10
+ a0 = 1.660311410e+00 la0 = 2.679089722e-05 wa0 = 9.928621024e-08 pa0 = -4.488291462e-11
+ ags = 3.605413385e-01 lags = 1.034736446e-05 wags = 1.508240068e-07 pags = -1.631521111e-11
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.037688366e-01 lketa = -3.226490678e-07 wketa = 7.670008359e-08 pketa = 1.246780554e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 7.007552736e-01 lpclm = -1.774108786e-05 wpclm = -7.777937054e-07 ppclm = 2.326593898e-11
+ pdiblc1 = 0.39
+ pdiblc2 = -2.946037909e-04 lpdiblc2 = 9.710049716e-09 wpdiblc2 = 6.749562121e-10 ppdiblc2 = -1.047403796e-14
+ pdiblcb = -1.254540710e-01 lpdiblcb = 1.178251771e-05 wpdiblcb = 1.911706520e-07 ppdiblcb = -1.840194732e-11
+ drout = 0.56
+ pscbe1 = 4.382143701e+08 lpscbe1 = 6.474742486e+03 wpscbe1 = 4.114699032e+02 ppscbe1 = -7.334113233e-3
+ pscbe2 = 7.611185491e-09 lpscbe2 = 2.732807441e-13 wpscbe2 = 3.220034435e-15 ppscbe2 = -4.378162583e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.982141126e-09 lalpha0 = -3.775230668e-14 walpha0 = -2.215133299e-15 palpha0 = 4.443152028e-20
+ alpha1 = -4.011274724e-10 lalpha1 = 1.005170003e-14 walpha1 = 5.897879470e-16 palpha1 = -1.183006691e-20
+ beta0 = 6.559987913e+00 lbeta0 = -2.698615475e-04 wbeta0 = -5.157294780e-06 pbeta0 = 4.144089383e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.414777873e-10 lagidl = -1.801932659e-14 wagidl = -8.303768856e-17 pagidl = 3.004045206e-20
+ bgidl = 3.263355063e+09 lbgidl = -4.539876062e+04 wbgidl = -2.663792367e+03 pbgidl = 5.343080015e-2
+ cgidl = 300.0
+ egidl = 6.942959155e-01 legidl = -5.946416174e-05 wegidl = -9.312153444e-07 pegidl = 9.317570324e-11
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.245168791e-01 lkt1 = -3.522028970e-06 wkt1 = -1.585619751e-07 pkt1 = 4.581205040e-12
+ kt2 = -4.885458026e-02 lkt2 = 1.089991706e-06 wkt2 = 1.706939057e-08 pkt2 = -1.707931983e-12
+ at = 0.0
+ ute = -2.860411391e-01 lute = -1.282568576e-05 wute = -1.096283809e-07 pute = 2.092392817e-11
+ ua1 = 5.426145170e-10 lua1 = 8.018488909e-14 wua1 = 2.502219990e-15 pua1 = -1.143418883e-19
+ ub1 = 2.869569686e-18 lub1 = -1.496786575e-22 wub1 = -5.640162214e-24 pub1 = 2.046498700e-28
+ uc1 = -1.440816848e-09 luc1 = 6.375158351e-14 wuc1 = 2.325213259e-15 puc1 = -8.786376900e-20
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.55 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-9.771625102e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} wvth0 = -1.674942308e-7
+ k1 = 6.016490171e-01 wk1 = -1.814005498e-7
+ k2 = 2.087985953e-02 wk2 = -1.461442335e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-8.922772115e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} wvoff = -1.225519450e-7
+ nfactor = {5.602497546e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} wnfactor = 1.260728433e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 5.705561047e-03 wu0 = 4.270507322e-9
+ ua = 1.039187269e-09 wua = -2.076170803e-15
+ ub = -2.257777857e-18 wub = 3.915759509e-24
+ uc = -2.221430873e-10 wuc = 1.769692633e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.603200444e+05 wvsat = -1.182144214e-5
+ a0 = 2.995971504e+00 wa0 = -2.138351352e-6
+ ags = 8.764091601e-01 wags = -6.625707899e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.198545049e-01 wketa = 1.388583240e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.837266039e-01 wpclm = 3.821296067e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 1.894907061e-04 wpdiblc2 = 1.527730835e-10
+ pdiblcb = 4.619633111e-01 wpdiblcb = -7.262583715e-7
+ drout = 0.56
+ pscbe1 = 7.610126356e+08 wpscbe1 = 4.582771189e+1
+ pscbe2 = 2.123559610e-08 wpscbe2 = -1.860729370e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -6.893958657e+00 wbeta0 = 1.550306149e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -7.568756812e-10 wagidl = 1.414628951e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -2.270289674e+00 wegidl = 3.714059037e-6
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.001076219e-01 wkt1 = 6.983398731e-8
+ kt2 = 5.486952670e-03 wkt2 = -6.807955289e-8
+ at = 0.0
+ ute = -9.254656608e-01 wute = 9.335339899e-7
+ ua1 = 4.540231902e-09 wua1 = -3.198294481e-15
+ ub1 = -4.592659295e-18 wub1 = 4.562656391e-24
+ uc1 = 1.737518140e-09 wuc1 = -2.055234658e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.56 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.039464975e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.020438552e-07 wvth0 = -9.396968477e-08 pvth0 = -5.924732914e-13
+ k1 = 4.395544491e-01 lk1 = 1.306185585e-06 wk1 = 1.905279541e-08 pk1 = -1.615287133e-12
+ k2 = 6.397728488e-02 lk2 = -3.472863801e-07 wk2 = -5.485942816e-08 pk2 = 4.302900475e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.854203722e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 7.751367346e-07 wvoff = -1.474224216e-09 pvoff = -9.756648570e-13
+ nfactor = {-3.367904986e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.165373869e-05 wnfactor = 6.221075191e-06 pnfactor = -3.997131744e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.527022300e-02 lu0 = -7.707367197e-08 wu0 = -7.133459154e-09 pu0 = 9.189510054e-14
+ ua = 3.803384462e-09 lua = -2.227437089e-14 wua = -5.384229918e-15 pua = 2.665690272e-20
+ ub = -4.144462113e-18 lub = 1.520322247e-23 wub = 6.218410791e-24 pub = -1.855515548e-29
+ uc = -3.604146801e-10 luc = 1.114216001e-15 wuc = 3.408186574e-16 puc = -1.320326272e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.223464537e+04 lvsat = 6.292254197e-01 wvsat = 2.194977663e-01 pvsat = -1.768845574e-6
+ a0 = 2.762766210e+00 la0 = 1.879207907e-06 wa0 = -1.723582741e-06 pa0 = -3.342275976e-12
+ ags = 9.393669959e-01 lags = -5.073249439e-07 wags = -7.515497339e-07 pags = 7.170074576e-13
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.483424359e-01 lketa = 2.295605913e-07 wketa = 1.736135090e-07 pketa = -2.800631891e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -2.821641705e+00 lpclm = 2.125676833e-05 wpclm = 3.605164007e-06 ppclm = -2.597175911e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 5.708932858e-03 lpdiblc2 = -4.447660316e-08 wpdiblc2 = -8.381319818e-09 ppdiblc2 = 6.876917140e-14
+ pdiblcb = 7.533649678e-01 lpdiblcb = -2.348164088e-06 wpdiblcb = -1.181133380e-06 ppdiblcb = 3.665460146e-12
+ drout = 0.56
+ pscbe1 = -5.791620826e+08 lpscbe1 = 1.079935571e+04 wpscbe1 = 2.130292561e+03 ppscbe1 = -1.679697211e-2
+ pscbe2 = 8.899760198e-08 lpscbe2 = -5.460377629e-13 wpscbe2 = -1.251159007e-13 ppscbe2 = 8.582644619e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -1.327249603e+01 lbeta0 = 5.139933852e-05 wbeta0 = 1.962816027e-05 pbeta0 = -3.324074724e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.320978648e-09 lagidl = 4.545637605e-15 wagidl = 2.371552542e-15 pagidl = -7.711052973e-21
+ bgidl = 1.917177767e+08 lbgidl = 6.513275563e+03 wbgidl = 9.512851308e+02 pbgidl = -7.665617303e-3
+ cgidl = 300.0
+ egidl = -4.675049286e+00 legidl = 1.937796176e-05 wegidl = 7.482129778e-06 pegidl = -3.036375460e-11
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -8.287776298e-01 lkt1 = 2.648478797e-06 wkt1 = 4.977976877e-07 pkt1 = -3.448604251e-12
+ kt2 = 2.027837890e-02 lkt2 = -1.191918271e-07 wkt2 = -8.078038200e-08 pkt2 = 1.023454401e-13
+ at = -4.536901304e+05 lat = 3.655912198e+00 wat = 4.256873615e-01 pat = -3.430261126e-6
+ ute = 1.182020579e+00 lute = -1.698248239e-05 wute = -1.585339884e-06 pute = 2.029751389e-11
+ ua1 = 1.991586369e-08 lua1 = -1.238994548e-13 wua1 = -2.278088073e-14 pua1 = 1.577998091e-19
+ ub1 = -1.967699579e-17 lub1 = 1.215521478e-22 wub1 = 2.414358958e-23 pub1 = -1.577864884e-28
+ uc1 = 3.235088994e-09 luc1 = -1.206768052e-14 wuc1 = -3.821186073e-15 puc1 = 1.423033671e-20
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.57 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-8.063874734e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.438242710e-07 wvth0 = -3.647712847e-07 pvth0 = 5.064856376e-13
+ k1 = 1.076123634e+00 lk1 = -1.277120382e-06 wk1 = -7.452955163e-07 pk1 = 1.486568255e-12
+ k2 = -8.961907422e-02 lk2 = 2.760337565e-07 wk2 = 1.309448337e-07 pk2 = -3.237352339e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -3.676219425e-01 ldsub = 3.764447538e-06 wdsub = 1.453511229e-06 pdsub = -5.898595666e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {1.411620170e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.501901197e-07 wvoff = -4.105008645e-07 pvoff = 6.842347836e-13
+ nfactor = {9.562862265e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.082151305e-05 wnfactor = -1.028900844e-05 pnfactor = 2.702940866e-11
+ eta0 = -1.668888352e-01 leta0 = 1.001916864e-06 weta0 = 3.868555474e-07 peta0 = -1.569925577e-12
+ etab = 1.458375140e-01 letab = -8.759053242e-07 wetab = -3.382005491e-07 petab = 1.372475322e-12
+ u0 = -1.059830024e-02 lu0 = 2.790519297e-08 wu0 = 2.302070708e-08 pu0 = -3.047563227e-14
+ ua = -3.320259392e-09 lua = 6.634586884e-15 wua = 2.885348929e-15 pua = -6.902454066e-21
+ ub = 6.714065832e-19 lub = -4.340391398e-24 wub = 5.585352280e-25 pub = 4.413581735e-30
+ uc = -3.941968353e-11 luc = -1.884362642e-16 wuc = -4.264422111e-17 puc = 2.358312778e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.264815510e+05 lvsat = -7.677870454e-01 wvsat = -4.390431621e-01 pvsat = 9.036254650e-7
+ a0 = 4.972802579e+00 la0 = -7.089495388e-06 wa0 = -4.606505024e-06 pa0 = 8.357112745e-12
+ ags = 1.746389676e+00 lags = -3.782360175e-06 wags = -1.855392226e-06 pags = 5.196587942e-12
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.880666405e-01 lketa = 3.907681668e-07 wketa = 2.292729425e-07 pketa = -5.059386320e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.501843674e+00 lpclm = -1.252135033e-05 wpclm = -7.141623786e-06 ppclm = 1.764053271e-11
+ pdiblc1 = 0.39
+ pdiblc2 = -1.020795804e-02 lpdiblc2 = 2.011684598e-08 wpdiblc2 = 1.633196226e-08 ppdiblc2 = -3.152152853e-14
+ pdiblcb = 3.802866368e-01 lpdiblcb = -8.341487972e-07 wpdiblcb = -5.638899512e-07 ppdiblcb = 1.160581381e-12
+ drout = 0.56
+ pscbe1 = 3.377143385e+09 lpscbe1 = -5.256004451e+03 wpscbe1 = -4.038182667e+03 ppscbe1 = 8.235749006e-3
+ pscbe2 = -7.322712350e-08 lpscbe2 = 1.122977513e-13 wpscbe2 = 1.413288522e-13 ppscbe2 = -2.230136411e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -1.254159816e+01 lbeta0 = 4.843323070e-05 wbeta0 = 2.831161912e-05 pbeta0 = -6.847969947e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -4.163727948e-10 lagidl = 8.745932692e-16 wagidl = 8.091158923e-16 pagidl = -1.370419435e-21
+ bgidl = 1.566854406e+09 lbgidl = 9.327373477e+02 wbgidl = -6.671434214e+02 pbgidl = -1.097759105e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 8.171089057e-02 lkt1 = -1.046438401e-06 wkt1 = -6.631183608e-07 pkt1 = 1.262590429e-12
+ kt2 = 2.134028729e-02 lkt2 = -1.235012319e-07 wkt2 = -9.614846990e-08 pkt2 = 1.647117534e-13
+ at = 8.072877814e+05 lat = -1.461350534e+00 wat = -8.294872926e-01 pat = 1.663451000e-6
+ ute = -6.302887656e+00 lute = 1.339254766e-05 wute = 7.261125675e-06 pute = -1.560294725e-11
+ ua1 = -2.361064703e-08 lua1 = 5.273852520e-14 wua1 = 3.170475177e-14 pua1 = -6.331215021e-20
+ ub1 = 2.166707672e-17 lub1 = -4.622912693e-23 wub1 = -2.885765556e-23 pub1 = 5.730157462e-29
+ uc1 = 3.185848902e-10 luc1 = -2.320110656e-16 wuc1 = -3.530619833e-16 puc1 = 1.560995761e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.58 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.033639938e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 2.389993400e-08 wvth0 = -1.100380727e-07 pvth0 = -1.779861753e-14
+ k1 = 6.744292113e-01 lk1 = -4.503649728e-07 wk1 = -3.803496739e-07 pk1 = 7.354476710e-13
+ k2 = -4.927085626e-02 lk2 = 1.929902648e-07 wk2 = 1.253007153e-07 pk2 = -3.121186788e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.383759653e+00 ldsub = -1.898363520e-06 wdsub = -3.139940315e-06 pdsub = 3.555508498e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.511778049e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.149493150e-08 wvoff = -5.013387679e-08 pvoff = -5.746173939e-14
+ nfactor = {-3.029468112e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.095643564e-06 wnfactor = 6.098905540e-06 pnfactor = -6.699704262e-12
+ eta0 = 4.299043781e-01 leta0 = -2.263850235e-07 weta0 = -7.787371493e-07 peta0 = 8.290623437e-13
+ etab = 3.275041966e-01 letab = -1.249806240e-06 wetab = 6.418873531e-07 petab = -6.447121953e-13
+ u0 = 5.732841310e-03 lu0 = -5.707072640e-09 wu0 = 4.716949512e-09 pu0 = 7.196612457e-15
+ ua = 1.229162538e-10 lua = -4.520539346e-16 wua = -2.477635436e-16 pua = -4.539759690e-22
+ ub = -7.937043777e-19 lub = -1.324943972e-24 wub = 1.074706720e-24 pub = 3.351213056e-30
+ uc = -2.710302850e-10 luc = 2.882577274e-16 wuc = 2.303955462e-16 puc = -3.261309801e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.203899956e+04 lvsat = 1.553444962e-01 wvsat = 9.637507484e-02 pvsat = -1.983562878e-7
+ a0 = 2.922677786e-01 la0 = 2.543840923e-06 wa0 = 1.357902801e-06 pa0 = -3.918652509e-12
+ ags = -1.781520799e-01 lags = 1.786739316e-07 wags = 4.017433743e-07 pags = 5.510191644e-13
+ a1 = 0.0
+ a2 = 1.438626299e+00 la2 = -1.314401490e-06 wa2 = -1.000677598e-06 pa2 = 2.059564612e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.360304892e-02 lketa = -4.488403794e-08 wketa = -4.043057508e-08 pketa = 4.915705667e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.271379880e+00 lpclm = 1.419095191e-06 wpclm = 2.024765156e-06 ppclm = -1.225454023e-12
+ pdiblc1 = -6.499984342e-01 lpdiblc1 = 2.140493577e-06 wpdiblc1 = 1.661126664e-06 ppdiblc1 = -3.418881066e-12
+ pdiblc2 = -1.347880124e-03 lpdiblc2 = 1.881299411e-09 wpdiblc2 = 2.092426231e-09 ppdiblc2 = -2.214142665e-15
+ pdiblcb = -0.025
+ drout = 1.352900990e-01 ldrout = 8.741251769e-07 wdrout = -4.811833710e-08 pdrout = 9.903571788e-14
+ pscbe1 = 8.044538782e+08 lpscbe1 = 3.902791177e+01 wpscbe1 = -6.978879745e+00 ppscbe1 = -6.115369356e-5
+ pscbe2 = -4.859844029e-08 lpscbe2 = 6.160773434e-14 wpscbe2 = 6.842038181e-14 ppscbe2 = -7.295561463e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.410205480e+00 lbeta0 = 3.252687005e-06 wbeta0 = -4.211986959e-06 pbeta0 = -1.540589138e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.214854894e-09 lagidl = -2.482750623e-15 wagidl = -1.746890660e-15 pagidl = 3.890276571e-21
+ bgidl = 2.085411307e+09 lbgidl = -1.345409086e+02 wbgidl = -1.277444446e+03 pbgidl = 1.583441552e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.991137551e-01 lkt1 = -5.681954036e-08 wkt1 = -6.952241299e-08 pkt1 = 4.086905725e-14
+ kt2 = -7.576154122e-02 lkt2 = 7.635083850e-08 wkt2 = 2.280346661e-08 pkt2 = -8.011155380e-14
+ at = -3.904681587e+04 lat = 2.805499439e-01 wat = 1.608652190e-01 pat = -3.748628287e-7
+ ute = -2.926946054e+00 lute = 6.444285930e-06 wute = 4.586296165e-06 pute = -1.009769340e-11
+ ua1 = -7.451543229e-09 lua1 = 1.948034253e-14 wua1 = 1.612445111e-14 pua1 = -3.124524280e-20
+ ub1 = 6.996514733e-18 lub1 = -1.603461637e-23 wub1 = -1.336501047e-23 pub1 = 2.541507726e-29
+ uc1 = 1.047074008e-09 luc1 = -1.731365513e-15 wuc1 = -1.387574971e-15 puc1 = 2.285303171e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.59 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.040807964e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.148492416e-08 wvth0 = -1.441428335e-07 pvth0 = 1.829001725e-14
+ k1 = -2.874354355e-01 lk1 = 5.674513405e-07 wk1 = 9.460036609e-07 pk1 = -6.680596374e-13
+ k2 = 4.011450935e-01 lk2 = -2.836263807e-07 wk2 = -5.159130830e-07 pk2 = 3.663945261e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.352572396e+00 ldsub = 3.113480964e-06 wdsub = 4.358620356e-06 pdsub = -4.379243446e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-3.833596256e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.791092078e-08 wvoff = -2.139913658e-07 pvoff = 1.159273397e-13
+ nfactor = {-2.167251158e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.119283308e-06 wnfactor = 3.534118373e-06 pnfactor = -3.985723425e-12
+ eta0 = 1.764363245e+00 leta0 = -1.638469363e-06 weta0 = -2.172333258e-06 peta0 = 2.303723938e-12
+ etab = -1.806366128e+00 letab = 1.008191321e-06 wetab = 6.968843902e-08 petab = -3.922847039e-14
+ u0 = -1.070629995e-02 lu0 = 1.168833347e-08 wu0 = 3.328475497e-08 pu0 = -2.303298224e-14
+ ua = -1.429568124e-09 lua = 1.190738459e-15 wua = 1.847459842e-15 pua = -2.671078498e-21
+ ub = -3.326718301e-18 lub = 1.355415372e-24 wub = 6.107071643e-24 pub = -1.973884535e-30
+ uc = 4.613567420e-11 luc = -4.735777563e-17 wuc = -1.764649340e-16 puc = 1.043965742e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.515326182e+06 lvsat = -1.471449218e+00 wvsat = -2.263470467e+00 pvsat = 2.298761469e-6
+ a0 = 2.825207985e+00 la0 = -1.364404159e-07 wa0 = -2.514151653e-06 pa0 = 1.786393537e-13
+ ags = -1.428114513e+00 lags = 1.501346679e-06 wags = 1.967572130e-06 pags = -1.105893850e-12
+ a1 = 0.0
+ a2 = -7.338616289e-01 la2 = 9.844600606e-07 wa2 = 2.053615482e-06 pa2 = -1.172396697e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = 4.375105758e-02 lketa = -6.620405626e-08 wketa = -3.604702801e-08 pketa = 4.451851866e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -2.941691079e+00 lpclm = 3.186568392e-06 wpclm = 5.433356683e-06 ppclm = -4.832323319e-12
+ pdiblc1 = -1.542745999e+00 lpdiblc1 = 3.085172268e-06 wpdiblc1 = 1.898378950e-06 ppdiblc1 = -3.669934318e-12
+ pdiblc2 = -3.518687094e-03 lpdiblc2 = 4.178382222e-09 wpdiblc2 = 5.159518347e-09 ppdiblc2 = -5.459647529e-15
+ pdiblcb = -1.172019504e-01 lpdiblcb = 9.756533787e-08 wpdiblcb = 1.013266518e-07 ppdiblcb = -1.072208231e-13
+ drout = 1.047288964e+00 ldrout = -9.092466248e-08 wdrout = -5.565542258e-08 pdrout = 1.070112356e-13
+ pscbe1 = 9.267076372e+08 lpscbe1 = -9.033734841e+01 wpscbe1 = -1.832428860e+02 ppscbe1 = 1.253635900e-4
+ pscbe2 = 1.035765614e-08 lpscbe2 = -7.778382134e-16 wpscbe2 = -1.588736616e-15 ppscbe2 = 1.125934222e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.427244749e+01 lbeta0 = -1.892391623e-06 wbeta0 = -9.195996549e-06 pbeta0 = 3.733340290e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.194236717e-09 lagidl = 1.124647847e-15 wagidl = 3.594889985e-15 pagidl = -1.762235454e-21
+ bgidl = 2.150490193e+09 lbgidl = -2.034054333e+02 wbgidl = -1.354037219e+03 pbgidl = 2.393923294e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.668637701e-01 lkt1 = 1.206884929e-07 wkt1 = 1.808563821e-07 pkt1 = -2.240742724e-13
+ kt2 = 9.582029589e-02 lkt2 = -1.052119141e-07 wkt2 = -1.908058746e-07 pkt2 = 1.459234428e-13
+ at = 4.396982134e+05 lat = -2.260436837e-01 wat = -4.097605215e-01 pat = 2.289562111e-7
+ ute = 6.114980409e+00 lute = -3.123609395e-06 wute = -9.546712978e-06 pute = 4.857432886e-12
+ ua1 = 2.218784354e-08 lua1 = -1.188316736e-14 wua1 = -3.055738076e-14 pua1 = 1.815207123e-20
+ ub1 = -1.797107983e-17 lub1 = 1.038534317e-23 wub1 = 2.658345338e-23 pub1 = -1.685718873e-29
+ uc1 = -1.589797975e-09 luc1 = 1.058893313e-15 wuc1 = 2.294380678e-15 puc1 = -1.610831837e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.60 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.010792788e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.473135326e-08 wvth0 = -8.016542866e-08 pvth0 = -1.742025082e-14
+ k1 = -1.138314552e+00 lk1 = 1.042386537e-06 wk1 = 1.917557101e-06 pk1 = -1.210351621e-12
+ k2 = 5.474270088e-01 lk2 = -3.652765574e-07 wk2 = -5.947370334e-07 pk2 = 4.103916906e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 7.444758193e+00 ldsub = -2.355095051e-06 wdsub = -9.253016554e-06 pdsub = 3.218363928e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {1.840204349e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -9.958037361e-08 wvoff = -1.956629873e-07 pvoff = 1.056969887e-13
+ nfactor = {2.193941989e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.737212502e-07 wnfactor = -3.272960725e-06 pnfactor = -1.862160849e-13
+ eta0 = -3.218632121e+00 leta0 = 1.142889161e-06 weta0 = 4.364770733e-06 peta0 = -1.345091397e-12
+ etab = 2.799881494e-03 letab = -1.630870621e-09 wetab = -4.928481208e-09 petab = 2.420455975e-15
+ u0 = 2.288220491e-02 lu0 = -7.059762289e-09 wu0 = -2.603391130e-08 pu0 = 1.007691771e-14
+ ua = 9.373963249e-09 lua = -4.839468647e-15 wua = -1.500658400e-14 pua = 6.736343154e-21
+ ub = -1.052435032e-17 lub = 5.372917637e-24 wub = 1.571049897e-23 pub = -7.334229565e-30
+ uc = -4.501954977e-11 luc = 3.522335731e-18 wuc = -2.520340710e-17 puc = 1.996692773e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.891720496e+06 lvsat = 9.884320263e-01 wvsat = 4.512888165e+00 pvsat = -1.483598628e-6
+ a0 = 4.213742446e+00 la0 = -9.114786958e-07 wa0 = -3.936983054e-06 pa0 = 9.728211563e-13
+ ags = 2.308663515e+00 lags = -5.844107123e-07 wags = -1.648697636e-06 pags = 9.125994455e-13
+ a1 = 0.0
+ a2 = 1.992345751e+00 la2 = -5.372271129e-07 wa2 = -9.038008924e-07 pa2 = 4.783444010e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = 7.074518612e-02 lketa = -8.127136899e-08 wketa = -1.340447947e-07 pketa = 9.921793207e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.915265502e+00 lpclm = -1.198949062e-06 wpclm = -6.638148291e-06 ppclm = 1.905628612e-12
+ pdiblc1 = 8.131110992e+00 lpdiblc1 = -2.314484489e-06 wpdiblc1 = -1.013384517e-05 ppdiblc1 = 3.046092222e-12
+ pdiblc2 = -5.872621502e-03 lpdiblc2 = 5.492277791e-09 wpdiblc2 = -6.320423112e-09 ppdiblc2 = 9.481113950e-16
+ pdiblcb = 4.357062023e-01 lpdiblcb = -2.110514057e-07 wpdiblcb = -2.500358441e-07 ppdiblcb = 8.889918121e-14
+ drout = 4.042210614e-01 ldrout = 2.680165489e-07 wdrout = 1.442432841e-06 pdrout = -7.291766907e-13
+ pscbe1 = 7.214405196e+08 lpscbe1 = 2.423659862e+01 wpscbe1 = 9.250038050e+01 ppscbe1 = -2.854802912e-5
+ pscbe2 = 7.911284505e-09 lpscbe2 = 5.876530413e-16 wpscbe2 = 1.918904914e-15 ppscbe2 = -8.319260511e-22
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.330645925e+01 lbeta0 = -1.353205969e-06 wbeta0 = -5.658306017e-06 pbeta0 = 1.758707566e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.616000796e-09 lagidl = 8.018939029e-16 wagidl = 2.262844056e-15 pagidl = -1.018727378e-21
+ bgidl = 3.723602198e+09 lbgidl = -1.081469361e+03 wbgidl = -3.583200818e+03 pbgidl = 1.483644576e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.526319122e-01 lkt1 = -1.105233032e-07 wkt1 = -4.836097038e-07 pkt1 = 1.468107628e-13
+ kt2 = -1.623589917e-01 lkt2 = 3.889601885e-08 wkt2 = 1.821172533e-07 pkt2 = -6.223105950e-14
+ at = 2.966940766e+05 lat = -1.462230646e-01 wat = -3.615160389e-01 pat = 2.020275883e-7
+ ute = -1.957045185e+00 lute = 1.381953131e-06 wute = 3.035198714e-06 pute = -2.165412763e-12
+ ua1 = -1.140432391e-09 lua1 = 1.137976413e-15 wua1 = 7.664837681e-15 pua1 = -3.182424434e-21
+ ub1 = 3.094014055e-18 lub1 = -1.372560284e-24 wub1 = -9.796890583e-24 pub1 = 3.449227862e-30
+ uc1 = 4.305508245e-10 luc1 = -6.880477608e-17 wuc1 = -8.696182097e-16 puc1 = 1.552174218e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.61 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -3.7585e-8
+ vth0 = {-7.317914118e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.517887854e-08 wvth0 = -4.989638002e-07 pvth0 = 1.177994387e-13
+ k1 = 8.216894870e+00 lk1 = -1.942144327e-06 wk1 = -1.136875026e-05 pk1 = 3.043188674e-12
+ k2 = -2.781324024e+00 lk2 = 6.969831694e-07 wk2 = 4.095575560e-06 pk2 = -1.092118262e-12
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -5.212353646e+00 ldsub = 1.630700701e-06 wdsub = 9.048437176e-06 pdsub = -2.555180804e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-7.282093693e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.377019722e-07 wvoff = 8.108749615e-07 pvoff = -2.157682496e-13
+ nfactor = {-2.625609989e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.383576803e-06 wnfactor = 7.608702267e-06 pnfactor = -3.734878931e-12
+ eta0 = -3.106474351e+00 leta0 = 1.169465565e-06 weta0 = 5.635394784e-06 peta0 = -1.832461322e-12
+ etab = -2.957267567e-01 letab = 9.535107039e-08 wetab = 4.624014348e-07 petab = -1.494076899e-13
+ u0 = -2.992973102e-02 lu0 = 9.723647668e-09 wu0 = 5.352140391e-08 pu0 = -1.523619745e-14
+ ua = -2.482735616e-08 lua = 6.014808208e-15 wua = 3.583661956e-14 pua = -9.424735307e-21
+ ub = 2.668706958e-17 lub = -6.430726223e-24 wub = -3.907703992e-23 pub = 1.007644640e-29
+ uc = -2.147148160e-10 luc = 5.889645284e-17 wuc = 3.233974421e-16 puc = -9.228614768e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.982764665e+05 lvsat = -1.569180684e-01 wvsat = -1.057486614e+00 pvsat = 2.458783736e-7
+ a0 = 1.979645128e+00 la0 = -2.352984075e-07 wa0 = -1.914065937e-06 pa0 = 3.686942513e-13
+ ags = -2.641481580e+00 lags = 9.929893268e-07 wags = 6.097648058e-06 pags = -1.555936822e-12
+ a1 = 0.0
+ a2 = -1.389548314e+00 la2 = 5.328275920e-07 wa2 = 3.215986414e-06 pa2 = -8.348992761e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.493612421e-01 lketa = 5.085135544e-08 wketa = 4.329550303e-07 pketa = -7.968010757e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.942708962e+00 lpclm = -2.985021066e-07 wpclm = -1.892870830e-06 ppclm = 4.677295179e-13
+ pdiblc1 = 3.525118905e-01 lpdiblc1 = 8.720553172e-08 wpdiblc1 = 1.708330172e-07 ppdiblc1 = -1.366442662e-13
+ pdiblc2 = -2.746552275e-03 lpdiblc2 = 4.778751835e-09 wpdiblc2 = 1.978390611e-08 ppdiblc2 = -7.487931383e-15
+ pdiblcb = -3.427918463e-01 lpdiblcb = 3.045028956e-08 wpdiblcb = 1.851718197e-07 ppdiblcb = -4.771322862e-14
+ drout = 2.839225247e+00 ldrout = -5.089888014e-07 wdrout = -3.376421926e-06 pdrout = 7.975457506e-13
+ pscbe1 = 8.004058320e+08 lpscbe1 = -1.035556232e-01 wpscbe1 = -6.359062991e-01 ppscbe1 = 1.622635843e-7
+ pscbe2 = 1.065821759e-08 lpscbe2 = -2.731496869e-16 wpscbe2 = -2.096911338e-15 ppscbe2 = 4.280042537e-22
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.169660883e+00 lbeta0 = 1.868328019e-06 wbeta0 = 9.051691261e-06 pbeta0 = -2.927524276e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.801304625e-08 lagidl = -5.536647362e-15 wagidl = -2.772276155e-14 pagidl = 8.675494557e-21
+ bgidl = -2.649916736e+09 lbgidl = 9.313492282e+02 wbgidl = 5.719134793e+03 pbgidl = -1.459351595e-3
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -2.8385e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -8.080083783e-01 lkt1 = 9.648851534e-08 wkt1 = 4.577423939e-07 pkt1 = -1.511899774e-13
+ kt2 = -3.787465448e-02 lkt2 = 5.631208133e-10 wkt2 = -1.710662809e-08 pkt2 = -8.823663910e-16
+ at = -6.485230269e+05 lat = 1.530668795e-01 wat = 1.031651139e+00 pat = -2.398438609e-7
+ ute = 8.963980259e+00 lute = -2.093002156e-06 wute = -1.407719631e-05 pute = 3.279571125e-12
+ ua1 = 4.094007903e-09 lua1 = -5.013308004e-16 wua1 = -5.077811068e-15 pua1 = 7.855462605e-22
+ ub1 = -1.005319057e-18 lub1 = -1.152965416e-25 wub1 = 8.401350134e-25 pub1 = 1.806606876e-31
+ uc1 = 7.711680226e-10 luc1 = -1.833588416e-16 wuc1 = -1.249509072e-15 puc1 = 2.873090028e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.62 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.26e-06 wmax = 1.65e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -3.7585e-8
+ vth0 = {-9.979491039e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.263420252e-09 wvth0 = -7.081409755e-08 pvth0 = 8.548479089e-15
+ k1 = -3.235842785e+00 lk1 = 9.802507399e-07 wk1 = 5.078588124e-06 pk1 = -1.153678661e-12
+ k2 = 1.340176991e+00 lk2 = -3.547002446e-07 wk2 = -1.820373740e-06 pk2 = 4.174545213e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 9.212718346e+00 ldsub = -2.050144919e-06 wdsub = -1.042109867e-05 pdsub = 2.412860659e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-7.357612698e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.396289906e-07 wvoff = 6.093002516e-07 pvoff = -1.643324309e-13
+ nfactor = {2.200899237e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.902434681e-06 wnfactor = -2.502734492e-05 pnfactor = 4.592861229e-12
+ eta0 = 1.166238683e+01 leta0 = -2.599104742e-06 weta0 = -1.353380564e-05 peta0 = 3.058943551e-12
+ etab = 1.428653197e+00 letab = -3.446589625e-07 wetab = -1.712793162e-06 petab = 4.056367154e-13
+ u0 = 1.157207661e-02 lu0 = -8.663685869e-10 wu0 = -1.018453997e-08 pu0 = 1.019648250e-15
+ ua = -4.754208825e-09 lua = 8.927432022e-16 wua = 3.019101073e-15 pua = -1.050689115e-21
+ ub = 8.466910935e-18 lub = -1.781488343e-24 wub = -7.804658481e-24 pub = 2.096672823e-30
+ uc = 1.218607767e-10 luc = -2.698754115e-17 wuc = -1.627426942e-16 puc = 3.176223090e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.942857221e+06 lvsat = -4.489807396e-01 wvsat = -2.164736434e+00 pvsat = 5.284153100e-7
+ a0 = 4.213334363e+00 la0 = -8.052688895e-07 wa0 = -4.183315538e-06 pa0 = 9.477386719e-13
+ ags = 1.249999068e+00 lags = 2.099152319e-13 wags = 1.097188147e-12 pags = -2.470538547e-19
+ a1 = 0.0
+ a2 = -3.808730910e-01 la2 = 2.754439353e-07 wa2 = 1.214484479e-06 pa2 = -3.241760272e-13
+ b0 = -6.354749858e-23 lb0 = 1.621541521e-29 wb0 = 7.479044913e-29 pb0 = -1.908427890e-35
+ b1 = 0.0
+ keta = -1.817818101e+00 lketa = 4.255574922e-07 wketa = 2.083493367e-06 pketa = -5.008479748e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.826488480e+00 lpclm = -5.240161260e-07 wpclm = -2.476781906e-06 ppclm = 6.167261071e-13
+ pdiblc1 = 9.604156600e+00 lpdiblc1 = -2.273536649e-06 wpdiblc1 = -1.085091549e-05 ppdiblc1 = 2.675775300e-12
+ pdiblc2 = 1.930039166e-01 lpdiblc2 = -4.517089532e-08 wpdiblc2 = -2.179029373e-07 ppdiblc2 = 5.316262046e-14
+ pdiblcb = -4.735270882e+00 lpdiblcb = 1.151279165e-06 wpdiblcb = 5.308237027e-06 ppdiblcb = -1.354965778e-12
+ drout = -8.672267067e+00 ldrout = 2.428398692e-06 wdrout = 1.094964147e-05 pdrout = -2.858035846e-12
+ pscbe1 = 8.112645225e+08 lpscbe1 = -2.874367686e+00 wpscbe1 = -1.325746440e+01 ppscbe1 = 3.382906566e-6
+ pscbe2 = 5.648242051e-08 lpscbe2 = -1.196611155e-14 wpscbe2 = -5.561094386e-14 ppscbe2 = 1.408317993e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.134020937e+01 lbeta0 = -5.319950837e-06 wbeta0 = -2.695838616e-05 pbeta0 = 6.261167180e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.423832843e-08 lagidl = 2.692935916e-15 wagidl = 1.869676300e-14 pagidl = -3.169375524e-21
+ bgidl = 9.999991591e+08 lbgidl = 1.893471966e-04 wbgidl = 9.896828232e-04 pbgidl = -2.228468800e-10
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -2.8385e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 4.295686792e-01 lkt1 = -2.193040224e-07 wkt1 = -1.146261627e-06 pkt1 = 2.581037287e-13
+ kt2 = 9.548021826e-02 lkt2 = -3.346504206e-08 wkt2 = -1.749155814e-07 pkt2 = 3.938574424e-14
+ at = -6.335523440e+05 lat = 1.492468103e-01 wat = 7.800854911e-01 pat = -1.756518545e-7
+ ute = 8.571970088e+00 lute = -1.992972921e-06 wute = -1.041690142e-05 pute = 2.345573676e-12
+ ua1 = 1.345013646e-08 lua1 = -2.888734124e-15 wua1 = -1.532301419e-14 pua1 = 3.399814742e-21
+ ub1 = -1.133019940e-17 lub1 = 2.519303175e-24 wub1 = 1.316793224e-23 pub1 = -2.965023331e-30
+ uc1 = 8.405662892e-10 luc1 = -2.010671973e-16 wuc1 = -1.050941079e-15 puc1 = 2.366404080e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.63 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 1.12e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-5.235572575e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.195307956e-05 wvth0 = -6.492111968e-07 pvth0 = 1.302198855e-11
+ k1 = 9.978156426e-01 lk1 = -1.103796988e-05 wk1 = -5.911876878e-07 pk1 = 1.185814314e-11
+ k2 = -2.249039941e-01 lk2 = 4.905067096e-06 wk2 = 2.882619299e-07 pk2 = -5.782006795e-12
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 9.962867658e-05 lcit = -1.797787232e-09 wcit = -1.054859613e-10 pcit = 2.115855344e-15
+ voff = {-1.626663355e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.155969615e-07 wvoff = 2.030055819e-09 pvoff = -4.071920473e-14
+ nfactor = {-6.217119814e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.519446452e-05 wnfactor = 2.259339830e-06 pnfactor = -4.531822240e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 9.694147868e-03 lu0 = -7.221901346e-09 wu0 = -1.753159258e-09 pu0 = 3.516516644e-14
+ ua = 4.043268237e-09 lua = -9.564034879e-14 wua = -4.965426806e-15 pua = 9.959737499e-20
+ ub = -3.601511520e-18 lub = 9.368875610e-23 wub = 4.278251384e-24 pub = -8.581389357e-29
+ uc = -1.513736216e-10 luc = 1.596564392e-15 wuc = 3.858850465e-17 puc = -7.740147864e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.028522955e+05 lvsat = -1.489403960e+01 wvsat = -8.739106835e-01 pvsat = 1.752904905e-5
+ a0 = 3.294371801e+00 la0 = -4.242908313e-05 wa0 = -1.823875413e-06 pa0 = 3.658360309e-11
+ ags = 3.640828848e+00 lags = -6.674133116e-05 wags = -3.709818529e-06 pags = 7.441217072e-11
+ a1 = 0.0
+ a2 = -7.748150016e-01 la2 = 3.158790702e-05 wa2 = 1.853434421e-06 pa2 = -3.717650271e-11
+ b0 = -5.306756011e-08 lb0 = 1.064438142e-12 wb0 = 6.245637898e-14 pb0 = -1.252760667e-18
+ b1 = -3.304702963e-07 lb1 = 6.628629383e-12 wb1 = 3.889377620e-13 pb1 = -7.801379750e-18
+ keta = -5.443666722e-01 lketa = 1.088148646e-05 wketa = 5.952493694e-07 pketa = -1.193961304e-11
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.581010114e-01 lpclm = -6.361288781e-06 wpclm = -4.922085659e-07 ppclm = 9.872803090e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -8.893660407e-03 lpdiblc2 = 1.847950863e-07 wpdiblc2 = 1.079537512e-08 ppdiblc2 = -2.165354694e-13
+ pdiblcb = 2.107116307e+00 lpdiblcb = -4.537631100e-05 wpdiblcb = -2.436390542e-06 ppdiblcb = 4.886953569e-11
+ drout = 0.56
+ pscbe1 = 6.975982990e+08 lpscbe1 = 2.053012890e+03 wpscbe1 = 1.061952508e+02 ppscbe1 = -2.130082394e-3
+ pscbe2 = 3.861803511e-09 lpscbe2 = 3.136414383e-14 wpscbe2 = 7.632764572e-15 ppscbe2 = -1.530992894e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.026361766e-09 lalpha0 = -1.858112178e-14 walpha0 = -1.090255542e-15 palpha0 = 2.186853100e-20
+ alpha1 = 1.026361766e-09 lalpha1 = -1.858112178e-14 walpha1 = -1.090255542e-15 palpha1 = 2.186853100e-20
+ beta0 = -2.479397080e+02 lbeta0 = 5.099153824e-03 wbeta0 = 2.943689963e-04 pbeta0 = -5.904503371e-9
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.618047850e-08 lagidl = 3.334786344e-13 wagidl = 1.912663175e-14 pagidl = -3.836452312e-19
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -9.693353258e-02 legidl = 1.970480888e-05 pegidl = -1.421085472e-26
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -6.194108128e-01 lkt1 = 3.583177705e-06 wkt1 = 1.885051832e-07 pkt1 = -3.781069011e-12
+ kt2 = 1.563404062e-01 lkt2 = -4.186117578e-06 wkt2 = -2.244291033e-07 pkt2 = 4.501637107e-12
+ at = -6.576242174e+05 lat = 1.319073835e+01 wat = 7.739724092e-01 pat = -1.552447016e-5
+ ute = -2.664616634e+00 lute = 5.079431711e-05 wute = 2.689769448e-06 pute = -5.395185284e-11
+ ua1 = 6.456578994e-09 lua1 = -9.294664522e-14 wua1 = -4.458054911e-15 pua1 = 8.942042327e-20
+ ub1 = -6.108958210e-18 lub1 = 1.081751014e-22 wub1 = 4.926864794e-24 pub1 = -9.882389161e-29
+ uc1 = 4.755999750e-09 luc1 = -9.557238659e-14 wuc1 = -4.967956525e-15 puc1 = 9.964811654e-20
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.64 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.12e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.119478+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.44751769
+ k2 = 0.01963811
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.19335692+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.6314579+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0093341
+ ua = -7.2488104e-10
+ ub = 1.06934111e-18
+ uc = -7.1776909e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 160310.0
+ a0 = 1.17907
+ ags = 0.31344
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.0018702
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.14095898
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00031929802
+ pdiblcb = -0.15511953
+ drout = 0.56
+ pscbe1 = 799951250.0
+ pscbe2 = 5.4254628e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.2785893
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 4.4509773e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.88544965
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.4407715
+ kt2 = -0.052358472
+ at = 0.0
+ ute = -0.13226612
+ ua1 = 1.8227243e-9
+ ub1 = -7.1588888e-19
+ uc1 = -8.7612717e-12
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.65 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.12e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.119308571e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.365284442e-9
+ k1 = 4.557431136e-01 lk1 = -6.628186177e-8
+ k2 = 1.736465621e-02 lk2 = 1.831987716e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.866729821e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.386030771e-8
+ nfactor = {1.917980732e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.308849687e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 9.209108364e-03 lu0 = 1.007203851e-9
+ ua = -7.714556020e-10 lua = 3.753057380e-16
+ ub = 1.139159733e-18 lub = -5.626103368e-25
+ uc = -7.082993503e-11 luc = -7.630877232e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.687361861e+05 lvsat = -8.737166397e-1
+ a0 = 1.298282802e+00 la0 = -9.606370240e-7
+ ags = 3.007947423e-01 lags = 1.018976364e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.275546727e-04 lketa = -8.401813297e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.415723457e-01 lpclm = -8.107596053e-07 wpclm = 4.440892099e-22
+ pdiblc1 = 0.39
+ pdiblc2 = -1.412456511e-03 lpdiblc2 = 1.395477241e-08 wpdiblc2 = 8.673617380e-25 ppdiblc2 = -3.469446952e-30
+ pdiblcb = -2.502133320e-01 lpdiblcb = 7.662820228e-7
+ drout = 0.56
+ pscbe1 = 1.230892076e+09 lpscbe1 = -3.472594437e+03 wpscbe1 = 1.907348633e-12
+ pscbe2 = -1.731012336e-08 lpscbe2 = 1.832072184e-13 ppscbe2 = 1.058791184e-34
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.405041024e+00 lbeta0 = 2.315554051e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.940678393e-10 lagidl = -2.006243465e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 1.682321702e+00 legidl = -6.421330460e-6
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.058118873e-01 lkt1 = -2.817105026e-7
+ kt2 = -4.835860979e-02 lkt2 = -3.223156969e-8
+ at = -9.199465573e+04 lat = 7.413085750e-1
+ ute = -1.650014701e-01 lute = 2.637870157e-7
+ ua1 = 5.595420866e-10 lua1 = 1.017893702e-14
+ ub1 = 8.371840607e-19 lub1 = -1.251492578e-23
+ uc1 = -1.167338578e-11 luc1 = 2.346631032e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.66 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.12e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.116324143e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.347660345e-8
+ k1 = 4.428654258e-01 lk1 = -1.402201541e-8
+ k2 = 2.164134381e-02 lk2 = 9.643518320e-10
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.673887289e-01 ldsub = -1.247435718e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.076298863e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.118637217e-8
+ nfactor = {8.205595117e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.144672185e-6
+ eta0 = 1.618122575e-01 leta0 = -3.320080490e-7
+ etab = -1.415226926e-01 letab = 2.902512456e-7
+ u0 = 8.961795573e-03 lu0 = 2.010841203e-9
+ ua = -8.686534836e-10 lua = 7.697512652e-16
+ ub = 1.145979433e-18 lub = -5.902858386e-25
+ uc = -7.565336861e-11 luc = 1.194343622e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 53438.0
+ a0 = 1.058775121e+00 la0 = 1.132585948e-8
+ ags = 1.699111794e-01 lags = 6.330453849e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.740613018e-03 lketa = -3.911472438e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.662082328e-01 lpclm = 2.467351305e-06 wpclm = 1.110223025e-22 ppclm = 1.110223025e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 3.668885335e-03 lpdiblc2 = -6.666176630e-9
+ pdiblcb = -9.883598245e-02 lpdiblcb = 1.519670040e-7
+ drout = 0.56
+ pscbe1 = -5.399535418e+07 lpscbe1 = 1.741697186e+3
+ pscbe2 = 4.685632485e-08 lpscbe2 = -7.719113680e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.151404795e+01 lbeta0 = -9.752188105e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.711119258e-10 lagidl = -2.898164661e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.817235263e-01 lkt1 = 2.635183383e-8
+ kt2 = -6.035456582e-02 lkt2 = 1.645005918e-8
+ at = 1.024940121e+05 lat = -4.795950233e-2
+ ute = -1.332981033e-01 lute = 1.351293641e-7
+ ua1 = 3.328055597e-09 lua1 = -1.056161454e-15
+ ub1 = -2.852522340e-18 lub1 = 2.458530043e-24
+ uc1 = 1.859730957e-11 luc1 = -9.937731742e-17 puc1 = 2.584939414e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.67 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.12e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.127136425e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.776911808e-9
+ k1 = 3.512559901e-01 lk1 = 1.745257769e-7
+ k2 = 5.719390124e-02 lk2 = -7.220885529e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.841659314e-01 ldsub = 1.122659537e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.937752555e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.671186683e-9
+ nfactor = {2.152613232e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.969208211e-7
+ eta0 = -2.317683150e-01 leta0 = 4.780476779e-07 weta0 = -2.168404345e-22 peta0 = 3.278627370e-28
+ etab = 8.728991787e-01 letab = -1.797601417e-06 wetab = 1.838806885e-22 petab = 7.459310947e-29
+ u0 = 9.740710576e-03 lu0 = 4.077017098e-10
+ ua = -8.760198240e-11 lua = -8.377855030e-16
+ ub = 1.194459582e-19 lub = 1.522494564e-24
+ uc = -7.526918424e-11 luc = 1.115271947e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.984839386e+04 lvsat = -1.319368033e-2
+ a0 = 1.446042456e+00 la0 = -7.857361509e-7
+ ags = 1.631988120e-01 lags = 6.468605781e-7
+ a1 = 0.0
+ a2 = 5.883765817e-01 la2 = 4.355569708e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.074975873e-02 lketa = -3.116565955e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.490103892e-01 lpclm = 3.778587940e-7
+ pdiblc1 = 7.614176700e-01 lpdiblc1 = -7.644407059e-7
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 9.440520000e-02 ldrout = 9.582732495e-7
+ pscbe1 = 7.985241057e+08 lpscbe1 = -1.293279044e+1
+ pscbe2 = 9.536577846e-09 lpscbe2 = -3.807531059e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.831389756e+00 lbeta0 = 1.943688500e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.694326460e-10 lagidl = 8.227161552e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.581851405e-01 lkt1 = -2.209416583e-8
+ kt2 = -5.638602898e-02 lkt2 = 8.282135728e-9
+ at = 9.763617505e+04 lat = -3.796124776e-2
+ ute = 9.699104623e-01 lute = -2.135461409e-06 wute = -2.220446049e-22 pute = -2.220446049e-28
+ ua1 = 6.248983323e-09 lua1 = -7.067927273e-15 pua1 = 6.617444900e-36
+ ub1 = -4.359386902e-18 lub1 = 5.559913481e-24
+ uc1 = -1.319123403e-10 luc1 = 2.103971287e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.68 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.12e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.163282379e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.702547591e-8
+ k1 = 5.163592603e-01 lk1 = -1.815505386e-10
+ k2 = -3.721282912e-02 lk2 = 2.768951457e-08 wk2 = 2.775557562e-23 pk2 = -1.387778781e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.350833910e+00 ldsub = -6.074482450e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.201588580e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.058952338e-8
+ nfactor = {2.786123308e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.267282178e-06 wnfactor = -3.552713679e-21
+ eta0 = -8.141180000e-02 leta0 = 3.189449244e-7
+ etab = -1.747153674e+00 letab = 9.748599102e-7
+ u0 = 1.757489028e-02 lu0 = -7.882192232e-09 pu0 = -1.387778781e-29
+ ua = 1.401704327e-10 lua = -1.078807440e-15
+ ub = 1.862301569e-18 lub = -3.217429574e-25
+ uc = -1.038019886e-10 luc = 4.134527707e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -4.078857788e+05 lvsat = 4.817485892e-01 wvsat = 1.164153218e-16
+ a0 = 6.889987434e-01 la0 = 1.534479470e-8
+ ags = 2.436803300e-01 lags = 5.616974502e-7
+ a1 = 0.0
+ a2 = 1.011042012e+00 la2 = -1.169490711e-8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.312283582e-02 lketa = -2.837782933e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.674890720e+00 lpclm = -9.193309952e-7
+ pdiblc1 = 7.025719961e-02 lpdiblc1 = -3.307543091e-08 ppdiblc1 = -5.551115123e-29
+ pdiblc2 = 8.652213951e-04 lpdiblc2 = -4.605382236e-10
+ pdiblcb = -3.110733092e-02 lpdiblcb = 6.462594361e-09 wpdiblcb = -5.551115123e-23
+ drout = 1.0
+ pscbe1 = 7.710109249e+08 lpscbe1 = 1.618083203e+1
+ pscbe2 = 9.007747976e-09 lpscbe2 = 1.788387980e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.458848501e+00 lbeta0 = 1.279730480e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 8.602477646e-10 lagidl = -3.726777648e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.131948081e-01 lkt1 = -6.970158589e-8
+ kt2 = -6.630249102e-02 lkt2 = 1.877543836e-8
+ at = 9.153536024e+04 lat = -3.150554856e-2
+ ute = -1.996613204e+00 lute = 1.003624939e-6
+ ua1 = -3.775967790e-09 lua1 = 3.540175246e-15 wua1 = 1.654361225e-30 pua1 = 3.308722450e-36
+ ub1 = 4.616188809e-18 lub1 = -3.937771469e-24 wub1 = -3.081487911e-39 pub1 = -3.081487911e-45
+ uc1 = 3.596775873e-10 luc1 = -3.097885850e-16 wuc1 = 2.067951531e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.69 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.12e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.078907267e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.018058955e-11
+ k1 = 4.909838222e-01 lk1 = 1.398225775e-8
+ k2 = 4.209442650e-02 lk2 = -1.657741630e-08 pk2 = 1.387778781e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -4.172892105e-01 ldsub = 3.794650372e-07 pdsub = -2.220446049e-28
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.478477057e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -9.772392518e-9
+ nfactor = {-5.870075767e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.154982881e-7
+ eta0 = 0.49
+ etab = -1.387720750e-03 letab = 4.257278410e-10
+ u0 = 7.618678736e-04 lu0 = 1.502332487e-9
+ ua = -3.376740709e-09 lua = 8.842268524e-16
+ ub = 2.824451866e-18 lub = -8.587863887e-25
+ uc = -6.643422899e-11 luc = 2.048771468e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.427631531e+05 lvsat = -2.721431252e-1
+ a0 = 8.685903852e-01 la0 = -8.489787201e-8
+ ags = 9.078080320e-01 lags = 1.910012908e-7
+ a1 = 0.0
+ a2 = 1.224409650e+00 la2 = -1.307903218e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -4.314918808e-02 lketa = 3.031526251e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -7.249963768e-01 lpclm = 4.202139854e-07 wpclm = 4.440892099e-22 ppclm = -1.665334537e-28
+ pdiblc1 = -4.793535710e-01 lpdiblc1 = 2.737008129e-07 wpdiblc1 = 1.387778781e-22 ppdiblc1 = 8.326672685e-29
+ pdiblc2 = -1.124292056e-02 lpdiblc2 = 6.297863373e-09 wpdiblc2 = 1.951563910e-24 ppdiblc2 = 4.336808690e-31
+ pdiblcb = 2.232572515e-01 lpdiblcb = -1.355160846e-07 wpdiblcb = 1.110223025e-22 ppdiblcb = -5.551115123e-29
+ drout = 1.629818715e+00 ldrout = -3.515459120e-7
+ pscbe1 = 8.000356861e+08 lpscbe1 = -1.991890262e-2
+ pscbe2 = 9.541728081e-09 lpscbe2 = -1.192128777e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.498743859e+00 lbeta0 = 1.411220881e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 3.066789197e-10 lagidl = -6.369224268e-17
+ bgidl = 6.790496970e+08 lbgidl = 1.791448306e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.635424940e-01 lkt1 = 1.421798196e-8
+ kt2 = -7.618700202e-03 lkt2 = -1.398009316e-8
+ at = -1.047669511e+04 lat = 2.543452038e-2
+ ute = 6.218841866e-01 lute = -4.579417499e-07 wute = 4.440892099e-22 pute = -2.220446049e-28
+ ua1 = 5.372180747e-09 lua1 = -1.566046823e-15
+ ub1 = -5.230148959e-18 lub1 = 1.558158882e-24
+ uc1 = -3.083411409e-10 luc1 = 6.307942852e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.70 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.12e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-4.572302168e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.916523970e-07 wvth0 = -8.160937497e-07 pvth0 = 2.514956109e-13
+ k1 = -4.718648500e+00 lk1 = 1.619434650e-06 wk1 = 4.010562175e-06 pk1 = -1.235934945e-12
+ k2 = 2.112067099e+00 lk2 = -6.544808947e-07 wk2 = -1.719256481e-06 pk2 = 5.298232698e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.853921239e+01 ldsub = -5.462360060e-06 wdsub = -1.903560441e-05 pdsub = 5.866202211e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {1.810835964e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.133799389e-07 wvoff = -2.188386413e-06 pvoff = 6.743950409e-13
+ nfactor = {3.418819145e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.010117480e-05 wnfactor = -3.590873003e-05 pnfactor = 1.106599333e-11
+ eta0 = 7.767654285e+00 leta0 = -2.242754721e-06 weta0 = -7.256052475e-06 peta0 = 2.236097691e-12
+ etab = 7.624397952e-01 letab = -2.349629977e-07 wetab = -7.905970781e-07 petab = 2.436383016e-13
+ u0 = -4.849529805e-03 lu0 = 3.231596910e-09 wu0 = 2.322699618e-08 pu0 = -7.157863414e-15
+ ua = 3.718909529e-09 lua = -1.302439681e-15 wua = 1.759278767e-15 pua = -5.421569377e-22
+ ub = -1.034097811e-17 lub = 3.198404168e-24 wub = 5.015930594e-24 pub = -1.545759331e-30
+ uc = 2.220670608e-10 luc = -6.841972778e-17 wuc = -1.953668734e-16 puc = 6.020620936e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.595835329e+05 lvsat = -2.465096616e-01 wvsat = -1.117101726e+00 pvsat = 3.442572388e-7
+ a0 = 6.838477503e+00 la0 = -1.924637985e-06 wa0 = -7.613731156e-06 pa0 = 2.346323530e-12
+ ags = 2.472114171e+00 lags = -2.910709322e-7
+ a1 = 0.0
+ a2 = -7.473993509e-01 la2 = 4.768620580e-07 wa2 = 2.417651634e-06 pa2 = -7.450477040e-13
+ b0 = 0.0
+ b1 = 0.0
+ keta = -6.989355254e-02 lketa = 1.127333704e-08 wketa = 9.998008542e-08 pketa = -3.081086292e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.129943055e-01 lpclm = 3.856983071e-07 wpclm = 1.138844354e-06 ppclm = -3.509576646e-13
+ pdiblc1 = 8.415054587e-01 lpdiblc1 = -1.333483143e-07 wpdiblc1 = -4.116424209e-07 ppdiblc1 = 1.268558449e-13
+ pdiblc2 = 6.617479122e-02 lpdiblc2 = -1.755995287e-08 wpdiblc2 = -6.171298503e-08 ppdiblc2 = 1.901809060e-14
+ pdiblcb = 2.114639687e+00 lpdiblcb = -7.183834098e-07 wpdiblcb = -2.709466543e-06 ppdiblcb = 8.349763046e-13
+ drout = -3.568266218e+00 ldrout = 1.250347922e-06 wdrout = 4.205366446e-06 pdrout = -1.295967778e-12
+ pscbe1 = 7.998725497e+08 lpscbe1 = 3.035483965e-2
+ pscbe2 = -5.598119199e-08 lpscbe2 = 2.007298540e-14 wpscbe2 = 7.635430186e-14 ppscbe2 = -2.353010520e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.144646343e+01 lbeta0 = -6.930676652e-06 wbeta0 = -2.437718832e-05 pbeta0 = 7.512318125e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -4.103040705e-08 lagidl = 1.267515754e-14 wagidl = 4.220918287e-14 pagidl = -1.300760389e-20
+ bgidl = 2.146251082e+09 lbgidl = -2.730026202e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.744252098e-01 lkt1 = -7.487929149e-08 wkt1 = -1.779532817e-07 pkt1 = 5.483986281e-14
+ kt2 = 2.029830968e-01 lkt2 = -7.888124893e-08 wkt2 = -3.006224105e-07 pkt2 = 9.264280824e-14
+ at = 7.700442191e+05 lat = -2.150986098e-01 wat = -6.501226557e-01 pat = 2.003482988e-7
+ ute = -2.066174858e+00 lute = 3.704374060e-07 wute = -9.283229527e-07 pute = 2.860812843e-13
+ ua1 = -6.132720519e-09 lua1 = 1.979418600e-15 wua1 = 6.998309390e-15 pua1 = -2.156669005e-21
+ ub1 = 1.257181891e-17 lub1 = -3.927873555e-24 wub1 = -1.512988460e-23 pub1 = 4.662576536e-30
+ uc1 = 1.563456106e-10 luc1 = -8.012308769e-17 wuc1 = -5.112597782e-16 puc1 = 1.575549259e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.71 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.12e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -3.7585e-8
+ vth0 = {-2.848938876e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.049602158e-07 wvth0 = 2.107656487e-06 pvth0 = -4.766065871e-13
+ k1 = 9.526687473e+00 lk1 = -1.899956392e-06 wk1 = -9.941914512e-06 pk1 = 2.236100476e-12
+ k2 = -3.993465707e+00 lk2 = 8.567526440e-07 wk2 = 4.456907691e-06 pk2 = -1.008331035e-12
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -4.316718685e+01 ldsub = 9.893371752e-06 wdsub = 5.122596412e-05 pdsub = -1.164372687e-11
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-4.604894873e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 9.799405185e-07 wvoff = 5.162968710e-06 pvoff = -1.153313555e-12
+ nfactor = {-5.945620173e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.307306753e-05 wnfactor = 7.085083425e-05 pnfactor = -1.538598078e-11
+ eta0 = -1.309098965e+01 leta0 = 2.919663030e-06 weta0 = 1.559898770e-05 peta0 = -3.436215653e-12
+ etab = -8.669614402e-01 letab = 1.640402236e-07 wetab = 9.889662081e-07 petab = -1.930625480e-13
+ u0 = 4.684905036e-02 lu0 = -9.729666201e-09 wu0 = -5.170278647e-08 pu0 = 1.145105820e-14
+ ua = 3.671726321e-09 lua = -1.383364944e-15 wua = -6.897567371e-15 pua = 1.628112637e-21
+ ub = 4.919305646e-18 lub = -4.672680658e-25 wub = -3.629403769e-24 pub = 5.499380665e-31
+ uc = 4.821827957e-10 luc = -1.396770950e-16 wuc = -5.868136054e-16 puc = 1.643890460e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.545403945e+06 lvsat = 6.047457283e-01 wvsat = 3.117596875e+00 pvsat = -7.117385521e-7
+ a0 = -1.174631282e+00 la0 = -1.730903262e-08 wa0 = 2.157899765e-06 pa0 = 2.037138129e-14
+ ags = 1.25
+ a1 = 0.0
+ a2 = 1.442889154e+01 la2 = -3.361634825e-06 wa2 = -1.621545333e-05 pa2 = 3.956381981e-12
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.777949702e+00 lketa = -7.146061625e-07 wketa = -3.325366867e-06 pketa = 8.410357140e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -2.407218296e+00 lpclm = 8.710606572e-07 wpclm = 3.682882740e-06 ppclm = -1.025170451e-12
+ pdiblc1 = -1.334820138e+01 lpdiblc1 = 3.477921100e-06 wpdiblc1 = 1.616221958e-05 ppdiblc1 = -4.093241857e-12
+ pdiblc2 = -4.024634266e-01 lpdiblc2 = 1.007690741e-07 wpdiblc2 = 4.829156792e-07 ppdiblc2 = -1.185973402e-13
+ pdiblcb = -1.223411646e+01 lpdiblcb = 2.891712221e-06 wpdiblcb = 1.413379336e-05 ppdiblcb = -3.403319731e-12
+ drout = 3.005724414e+01 ldrout = -7.240626739e-06 wdrout = -3.463197232e-05 pdrout = 8.521652903e-12
+ pscbe1 = 800000000.0
+ pscbe2 = 1.217401629e-07 lpscbe2 = -2.384341146e-14 wpscbe2 = -1.324142166e-13 ppscbe2 = 2.806183550e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -5.473606614e+01 lbeta0 = 1.456582444e-05 wbeta0 = 7.434667616e-05 pbeta0 = -1.714283923e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.951684681e-08 lagidl = -4.421663060e-15 wagidl = -3.279966535e-14 pagidl = 5.203952532e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -2.8385e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.00081386752815302
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207367379934e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.139261571e+00 lkt1 = 3.956262997e-07 wkt1 = 1.877051209e-06 pkt1 = -4.656212959e-13
+ kt2 = -3.088674796e+00 lkt2 = 7.554207424e-07 wkt2 = 3.572586507e-06 pkt2 = -8.890712910e-13
+ at = -1.741178401e+06 lat = 4.103368464e-01 wat = 2.083674966e+00 pat = -4.829344620e-7
+ ute = 1.298119362e+01 lute = -3.442758680e-06 wute = -1.560621360e-05 pute = 4.051858432e-12
+ ua1 = 3.269618732e-08 lua1 = -7.787267688e-15 wua1 = -3.797411487e-14 pua1 = 9.165006662e-21
+ ub1 = -5.067126034e-17 lub1 = 1.192950084e-23 wub1 = 5.946929237e-23 pub1 = -1.404009199e-29
+ uc1 = 5.545210808e-10 luc1 = -1.874445151e-16 wuc1 = -7.142881799e-16 puc1 = 2.206075736e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.72 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 1.0e-06 wmax = 1.12e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.149651792e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.052310473e-07 wvth0 = -1.776356839e-21
+ k1 = 4.276785563e-01 lk1 = 3.979367167e-7
+ k2 = 5.309370481e-02 lk2 = -6.710580081e-7
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -2.101213709e-06 lcit = 2.427282018e-10 wcit = -4.235164736e-28 pcit = -2.710505431e-32
+ voff = {-1.607085645e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.548662650e-07 wvoff = -2.220446049e-22
+ nfactor = {1.557178842e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.489901973e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 8.003413890e-03 lu0 = 2.669112821e-8
+ ua = -7.453530917e-10 lua = 4.106318926e-16
+ ub = 5.244028537e-19 lub = 1.093046418e-23
+ uc = -1.141591497e-10 luc = 8.501101883e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.005921802e+04 lvsat = 2.010847228e+0
+ a0 = 1.535439680e+00 la0 = -7.148123619e-6
+ ags = 6.310696593e-02 lags = 5.021222554e-6
+ a1 = 0.0
+ a2 = 1.012623611e+00 la2 = -4.264840540e-6
+ b0 = 7.164915408e-09 lb0 = -1.437150913e-13
+ b1 = 4.461843946e-08 lb1 = -8.949642438e-13
+ keta = 2.968747017e-02 lketa = -6.329891132e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.658133292e-02 lpclm = 3.159970378e-06 ppclm = 1.776356839e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 1.517320480e-03 lpdiblc2 = -2.403013816e-8
+ pdiblcb = -2.425209293e-01 lpdiblcb = 1.753112126e-6
+ drout = 0.56
+ pscbe1 = 8.000122229e+08 lpscbe1 = -1.223005743e+0
+ pscbe2 = 1.122278589e-08 lpscbe2 = -1.162836921e-13
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -2.507271250e-11 lalpha0 = 2.508729730e-15
+ alpha1 = -2.507271250e-11 lalpha1 = 2.508729730e-15
+ beta0 = 3.594760111e+01 lbeta0 = -5.951060825e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.265105400e-09 lagidl = -3.650602326e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -9.693353258e-02 legidl = 1.970480888e-05 pegidl = -1.065814104e-26
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.376177916e-01 lkt1 = -6.325762013e-8
+ kt2 = -6.009738111e-02 lkt2 = 1.552283545e-7
+ at = 8.878911860e+04 lat = -1.780947235e+0
+ ute = -7.062263283e-02 lute = -1.236455545e-6
+ ua1 = 2.157263413e-09 lua1 = -6.710242406e-15
+ ub1 = -1.357525803e-18 lub1 = 1.287006248e-23
+ uc1 = -3.506122186e-11 luc1 = 5.275288713e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.73 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.0e-06 wmax = 1.12e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.119478+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.44751769
+ k2 = 0.01963811
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.19335692+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.6314579+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0093341
+ ua = -7.2488104e-10
+ ub = 1.06934111e-18
+ uc = -7.1776909e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 160310.0
+ a0 = 1.17907
+ ags = 0.31344
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.0018702
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.14095898
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00031929802
+ pdiblcb = -0.15511953
+ drout = 0.56
+ pscbe1 = 799951250.0
+ pscbe2 = 5.4254628e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.2785893
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 4.4509773e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.88544965
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.4407715
+ kt2 = -0.052358472
+ at = 0.0
+ ute = -0.13226612
+ ua1 = 1.8227243e-9
+ ub1 = -7.1588888e-19
+ uc1 = -8.7612717e-12
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.74 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.0e-06 wmax = 1.12e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.119308571e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.365284442e-9
+ k1 = 4.557431136e-01 lk1 = -6.628186177e-8
+ k2 = 1.736465621e-02 lk2 = 1.831987716e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.866729821e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.386030771e-8
+ nfactor = {1.917980732e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.308849687e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 9.209108364e-03 lu0 = 1.007203851e-9
+ ua = -7.714556020e-10 lua = 3.753057380e-16
+ ub = 1.139159733e-18 lub = -5.626103368e-25
+ uc = -7.082993503e-11 luc = -7.630877232e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.687361861e+05 lvsat = -8.737166397e-01 wvsat = 4.656612873e-16
+ a0 = 1.298282802e+00 la0 = -9.606370240e-7
+ ags = 3.007947423e-01 lags = 1.018976364e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.275546728e-04 lketa = -8.401813297e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.415723457e-01 lpclm = -8.107596053e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -1.412456511e-03 lpdiblc2 = 1.395477241e-08 ppdiblc2 = 6.938893904e-30
+ pdiblcb = -2.502133320e-01 lpdiblcb = 7.662820228e-7
+ drout = 0.56
+ pscbe1 = 1.230892076e+09 lpscbe1 = -3.472594437e+3
+ pscbe2 = -1.731012336e-08 lpscbe2 = 1.832072184e-13 ppscbe2 = -5.293955920e-35
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.405041024e+00 lbeta0 = 2.315554051e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.940678393e-10 lagidl = -2.006243465e-15 wagidl = -8.271806126e-31 pagidl = 3.308722450e-36
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 1.682321702e+00 legidl = -6.421330460e-6
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.058118873e-01 lkt1 = -2.817105026e-7
+ kt2 = -4.835860979e-02 lkt2 = -3.223156969e-8
+ at = -9.199465573e+04 lat = 7.413085750e-1
+ ute = -1.650014701e-01 lute = 2.637870157e-7
+ ua1 = 5.595420866e-10 lua1 = 1.017893702e-14
+ ub1 = 8.371840607e-19 lub1 = -1.251492578e-23 pub1 = 6.162975822e-45
+ uc1 = -1.167338578e-11 luc1 = 2.346631032e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.75 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.0e-06 wmax = 1.12e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.116324143e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.347660345e-8
+ k1 = 4.428654258e-01 lk1 = -1.402201541e-8
+ k2 = 2.164134381e-02 lk2 = 9.643518320e-10
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.673887289e-01 ldsub = -1.247435718e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.076298863e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.118637217e-8
+ nfactor = {8.205595117e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.144672185e-6
+ eta0 = 1.618122575e-01 leta0 = -3.320080490e-7
+ etab = -1.415226926e-01 letab = 2.902512456e-7
+ u0 = 8.961795572e-03 lu0 = 2.010841203e-9
+ ua = -8.686534836e-10 lua = 7.697512652e-16
+ ub = 1.145979433e-18 lub = -5.902858386e-25
+ uc = -7.565336861e-11 luc = 1.194343622e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 53438.0
+ a0 = 1.058775121e+00 la0 = 1.132585948e-8
+ ags = 1.699111794e-01 lags = 6.330453849e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.740613019e-03 lketa = -3.911472438e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.662082328e-01 lpclm = 2.467351305e-06 wpclm = -1.110223025e-22 ppclm = 1.110223025e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 3.668885335e-03 lpdiblc2 = -6.666176630e-9
+ pdiblcb = -9.883598245e-02 lpdiblcb = 1.519670040e-7
+ drout = 0.56
+ pscbe1 = -5.399535418e+07 lpscbe1 = 1.741697186e+3
+ pscbe2 = 4.685632485e-08 lpscbe2 = -7.719113680e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.151404795e+01 lbeta0 = -9.752188105e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.711119258e-10 lagidl = -2.898164661e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.817235264e-01 lkt1 = 2.635183383e-8
+ kt2 = -6.035456581e-02 lkt2 = 1.645005918e-8
+ at = 1.024940121e+05 lat = -4.795950233e-2
+ ute = -1.332981033e-01 lute = 1.351293641e-7
+ ua1 = 3.328055597e-09 lua1 = -1.056161454e-15
+ ub1 = -2.852522339e-18 lub1 = 2.458530043e-24
+ uc1 = 1.859730957e-11 luc1 = -9.937731742e-17 wuc1 = 1.292469707e-32 puc1 = 2.584939414e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.76 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.0e-06 wmax = 1.12e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.127136425e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.776911808e-9
+ k1 = 3.512559901e-01 lk1 = 1.745257769e-7
+ k2 = 5.719390124e-02 lk2 = -7.220885529e-08 wk2 = 5.551115123e-23 pk2 = -5.551115123e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.841659314e-01 ldsub = 1.122659537e-06 pdsub = 8.881784197e-28
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.937752555e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.671186683e-9
+ nfactor = {2.152613232e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.969208211e-07 wnfactor = -3.552713679e-21
+ eta0 = -2.317683150e-01 leta0 = 4.780476779e-07 weta0 = -2.602085214e-23 peta0 = 1.994931997e-28
+ etab = 8.728991787e-01 letab = -1.797601417e-06 wetab = 3.209238431e-22 petab = 1.387778781e-28
+ u0 = 9.740710576e-03 lu0 = 4.077017098e-10
+ ua = -8.760198240e-11 lua = -8.377855030e-16
+ ub = 1.194459582e-19 lub = 1.522494564e-24
+ uc = -7.526918424e-11 luc = 1.115271947e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.984839386e+04 lvsat = -1.319368033e-2
+ a0 = 1.446042456e+00 la0 = -7.857361509e-7
+ ags = 1.631988120e-01 lags = 6.468605781e-7
+ a1 = 0.0
+ a2 = 5.883765817e-01 la2 = 4.355569708e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.074975873e-02 lketa = -3.116565955e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.490103892e-01 lpclm = 3.778587940e-7
+ pdiblc1 = 7.614176700e-01 lpdiblc1 = -7.644407059e-07 ppdiblc1 = -8.881784197e-28
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 9.440520000e-02 ldrout = 9.582732495e-7
+ pscbe1 = 7.985241057e+08 lpscbe1 = -1.293279044e+1
+ pscbe2 = 9.536577846e-09 lpscbe2 = -3.807531059e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.831389756e+00 lbeta0 = 1.943688500e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.694326460e-10 lagidl = 8.227161552e-16 pagidl = 4.135903063e-37
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.581851405e-01 lkt1 = -2.209416583e-8
+ kt2 = -5.638602898e-02 lkt2 = 8.282135728e-9
+ at = 9.763617505e+04 lat = -3.796124776e-2
+ ute = 9.699104623e-01 lute = -2.135461409e-06 wute = 2.220446049e-22 pute = 8.881784197e-28
+ ua1 = 6.248983323e-09 lua1 = -7.067927273e-15
+ ub1 = -4.359386902e-18 lub1 = 5.559913481e-24 pub1 = 6.162975822e-45
+ uc1 = -1.319123403e-10 luc1 = 2.103971287e-16 wuc1 = 1.033975766e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.77 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.0e-06 wmax = 1.12e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.163282379e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.702547591e-8
+ k1 = 5.163592603e-01 lk1 = -1.815505386e-10
+ k2 = -3.721282912e-02 lk2 = 2.768951457e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.350833910e+00 ldsub = -6.074482450e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.201588580e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.058952338e-8
+ nfactor = {2.786123308e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.267282178e-6
+ eta0 = -8.141180000e-02 leta0 = 3.189449244e-7
+ etab = -1.747153674e+00 letab = 9.748599102e-7
+ u0 = 1.757489028e-02 lu0 = -7.882192232e-9
+ ua = 1.401704327e-10 lua = -1.078807440e-15
+ ub = 1.862301569e-18 lub = -3.217429574e-25
+ uc = -1.038019886e-10 luc = 4.134527707e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -4.078857788e+05 lvsat = 4.817485892e-01 wvsat = -1.164153218e-16 pvsat = -1.164153218e-22
+ a0 = 6.889987434e-01 la0 = 1.534479470e-8
+ ags = 2.436803300e-01 lags = 5.616974502e-7
+ a1 = 0.0
+ a2 = 1.011042012e+00 la2 = -1.169490711e-8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.312283582e-02 lketa = -2.837782933e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.674890720e+00 lpclm = -9.193309952e-7
+ pdiblc1 = 7.025719961e-02 lpdiblc1 = -3.307543091e-8
+ pdiblc2 = 8.652213951e-04 lpdiblc2 = -4.605382236e-10
+ pdiblcb = -3.110733092e-02 lpdiblcb = 6.462594361e-9
+ drout = 1.0
+ pscbe1 = 7.710109249e+08 lpscbe1 = 1.618083203e+1
+ pscbe2 = 9.007747976e-09 lpscbe2 = 1.788387980e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.458848501e+00 lbeta0 = 1.279730480e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 8.602477646e-10 lagidl = -3.726777648e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.131948081e-01 lkt1 = -6.970158589e-8
+ kt2 = -6.630249102e-02 lkt2 = 1.877543836e-8
+ at = 9.153536024e+04 lat = -3.150554856e-02 wat = -1.164153218e-16
+ ute = -1.996613204e+00 lute = 1.003624939e-6
+ ua1 = -3.775967790e-09 lua1 = 3.540175246e-15
+ ub1 = 4.616188809e-18 lub1 = -3.937771469e-24 wub1 = 3.081487911e-39 pub1 = -1.540743956e-45
+ uc1 = 3.596775873e-10 luc1 = -3.097885850e-16 wuc1 = 2.067951531e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.78 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.0e-06 wmax = 1.12e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.078907267e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.018058955e-11
+ k1 = 4.909838222e-01 lk1 = 1.398225775e-8
+ k2 = 4.209442650e-02 lk2 = -1.657741630e-08 wk2 = -2.775557562e-23
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -4.172892105e-01 ldsub = 3.794650372e-07 pdsub = -2.220446049e-28
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.478477057e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -9.772392518e-9
+ nfactor = {-5.870075767e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.154982881e-7
+ eta0 = 0.49
+ etab = -1.387720750e-03 letab = 4.257278410e-10
+ u0 = 7.618678736e-04 lu0 = 1.502332487e-9
+ ua = -3.376740709e-09 lua = 8.842268524e-16
+ ub = 2.824451866e-18 lub = -8.587863887e-25
+ uc = -6.643422899e-11 luc = 2.048771468e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.427631531e+05 lvsat = -2.721431252e-1
+ a0 = 8.685903852e-01 la0 = -8.489787201e-8
+ ags = 9.078080320e-01 lags = 1.910012908e-7
+ a1 = 0.0
+ a2 = 1.224409650e+00 la2 = -1.307903218e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -4.314918808e-02 lketa = 3.031526251e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -7.249963768e-01 lpclm = 4.202139854e-07 wpclm = -2.775557562e-22 ppclm = -8.326672685e-29
+ pdiblc1 = -4.793535710e-01 lpdiblc1 = 2.737008129e-07 wpdiblc1 = -2.220446049e-22 ppdiblc1 = -1.318389842e-28
+ pdiblc2 = -1.124292056e-02 lpdiblc2 = 6.297863373e-09 wpdiblc2 = 6.505213035e-24 ppdiblc2 = 7.047314121e-31
+ pdiblcb = 2.232572515e-01 lpdiblcb = -1.355160846e-07 wpdiblcb = 1.110223025e-22 ppdiblcb = 1.387778781e-29
+ drout = 1.629818715e+00 ldrout = -3.515459120e-7
+ pscbe1 = 8.000356861e+08 lpscbe1 = -1.991890262e-2
+ pscbe2 = 9.541728081e-09 lpscbe2 = -1.192128777e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.498743859e+00 lbeta0 = 1.411220881e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 3.066789197e-10 lagidl = -6.369224268e-17 wagidl = -4.135903063e-31
+ bgidl = 6.790496970e+08 lbgidl = 1.791448306e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.635424940e-01 lkt1 = 1.421798196e-8
+ kt2 = -7.618700202e-03 lkt2 = -1.398009316e-8
+ at = -1.047669511e+04 lat = 2.543452038e-2
+ ute = 6.218841866e-01 lute = -4.579417499e-7
+ ua1 = 5.372180747e-09 lua1 = -1.566046823e-15 pua1 = 1.654361225e-36
+ ub1 = -5.230148959e-18 lub1 = 1.558158882e-24
+ uc1 = -3.083411409e-10 luc1 = 6.307942852e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.79 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.0e-06 wmax = 1.12e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.244265066e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.088813240e-8
+ k1 = -8.508916437e-01 lk1 = 4.275080201e-7
+ k2 = 4.540287111e-01 lk2 = -1.435232048e-07 wk2 = 1.665334537e-22 pk2 = -6.938893904e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.814145886e-01 ldsub = 1.949624874e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.996279025e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.700171071e-8
+ nfactor = {-4.419254060e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.707883156e-7
+ eta0 = 7.699702980e-01 leta0 = -8.627844675e-8
+ etab = -6.25e-6
+ u0 = 1.755041559e-02 lu0 = -3.671394264e-9
+ ua = 5.415545117e-09 lua = -1.825291870e-15 wua = 3.308722450e-30 pua = -8.271806126e-37
+ ub = -5.503651299e-18 lub = 1.707685164e-24 wub = -1.540743956e-39 pub = 4.333342375e-46
+ uc = 3.365667565e-11 luc = -1.035729940e-17 wuc = 9.289626020e-33 puc = 6.310887242e-39
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.177412087e+05 lvsat = 8.548950402e-02 pvsat = -5.820766091e-23
+ a0 = -5.041491900e-01 la0 = 3.381392829e-7
+ ags = 2.472114171e+00 lags = -2.910709322e-7
+ a1 = 0.0
+ a2 = 1.584166219e+00 la2 = -2.416565037e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.652651129e-02 lketa = -1.844043402e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.852988681e-01 lpclm = 4.723729973e-8
+ pdiblc1 = 4.445205159e-01 lpdiblc1 = -1.100946442e-8
+ pdiblc2 = 6.659239392e-03 lpdiblc2 = 7.809547401e-10
+ pdiblcb = -4.983500488e-01 lpdiblcb = 8.686163714e-8
+ drout = 4.873584535e-01 ldrout = 5.260666719e-10
+ pscbe1 = 7.998725497e+08 lpscbe1 = 3.035483965e-2
+ pscbe2 = 1.765433880e-08 lpscbe2 = -2.619276124e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.937281138e+00 lbeta0 = 3.141480549e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -3.241795111e-10 lagidl = 1.307193999e-16
+ bgidl = 2.146251082e+09 lbgidl = -2.730026202e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.460420544e-01 lkt1 = -2.199212851e-8
+ kt2 = -8.693495928e-02 lkt2 = 1.046279840e-8
+ at = 1.430706804e+05 lat = -2.188417433e-2
+ ute = -2.961442731e+00 lute = 6.463321062e-7
+ ua1 = 6.163979206e-10 lua1 = -1.004572290e-16
+ ub1 = -2.019331242e-18 lub1 = 5.686811864e-25 wub1 = -7.703719778e-40 pub1 = 3.851859889e-46
+ uc1 = -3.367095838e-10 luc1 = 7.182173155e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.80 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.0e-06 wmax = 1.12e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -3.7585e-8
+ vth0 = {-8.163313737e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -5.467543570e-08 wvth0 = 1.050561053e-12 pvth0 = -2.680716626e-19
+ k1 = -6.122276825e-02 lk1 = 2.565227042e-07 wk1 = 5.513146135e-13 pk1 = -1.406789494e-19
+ k2 = 3.047439370e-01 lk2 = -1.156745491e-07 wk2 = -4.492352623e-13 pk2 = 1.146313617e-19
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 6.234759321e+00 ldsub = -1.335753536e-06 wdsub = -7.160708293e-13 pdsub = 1.827197966e-19
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {3.742322261e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.323060854e-07 wvoff = 2.280268491e-12 pvoff = -5.818561108e-19
+ nfactor = {8.871857503e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.765068176e-06 wnfactor = -3.358624133e-11 pnfactor = 8.570201196e-18
+ eta0 = 1.952570675e+00 leta0 = -3.942009323e-07 weta0 = -1.095308938e-11 peta0 = 2.794899816e-18
+ etab = 8.678913516e-02 letab = -2.214757843e-08 wetab = 1.253977103e-12 petab = -3.199773374e-19
+ u0 = -3.012757077e-03 lu0 = 1.313655241e-09 wu0 = 1.862281274e-14 pu0 = -4.751983126e-21
+ ua = -2.980241684e-09 lua = 1.867761173e-16 wua = 4.596666804e-21 pua = -1.172931468e-27
+ ub = 1.419139632e-18 lub = 6.308704882e-26 wub = -4.625850347e-30 pub = 1.180378230e-36
+ uc = -8.373631094e-11 luc = 1.885858995e-17 wuc = 3.664653722e-22 puc = -9.351096903e-29
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.611846143e+05 lvsat = -8.164996368e-02 wvsat = -9.471086636e-07 pvsat = 2.416737173e-13
+ a0 = 9.064192342e-01 la0 = 2.340104320e-09 wa0 = 1.270166973e-11 pa0 = -3.241085066e-18
+ ags = 1.25
+ a1 = 0.0
+ a2 = -1.209170084e+00 la2 = 4.538702625e-07 wa2 = -3.194329146e-12 pa2 = 8.150969677e-19
+ b0 = 0.0
+ b1 = 0.0
+ keta = -4.290231040e-01 lketa = 9.648592761e-08 wketa = 1.378797894e-11 pketa = -3.518278587e-18
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.144525300e+00 lpclm = -1.176058244e-07 wpclm = 1.666924433e-12 ppclm = -4.253491070e-19
+ pdiblc1 = 2.238540380e+00 lpdiblc1 = -4.695753422e-07 wpdiblc1 = -1.586795589e-11 ppdiblc1 = 4.049026303e-18
+ pdiblc2 = 6.325670189e-02 lpdiblc2 = -1.360527710e-08 wpdiblc2 = 2.321298493e-13 ppdiblc2 = -5.923257368e-20
+ pdiblcb = 1.396363005e+00 lpdiblcb = -3.904123186e-07 wpdiblcb = 4.933473054e-11 ppdiblcb = -1.258874319e-17
+ drout = -3.341622739e+00 ldrout = 9.776047470e-07 wdrout = 4.752114189e-11 pdrout = -1.212596978e-17
+ pscbe1 = 800000000.0
+ pscbe2 = -5.958908092e-09 lpscbe2 = 3.219158476e-15 wpscbe2 = -2.404644881e-19 ppscbe2 = 6.135932343e-26
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.696329718e+01 lbeta0 = -1.966597328e-06 wbeta0 = 2.894960755e-11 pbeta0 = -7.387071378e-18
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.115301538e-09 lagidl = 5.970904430e-16 wagidl = 4.051726842e-19 pagidl = -1.033879138e-25
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -2.8385e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.290482065e-01 lkt1 = -5.341519375e-08 wkt1 = 1.145980534e-12 pkt1 = -2.924198537e-19
+ kt2 = 3.566996392e-01 lkt2 = -1.019926328e-07 wkt2 = 1.956205383e-12 pkt2 = -4.991649276e-19
+ at = 2.683032014e+05 lat = -5.540179629e-02 wat = -7.168273050e-07 pat = 1.829128234e-13
+ ute = -2.069320434e+00 lute = 4.648228862e-07 wute = -4.461409659e-12 pute = 1.138417903e-18
+ ua1 = -3.925739113e-09 lua1 = 1.051389483e-15 wua1 = -3.366643843e-20 pua1 = 8.590665094e-27
+ ub1 = 6.680453425e-18 lub1 = -1.610651776e-24 wub1 = 3.862871181e-29 pub1 = -9.856888391e-36
+ uc1 = -1.343358286e-10 luc1 = 2.530848236e-17 wuc1 = 2.704205952e-21 puc1 = -6.900322328e-28
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.81 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 9.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.149651792e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.052310473e-7
+ k1 = 4.276785563e-01 lk1 = 3.979367167e-7
+ k2 = 5.309370481e-02 lk2 = -6.710580081e-7
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -2.101213709e-06 lcit = 2.427282018e-10 wcit = 8.470329473e-28 pcit = 1.490777987e-31
+ voff = {-1.607085645e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.548662650e-7
+ nfactor = {1.557178842e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.489901973e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 8.003413890e-03 lu0 = 2.669112821e-8
+ ua = -7.453530917e-10 lua = 4.106318926e-16
+ ub = 5.244028537e-19 lub = 1.093046418e-23
+ uc = -1.141591497e-10 luc = 8.501101883e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.005921802e+04 lvsat = 2.010847228e+0
+ a0 = 1.535439680e+00 la0 = -7.148123619e-6
+ ags = 6.310696593e-02 lags = 5.021222554e-6
+ a1 = 0.0
+ a2 = 1.012623611e+00 la2 = -4.264840540e-6
+ b0 = 7.164915408e-09 lb0 = -1.437150913e-13
+ b1 = 4.461843946e-08 lb1 = -8.949642438e-13
+ keta = 2.968747017e-02 lketa = -6.329891132e-07 pketa = -8.881784197e-28
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.658133292e-02 lpclm = 3.159970378e-06 ppclm = 8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 1.517320480e-03 lpdiblc2 = -2.403013816e-8
+ pdiblcb = -2.425209293e-01 lpdiblcb = 1.753112126e-6
+ drout = 0.56
+ pscbe1 = 8.000122229e+08 lpscbe1 = -1.223005743e+0
+ pscbe2 = 1.122278589e-08 lpscbe2 = -1.162836921e-13
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -2.507271250e-11 lalpha0 = 2.508729730e-15
+ alpha1 = -2.507271250e-11 lalpha1 = 2.508729730e-15
+ beta0 = 3.594760111e+01 lbeta0 = -5.951060825e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.265105400e-09 lagidl = -3.650602326e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -9.693353258e-02 legidl = 1.970480888e-05 pegidl = 2.131628207e-26
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.376177916e-01 lkt1 = -6.325762013e-08 wkt1 = -8.881784197e-22
+ kt2 = -6.009738111e-02 lkt2 = 1.552283545e-7
+ at = 8.878911860e+04 lat = -1.780947235e+0
+ ute = -7.062263283e-02 lute = -1.236455545e-6
+ ua1 = 2.157263413e-09 lua1 = -6.710242406e-15
+ ub1 = -1.357525803e-18 lub1 = 1.287006248e-23
+ uc1 = -3.506122186e-11 luc1 = 5.275288713e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.82 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 9.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.119478+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.44751769
+ k2 = 0.01963811
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.19335692+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.6314579+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0093341
+ ua = -7.2488104e-10
+ ub = 1.06934111e-18
+ uc = -7.1776909e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 160310.0
+ a0 = 1.17907
+ ags = 0.31344
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.0018702
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.14095898
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00031929802
+ pdiblcb = -0.15511953
+ drout = 0.56
+ pscbe1 = 799951250.0
+ pscbe2 = 5.4254628e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.2785893
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 4.4509773e-10
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.88544965
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.4407715
+ kt2 = -0.052358472
+ at = 0.0
+ ute = -0.13226612
+ ua1 = 1.8227243e-9
+ ub1 = -7.1588888e-19
+ uc1 = -8.7612717e-12
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.83 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 9.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.119308571e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.365284442e-9
+ k1 = 4.557431136e-01 lk1 = -6.628186177e-8
+ k2 = 1.736465621e-02 lk2 = 1.831987716e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.866729821e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.386030771e-8
+ nfactor = {1.917980732e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.308849687e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 9.209108364e-03 lu0 = 1.007203851e-9
+ ua = -7.714556020e-10 lua = 3.753057380e-16
+ ub = 1.139159733e-18 lub = -5.626103368e-25
+ uc = -7.082993503e-11 luc = -7.630877232e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.687361861e+05 lvsat = -8.737166397e-1
+ a0 = 1.298282802e+00 la0 = -9.606370240e-7
+ ags = 3.007947423e-01 lags = 1.018976364e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.275546728e-04 lketa = -8.401813297e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.415723457e-01 lpclm = -8.107596053e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -1.412456511e-03 lpdiblc2 = 1.395477241e-08 ppdiblc2 = -6.938893904e-30
+ pdiblcb = -2.502133320e-01 lpdiblcb = 7.662820228e-7
+ drout = 0.56
+ pscbe1 = 1.230892076e+09 lpscbe1 = -3.472594437e+3
+ pscbe2 = -1.731012336e-08 lpscbe2 = 1.832072184e-13 ppscbe2 = -2.117582368e-34
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.405041024e+00 lbeta0 = 2.315554051e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.940678393e-10 lagidl = -2.006243465e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 1.682321702e+00 legidl = -6.421330460e-6
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.058118873e-01 lkt1 = -2.817105026e-7
+ kt2 = -4.835860979e-02 lkt2 = -3.223156969e-8
+ at = -9.199465573e+04 lat = 7.413085750e-1
+ ute = -1.650014701e-01 lute = 2.637870157e-7
+ ua1 = 5.595420866e-10 lua1 = 1.017893702e-14
+ ub1 = 8.371840607e-19 lub1 = -1.251492578e-23
+ uc1 = -1.167338578e-11 luc1 = 2.346631032e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.84 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 9.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.116324143e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.347660345e-8
+ k1 = 4.428654258e-01 lk1 = -1.402201541e-8
+ k2 = 2.164134381e-02 lk2 = 9.643518320e-10
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.673887289e-01 ldsub = -1.247435718e-06 pdsub = 3.552713679e-27
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.076298863e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.118637217e-8
+ nfactor = {8.205595117e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.144672185e-6
+ eta0 = 1.618122575e-01 leta0 = -3.320080490e-7
+ etab = -1.415226926e-01 letab = 2.902512456e-7
+ u0 = 8.961795573e-03 lu0 = 2.010841203e-9
+ ua = -8.686534836e-10 lua = 7.697512652e-16
+ ub = 1.145979433e-18 lub = -5.902858386e-25
+ uc = -7.565336861e-11 luc = 1.194343622e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 53438.0
+ a0 = 1.058775121e+00 la0 = 1.132585948e-8
+ ags = 1.699111794e-01 lags = 6.330453849e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.740613018e-03 lketa = -3.911472438e-08 pketa = -2.775557562e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.662082328e-01 lpclm = 2.467351305e-06 wpclm = 2.220446049e-22 ppclm = 1.332267630e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 3.668885335e-03 lpdiblc2 = -6.666176630e-9
+ pdiblcb = -9.883598245e-02 lpdiblcb = 1.519670040e-7
+ drout = 0.56
+ pscbe1 = -5.399535418e+07 lpscbe1 = 1.741697186e+3
+ pscbe2 = 4.685632485e-08 lpscbe2 = -7.719113680e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.151404795e+01 lbeta0 = -9.752188105e-06 wbeta0 = -2.842170943e-20
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.711119258e-10 lagidl = -2.898164661e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.817235263e-01 lkt1 = 2.635183383e-8
+ kt2 = -6.035456581e-02 lkt2 = 1.645005918e-8
+ at = 1.024940121e+05 lat = -4.795950233e-2
+ ute = -1.332981033e-01 lute = 1.351293641e-7
+ ua1 = 3.328055597e-09 lua1 = -1.056161454e-15
+ ub1 = -2.852522340e-18 lub1 = 2.458530043e-24
+ uc1 = 1.859730957e-11 luc1 = -9.937731742e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.85 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 9.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.127136425e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.776911808e-9
+ k1 = 3.512559901e-01 lk1 = 1.745257769e-7
+ k2 = 5.719390124e-02 lk2 = -7.220885529e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.841659314e-01 ldsub = 1.122659537e-06 pdsub = -8.881784197e-28
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.937752555e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.671186683e-9
+ nfactor = {2.152613232e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.969208211e-7
+ eta0 = -2.317683150e-01 leta0 = 4.780476779e-07 weta0 = 8.500145032e-23 peta0 = -3.191891196e-28
+ etab = 8.728991787e-01 letab = -1.797601417e-06 wetab = -2.289834988e-22 petab = -8.291978215e-28
+ u0 = 9.740710576e-03 lu0 = 4.077017098e-10
+ ua = -8.760198240e-11 lua = -8.377855030e-16
+ ub = 1.194459582e-19 lub = 1.522494564e-24
+ uc = -7.526918424e-11 luc = 1.115271947e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.984839386e+04 lvsat = -1.319368033e-2
+ a0 = 1.446042456e+00 la0 = -7.857361509e-7
+ ags = 1.631988120e-01 lags = 6.468605781e-7
+ a1 = 0.0
+ a2 = 5.883765817e-01 la2 = 4.355569708e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.074975873e-02 lketa = -3.116565955e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.490103892e-01 lpclm = 3.778587940e-7
+ pdiblc1 = 7.614176700e-01 lpdiblc1 = -7.644407059e-7
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 9.440520000e-02 ldrout = 9.582732495e-7
+ pscbe1 = 7.985241057e+08 lpscbe1 = -1.293279044e+1
+ pscbe2 = 9.536577846e-09 lpscbe2 = -3.807531059e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.831389756e+00 lbeta0 = 1.943688500e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.694326460e-10 lagidl = 8.227161552e-16 pagidl = 4.135903063e-37
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.581851405e-01 lkt1 = -2.209416583e-8
+ kt2 = -5.638602898e-02 lkt2 = 8.282135728e-9
+ at = 9.763617505e+04 lat = -3.796124776e-2
+ ute = 9.699104623e-01 lute = -2.135461409e-06 wute = 6.661338148e-22 pute = -1.776356839e-27
+ ua1 = 6.248983323e-09 lua1 = -7.067927273e-15
+ ub1 = -4.359386902e-18 lub1 = 5.559913481e-24 pub1 = 6.162975822e-45
+ uc1 = -1.319123403e-10 luc1 = 2.103971287e-16 puc1 = 1.033975766e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.86 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 9.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.163282379e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.702547591e-8
+ k1 = 5.163592603e-01 lk1 = -1.815505386e-10
+ k2 = -3.721282912e-02 lk2 = 2.768951457e-08 wk2 = -5.551115123e-23
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.350833910e+00 ldsub = -6.074482450e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.201588580e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.058952338e-8
+ nfactor = {2.786123308e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.267282178e-6
+ eta0 = -8.141180000e-02 leta0 = 3.189449244e-7
+ etab = -1.747153674e+00 letab = 9.748599102e-7
+ u0 = 1.757489028e-02 lu0 = -7.882192232e-9
+ ua = 1.401704327e-10 lua = -1.078807440e-15
+ ub = 1.862301569e-18 lub = -3.217429574e-25
+ uc = -1.038019886e-10 luc = 4.134527707e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -4.078857788e+05 lvsat = 4.817485892e-01 wvsat = 2.328306437e-16 pvsat = -3.492459655e-22
+ a0 = 6.889987434e-01 la0 = 1.534479470e-8
+ ags = 2.436803300e-01 lags = 5.616974502e-7
+ a1 = 0.0
+ a2 = 1.011042012e+00 la2 = -1.169490711e-8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.312283582e-02 lketa = -2.837782933e-08 pketa = 2.775557562e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.674890720e+00 lpclm = -9.193309952e-7
+ pdiblc1 = 7.025719961e-02 lpdiblc1 = -3.307543091e-8
+ pdiblc2 = 8.652213951e-04 lpdiblc2 = -4.605382236e-10
+ pdiblcb = -3.110733092e-02 lpdiblcb = 6.462594361e-9
+ drout = 1.0
+ pscbe1 = 7.710109249e+08 lpscbe1 = 1.618083203e+1
+ pscbe2 = 9.007747976e-09 lpscbe2 = 1.788387980e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.458848501e+00 lbeta0 = 1.279730480e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 8.602477646e-10 lagidl = -3.726777648e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.131948081e-01 lkt1 = -6.970158589e-8
+ kt2 = -6.630249102e-02 lkt2 = 1.877543836e-8
+ at = 9.153536024e+04 lat = -3.150554856e-2
+ ute = -1.996613204e+00 lute = 1.003624939e-6
+ ua1 = -3.775967790e-09 lua1 = 3.540175246e-15 wua1 = -1.654361225e-30 pua1 = 2.481541838e-36
+ ub1 = 4.616188809e-18 lub1 = -3.937771469e-24 wub1 = 3.081487911e-39 pub1 = 3.081487911e-45
+ uc1 = 3.596775873e-10 luc1 = -3.097885850e-16 wuc1 = -2.067951531e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.87 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 9.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.078907267e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.018058955e-11
+ k1 = 4.909838222e-01 lk1 = 1.398225775e-8
+ k2 = 4.209442650e-02 lk2 = -1.657741630e-08 wk2 = -5.551115123e-23
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -4.172892105e-01 ldsub = 3.794650372e-07 pdsub = -4.440892099e-28
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.478477057e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -9.772392518e-9
+ nfactor = {-5.870075767e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.154982881e-7
+ eta0 = 0.49
+ etab = -1.387720750e-03 letab = 4.257278410e-10
+ u0 = 7.618678736e-04 lu0 = 1.502332487e-9
+ ua = -3.376740709e-09 lua = 8.842268524e-16 wua = -6.617444900e-30
+ ub = 2.824451866e-18 lub = -8.587863887e-25
+ uc = -6.643422899e-11 luc = 2.048771468e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.427631531e+05 lvsat = -2.721431252e-1
+ a0 = 8.685903852e-01 la0 = -8.489787201e-8
+ ags = 9.078080320e-01 lags = 1.910012908e-7
+ a1 = 0.0
+ a2 = 1.224409650e+00 la2 = -1.307903218e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -4.314918808e-02 lketa = 3.031526251e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -7.249963768e-01 lpclm = 4.202139854e-07 wpclm = 7.771561172e-22 ppclm = -5.551115123e-29
+ pdiblc1 = -4.793535710e-01 lpdiblc1 = 2.737008129e-07 wpdiblc1 = 4.440892099e-22 ppdiblc1 = -1.249000903e-28
+ pdiblc2 = -1.124292056e-02 lpdiblc2 = 6.297863373e-09 wpdiblc2 = -1.322726650e-23 ppdiblc2 = -6.613633252e-30
+ pdiblcb = 2.232572515e-01 lpdiblcb = -1.355160846e-07 ppdiblcb = 8.326672685e-29
+ drout = 1.629818715e+00 ldrout = -3.515459120e-7
+ pscbe1 = 8.000356861e+08 lpscbe1 = -1.991890262e-2
+ pscbe2 = 9.541728081e-09 lpscbe2 = -1.192128777e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.498743859e+00 lbeta0 = 1.411220881e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 3.066789197e-10 lagidl = -6.369224268e-17
+ bgidl = 6.790496970e+08 lbgidl = 1.791448306e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.635424940e-01 lkt1 = 1.421798196e-8
+ kt2 = -7.618700202e-03 lkt2 = -1.398009316e-8
+ at = -1.047669511e+04 lat = 2.543452038e-2
+ ute = 6.218841866e-01 lute = -4.579417499e-07 wute = -8.881784197e-22
+ ua1 = 5.372180747e-09 lua1 = -1.566046823e-15
+ ub1 = -5.230148959e-18 lub1 = 1.558158882e-24
+ uc1 = -3.083411409e-10 luc1 = 6.307942852e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.88 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 9.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.244265066e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.088813240e-8
+ k1 = -8.508916437e-01 lk1 = 4.275080201e-7
+ k2 = 4.540287111e-01 lk2 = -1.435232048e-07 wk2 = 4.440892099e-22 pk2 = 5.551115123e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.814145886e-01 ldsub = 1.949624874e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.996279025e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.700171071e-8
+ nfactor = {-4.419254060e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.707883156e-7
+ eta0 = 7.699702980e-01 leta0 = -8.627844675e-8
+ etab = -6.25e-6
+ u0 = 1.755041559e-02 lu0 = -3.671394264e-9
+ ua = 5.415545117e-09 lua = -1.825291870e-15 wua = -3.308722450e-30 pua = 8.271806126e-37
+ ub = -5.503651299e-18 lub = 1.707685164e-24 wub = 7.703719778e-40 pub = -3.851859889e-46
+ uc = 3.365667565e-11 luc = -1.035729940e-17 wuc = -2.584939414e-32 puc = -1.241982609e-38
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.177412087e+05 lvsat = 8.548950402e-02 pvsat = 1.164153218e-22
+ a0 = -5.041491900e-01 la0 = 3.381392829e-7
+ ags = 2.472114171e+00 lags = -2.910709322e-7
+ a1 = 0.0
+ a2 = 1.584166219e+00 la2 = -2.416565037e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.652651129e-02 lketa = -1.844043402e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.852988681e-01 lpclm = 4.723729973e-8
+ pdiblc1 = 4.445205159e-01 lpdiblc1 = -1.100946442e-8
+ pdiblc2 = 6.659239392e-03 lpdiblc2 = 7.809547401e-10
+ pdiblcb = -4.983500488e-01 lpdiblcb = 8.686163714e-8
+ drout = 4.873584535e-01 ldrout = 5.260666719e-10
+ pscbe1 = 7.998725497e+08 lpscbe1 = 3.035483965e-2
+ pscbe2 = 1.765433880e-08 lpscbe2 = -2.619276124e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.937281138e+00 lbeta0 = 3.141480549e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -3.241795111e-10 lagidl = 1.307193999e-16
+ bgidl = 2.146251082e+09 lbgidl = -2.730026202e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.460420544e-01 lkt1 = -2.199212851e-8
+ kt2 = -8.693495928e-02 lkt2 = 1.046279840e-8
+ at = 1.430706804e+05 lat = -2.188417433e-2
+ ute = -2.961442731e+00 lute = 6.463321062e-7
+ ua1 = 6.163979206e-10 lua1 = -1.004572290e-16
+ ub1 = -2.019331242e-18 lub1 = 5.686811864e-25 pub1 = 7.703719778e-46
+ uc1 = -3.367095838e-10 luc1 = 7.182173155e-17 puc1 = 2.067951531e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.89 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 9.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -3.7585e-8
+ vth0 = {-1.809842643e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.988388349e-07 wvth0 = 9.109733906e-07 pvth0 = -2.324530801e-13
+ k1 = 1.110509677e+00 lk1 = -4.246826391e-08 wk1 = -1.074386706e-06 pk1 = 2.741512558e-13
+ k2 = -2.348795169e+00 lk2 = 5.614290246e-07 wk2 = 2.433087935e-06 pk2 = -6.208510483e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 6.492528619e+00 ldsub = -1.401528528e-06 wdsub = -2.363550562e-07 pdsub = 6.031071970e-14
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {7.676362523e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.326909908e-07 wvoff = -3.607185263e-07 pvoff = 9.204454635e-14
+ nfactor = {3.796926372e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -9.189853320e-06 wnfactor = -2.668008549e-05 pnfactor = 6.807957414e-12
+ eta0 = 2.577143952e+00 leta0 = -5.535732953e-07 weta0 = -5.726959312e-07 peta0 = 1.461348208e-13
+ etab = -4.793348855e-01 letab = 1.223102879e-07 wetab = 5.190928233e-07 petab = -1.324569157e-13
+ u0 = 6.600545432e-02 lu0 = -1.629772176e-08 wu0 = -6.328429781e-08 pu0 = 1.614825427e-14
+ ua = 4.108464464e-08 lua = -1.105726093e-14 wua = -4.040405910e-14 pua = 1.030990376e-20
+ ub = -3.613726974e-17 lub = 9.646356028e-24 wub = 3.443629337e-23 pub = -8.787108978e-30
+ uc = -8.124451085e-11 luc = 1.822275732e-17 wuc = -2.284419859e-18 puc = 5.829154154e-25
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.154102576e+07 lvsat = -8.012293030e+00 wvsat = -2.849779105e+01 pvsat = 7.271781343e-6
+ a0 = 8.593457615e+00 la0 = -1.959161479e-06 wa0 = -7.048401904e-06 pa0 = 1.798540714e-12
+ ags = 1.250000034e+00 lags = -8.762611969e-15 wags = -3.148736027e-14 pags = 8.034632515e-21
+ a1 = 0.0
+ a2 = -6.989463268e+00 la2 = 1.928827674e-06 wa2 = 5.300074792e-06 pa2 = -1.352420085e-12
+ b0 = -1.903053811e-05 lb0 = 4.856022408e-12 wb0 = 1.744951906e-11 pb0 = -4.452593779e-18
+ b1 = 1.742988472e-13 lb1 = -4.447583685e-20 wb1 = -1.598184476e-19 pb1 = 4.078087327e-26
+ keta = -3.829678722e-01 lketa = 8.473401412e-08 wketa = -4.221526723e-08 pketa = 1.077206974e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.139143292e+00 lpclm = -1.162324973e-07 wpclm = 4.936548958e-09 ppclm = -1.259659198e-15
+ pdiblc1 = 2.762203725e+00 lpdiblc1 = -6.031985180e-07 wpdiblc1 = -4.801743096e-07 ppdiblc1 = 1.225260786e-13
+ pdiblc2 = 9.997492380e-02 lpdiblc2 = -2.297466578e-08 wpdiblc2 = -3.366751334e-08 ppdiblc2 = 8.590939378e-15
+ pdiblcb = -1.153807211e-01 lpdiblcb = -4.660672123e-09 wpdiblcb = 1.386200415e-06 ppdiblcb = -3.537167600e-13
+ drout = -3.341571429e+00 ldrout = 9.775916543e-07 wdrout = 4.742114328e-13 pdrout = -1.210045326e-19
+ pscbe1 = 7.999999947e+08 lpscbe1 = 1.353385925e-06 wpscbe1 = 4.863220215e-06 ppscbe1 = -1.240947723e-12
+ pscbe2 = -4.034257020e-08 lpscbe2 = 1.199283754e-14 wpscbe2 = 3.152689577e-14 ppscbe2 = -8.044717992e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 2.133515389e+01 lbeta0 = -3.082164006e-06 wbeta0 = -4.008622653e-06 pbeta0 = 1.022880242e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -5.951120420e-08 lagidl = 1.524280293e-14 wagidl = 5.262797103e-14 pagidl = -1.342907937e-20
+ bgidl = 9.999999962e+08 lbgidl = 9.640083313e-07 wbgidl = 3.464065552e-06 pbgidl = -8.839225769e-13
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -2.8385e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 7.361788721e-01 lkt1 = -3.252291874e-07 wkt1 = -9.767289974e-07 pkt1 = 2.492319383e-13
+ kt2 = 3.567017659e-01 lkt2 = -1.019931754e-07 wkt2 = 6.243217499e-15 pkt2 = -1.593082111e-21
+ at = 9.491710644e+05 lat = -2.291388489e-01 wat = -6.243034395e-01 pat = 1.593035087e-7
+ ute = -3.681908811e+00 lute = 8.763070624e-07 wute = 1.478613298e-06 pute = -3.772977553e-13
+ ua1 = -3.925775991e-09 lua1 = 1.051398893e-15 wua1 = 1.476190227e-22 pua1 = -3.766794559e-29
+ ub1 = 6.680496438e-18 lub1 = -1.610662751e-24 wub1 = -8.109788086e-31 pub1 = 2.069374609e-37
+ uc1 = -1.343328680e-10 luc1 = 2.530772693e-17 wuc1 = -1.036405940e-23 puc1 = 2.644596921e-30
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.90 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 8.6e-07 wmax = 9.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.208394786e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.482947494e-06 wvth0 = 5.033816362e-08 pvth0 = -5.036744533e-12
+ k1 = 3.890552997e-01 lk1 = 4.262509089e-06 wk1 = 3.309711827e-08 pk1 = -3.311637087e-12
+ k2 = 1.182257837e-01 lk2 = -7.188054630e-06 wk2 = -5.581311130e-08 pk2 = 5.584557779e-12
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -2.566011949e-05 lcit = 2.599989202e-09 wcit = 2.018814466e-11 pcit = -2.019988810e-15
+ voff = {-9.714803661e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.014616369e-06 wvoff = -5.446641467e-08 pvoff = 5.449809779e-12
+ nfactor = {1.412570758e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.595912223e-05 wnfactor = 1.239178486e-07 pnfactor = -1.239899316e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 5.412805258e-03 lu0 = 2.859026871e-07 wu0 = 2.219949530e-09 pu0 = -2.221240875e-13
+ ua = -7.852085267e-10 lua = 4.398493784e-15 wua = 3.415299907e-17 pua = -3.417286587e-21
+ ub = -5.364947840e-19 lub = 1.170819404e-22 wub = 9.091065255e-25 pub = -9.096353528e-29
+ uc = -1.966698167e-10 luc = 9.105976534e-15 wuc = 7.070520579e-17 puc = -7.074633501e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.351111826e+05 lvsat = 2.153924035e+01 wvsat = 1.672458100e-01 pvsat = -1.673430969e-5
+ a0 = 2.229227915e+00 la0 = -7.656730485e-05 wa0 = -5.945224025e-07 pa0 = 5.948682362e-11
+ ags = -4.242468240e-01 lags = 5.378495092e-05 wags = 4.176241844e-07 pags = -4.178671164e-11
+ a1 = 0.0
+ a2 = 1.426563877e+00 la2 = -4.568294607e-05 wa2 = -3.547145208e-07 pa2 = 3.549208583e-11
+ b0 = 2.111372840e-08 lb0 = -1.539407793e-12 wb0 = -1.195304473e-14 pb0 = 1.195999782e-18
+ b1 = 1.314825869e-07 lb1 = -9.586431871e-12 wb1 = -7.443579892e-14 pb1 = 7.447909822e-18
+ keta = 9.112462815e-02 lketa = -6.780278710e-06 wketa = -5.264685229e-08 pketa = 5.267747696e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -3.232842371e-01 lpclm = 3.384810171e-05 wpclm = 2.628204661e-07 ppclm = -2.629733488e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 3.849656634e-03 lpdiblc2 = -2.573994256e-07 wpdiblc2 = -1.998630162e-09 ppdiblc2 = 1.999792766e-13
+ pdiblcb = -4.126758726e-01 lpdiblcb = 1.877850437e-05 wpdiblcb = 1.458095143e-07 ppdiblcb = -1.458943317e-11
+ drout = 0.56
+ pscbe1 = 8.001309264e+08 lpscbe1 = -1.310025659e+01 wpscbe1 = -1.017196052e-01 ppscbe1 = 1.017787755e-5
+ pscbe2 = 2.250914045e-08 lpscbe2 = -1.245575675e-12 wpscbe2 = -9.671525522e-15 ppscbe2 = 9.677151448e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -2.685669868e-10 lalpha0 = 2.687232122e-14 walpha0 = 2.086556005e-16 palpha0 = -2.087769755e-20
+ alpha1 = -2.685669868e-10 lalpha1 = 2.687232122e-14 walpha1 = 2.086556005e-16 palpha1 = -2.087769755e-20
+ beta0 = 9.370787793e+01 lbeta0 = -6.374493681e-03 wbeta0 = -4.949605194e-05 pbeta0 = 4.952484379e-9
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 5.808335878e-09 lagidl = -3.910351808e-13 wagidl = -3.036272148e-15 pagidl = 3.038038347e-19
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -2.009458458e+00 legidl = 2.110685530e-04 wegidl = 1.638884684e-06 pegidl = -1.639838023e-10
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.314780834e-01 lkt1 = -6.775855795e-07 wkt1 = -5.261250966e-09 pkt1 = 5.264311436e-13
+ kt2 = -7.516365750e-02 lkt2 = 1.662732400e-06 wkt2 = 1.291062370e-08 pkt2 = -1.291813381e-12
+ at = 2.616457039e+05 lat = -1.907666083e+01 wat = -1.481246108e-01 pat = 1.482107749e-5
+ ute = 4.938624738e-02 lute = -1.324432448e-05 wute = -1.028382496e-07 pute = 1.028980707e-11
+ ua1 = 2.808551428e-09 lua1 = -7.187692928e-14 wua1 = -5.581030280e-16 pua1 = 5.584276765e-20
+ ub1 = -2.606678507e-18 lub1 = 1.378579960e-22 wub1 = 1.070426433e-24 pub1 = -1.071049100e-28
+ uc1 = -8.626253628e-11 luc1 = 5.650638694e-15 wuc1 = 4.387553275e-17 puc1 = -4.390105515e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.91 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 8.6e-07 wmax = 9.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-7.278580422e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.155740195e-06 wvth0 = -3.355877575e-07 pvth0 = 2.704223199e-12
+ k1 = 7.050060672e-01 lk1 = -2.074885116e-06 wk1 = -2.206474552e-07 pk1 = 1.778014704e-12
+ k2 = -4.145757492e-01 lk2 = 3.498969094e-06 wk2 = 3.720874087e-07 pk2 = -2.998343594e-12
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.670593719e-04 lcit = -1.265611119e-09 wcit = -1.345876311e-10 pcit = 1.084530011e-15
+ voff = {-6.170937725e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.414543593e-06 wvoff = 3.631094312e-07 pvoff = -2.925997525e-12
+ nfactor = {2.595511794e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.768510165e-06 wnfactor = -8.261189907e-07 pnfactor = 6.657007267e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.660482421e-02 lu0 = -1.391704317e-07 wu0 = -1.479966354e-08 pu0 = 1.192582047e-13
+ ua = -4.591781400e-10 lua = -2.141079138e-15 wua = -2.276866605e-16 pua = 1.834737817e-21
+ ub = 8.141992028e-18 lub = -5.699262345e-23 wub = -6.060710170e-24 pub = 4.883823287e-29
+ uc = 4.782942044e-10 luc = -4.432566544e-15 wuc = -4.713680386e-16 puc = 3.798363788e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.461446004e+06 lvsat = -1.048477511e+01 wvsat = -1.114972067e+00 pvsat = 8.984634459e-6
+ a0 = -3.446184904e+00 la0 = 3.727109031e-05 wa0 = 3.963482683e-06 pa0 = -3.193841725e-11
+ ags = 3.562465266e+00 lags = -2.618119793e-05 wags = -2.784161229e-06 pags = 2.243524449e-11
+ a1 = 0.0
+ a2 = -1.959601775e+00 la2 = 2.223734023e-05 wa2 = 2.364763472e-06 pa2 = -1.905566607e-11
+ b0 = -9.299208664e-08 lb0 = 7.493460428e-13 wb0 = 7.968696486e-14 pb0 = -6.421311097e-19
+ b1 = -5.790943160e-07 lb1 = 4.666440444e-12 wb1 = 4.962386595e-13 pb1 = -3.998775478e-18
+ keta = -4.114512532e-01 lketa = 3.300473755e-06 wketa = 3.509790153e-07 pketa = -2.828248571e-12
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.185645008e+00 lpclm = -1.647642761e-05 wpclm = -1.752136441e-06 ppclm = 1.411901330e-11
+ pdiblc1 = 0.39
+ pdiblc2 = -1.522960968e-02 lpdiblc2 = 1.252957415e-07 wpdiblc2 = 1.332420108e-08 ppdiblc2 = -1.073686774e-13
+ pdiblcb = 9.792467585e-01 lpdiblcb = -9.140916395e-06 wpdiblcb = -9.720634287e-07 ppdiblcb = 7.833052359e-12
+ drout = 0.56
+ pscbe1 = 7.991598936e+08 lpscbe1 = 6.376884332e+00 wpscbe1 = 6.781307016e-01 ppscbe1 = -5.464492476e-6
+ pscbe2 = -6.981690093e-08 lpscbe2 = 6.063157582e-13 wpscbe2 = 6.447683681e-14 ppscbe2 = -5.195653121e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.723295162e-09 lalpha0 = -1.308078837e-14 walpha0 = -1.391037337e-15 palpha0 = 1.120921533e-20
+ alpha1 = 1.723295162e-09 lalpha1 = -1.308078837e-14 walpha1 = -1.391037337e-15 palpha1 = 1.120921533e-20
+ beta0 = -3.787899229e+02 lbeta0 = 3.102947533e-03 wbeta0 = 3.299736796e-04 pbeta0 = -2.658984006e-9
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.317643879e-08 lagidl = 1.903463569e-13 wagidl = 2.024181432e-14 pagidl = -1.631119809e-19
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 1.363561582e+01 legidl = -1.027430065e-04 wegidl = -1.092589789e-05 pegidl = 8.804274261e-11
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.817028875e-01 lkt1 = 3.298320788e-07 wkt1 = 3.507500644e-08 pkt1 = -2.826403647e-13
+ kt2 = 4.808337066e-02 lkt2 = -8.093774432e-07 wkt2 = -8.607082469e-08 pkt2 = 6.935733374e-13
+ at = -1.152377235e+06 lat = 9.286051666e+00 wat = 9.874974052e-01 pat = -7.957421966e-6
+ ute = -9.323253214e-01 lute = 6.447013055e-06 wute = 6.855883310e-07 pute = -5.524587321e-12
+ ua1 = -2.519195797e-09 lua1 = 3.498793027e-14 wua1 = 3.720686853e-15 pua1 = -2.998192718e-20
+ ub1 = 7.611795810e-18 lub1 = -6.710589894e-23 wub1 = -7.136176220e-24 pub1 = 5.750452113e-29
+ uc1 = 3.325808244e-10 luc1 = -2.750592639e-15 wuc1 = -2.925035517e-16 puc1 = 2.357043345e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.92 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 8.6e-07 wmax = 9.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.119308571e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.365284442e-9
+ k1 = 4.557431136e-01 lk1 = -6.628186177e-8
+ k2 = 1.736465621e-02 lk2 = 1.831987716e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.866729821e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.386030771e-8
+ nfactor = {1.917980732e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.308849687e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 9.209108364e-03 lu0 = 1.007203851e-9
+ ua = -7.714556020e-10 lua = 3.753057380e-16
+ ub = 1.139159733e-18 lub = -5.626103368e-25
+ uc = -7.082993503e-11 luc = -7.630877232e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.687361861e+05 lvsat = -8.737166397e-1
+ a0 = 1.298282802e+00 la0 = -9.606370240e-7
+ ags = 3.007947423e-01 lags = 1.018976364e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.275546727e-04 lketa = -8.401813297e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.415723457e-01 lpclm = -8.107596053e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -1.412456511e-03 lpdiblc2 = 1.395477241e-8
+ pdiblcb = -2.502133320e-01 lpdiblcb = 7.662820228e-7
+ drout = 0.56
+ pscbe1 = 1.230892076e+09 lpscbe1 = -3.472594437e+3
+ pscbe2 = -1.731012336e-08 lpscbe2 = 1.832072184e-13 ppscbe2 = -1.058791184e-34
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.405041024e+00 lbeta0 = 2.315554051e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.940678393e-10 lagidl = -2.006243465e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 1.682321702e+00 legidl = -6.421330460e-6
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.058118873e-01 lkt1 = -2.817105026e-7
+ kt2 = -4.835860979e-02 lkt2 = -3.223156969e-8
+ at = -9.199465573e+04 lat = 7.413085750e-1
+ ute = -1.650014701e-01 lute = 2.637870157e-7
+ ua1 = 5.595420866e-10 lua1 = 1.017893702e-14
+ ub1 = 8.371840607e-19 lub1 = -1.251492578e-23 pub1 = 6.162975822e-45
+ uc1 = -1.167338578e-11 luc1 = 2.346631032e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.93 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 8.6e-07 wmax = 9.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.116324143e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.347660345e-8
+ k1 = 4.428654258e-01 lk1 = -1.402201541e-8
+ k2 = 2.164134381e-02 lk2 = 9.643518320e-10
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.673887289e-01 ldsub = -1.247435718e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.076298863e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.118637217e-8
+ nfactor = {8.205595117e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.144672185e-6
+ eta0 = 1.618122575e-01 leta0 = -3.320080490e-7
+ etab = -1.415226926e-01 letab = 2.902512456e-7
+ u0 = 8.961795572e-03 lu0 = 2.010841203e-9
+ ua = -8.686534836e-10 lua = 7.697512652e-16
+ ub = 1.145979433e-18 lub = -5.902858386e-25
+ uc = -7.565336861e-11 luc = 1.194343622e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 53438.0
+ a0 = 1.058775121e+00 la0 = 1.132585948e-8
+ ags = 1.699111794e-01 lags = 6.330453849e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.740613019e-03 lketa = -3.911472438e-08 pketa = 2.775557562e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.662082328e-01 lpclm = 2.467351305e-06 wpclm = -1.110223025e-22 ppclm = 1.110223025e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 3.668885335e-03 lpdiblc2 = -6.666176630e-9
+ pdiblcb = -9.883598245e-02 lpdiblcb = 1.519670040e-7
+ drout = 0.56
+ pscbe1 = -5.399535418e+07 lpscbe1 = 1.741697186e+3
+ pscbe2 = 4.685632485e-08 lpscbe2 = -7.719113680e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.151404795e+01 lbeta0 = -9.752188105e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.711119258e-10 lagidl = -2.898164661e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.817235263e-01 lkt1 = 2.635183383e-8
+ kt2 = -6.035456581e-02 lkt2 = 1.645005918e-8
+ at = 1.024940121e+05 lat = -4.795950233e-2
+ ute = -1.332981033e-01 lute = 1.351293641e-7
+ ua1 = 3.328055597e-09 lua1 = -1.056161454e-15
+ ub1 = -2.852522339e-18 lub1 = 2.458530043e-24
+ uc1 = 1.859730957e-11 luc1 = -9.937731742e-17 wuc1 = 1.292469707e-32 puc1 = -2.584939414e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.94 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 8.6e-07 wmax = 9.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.127136425e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.776911808e-9
+ k1 = 3.512559901e-01 lk1 = 1.745257769e-7
+ k2 = 5.719390124e-02 lk2 = -7.220885529e-08 pk2 = 5.551115123e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.841659314e-01 ldsub = 1.122659537e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.937752555e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.671186683e-9
+ nfactor = {2.152613232e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.969208211e-07 wnfactor = 3.552713679e-21
+ eta0 = -2.317683150e-01 leta0 = 4.780476779e-07 weta0 = -8.153200337e-23 peta0 = 6.071532166e-29
+ etab = 8.728991787e-01 letab = -1.797601417e-06 wetab = -3.070460552e-22 petab = -8.847089727e-28
+ u0 = 9.740710576e-03 lu0 = 4.077017098e-10
+ ua = -8.760198240e-11 lua = -8.377855030e-16
+ ub = 1.194459582e-19 lub = 1.522494564e-24
+ uc = -7.526918424e-11 luc = 1.115271947e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.984839386e+04 lvsat = -1.319368033e-2
+ a0 = 1.446042456e+00 la0 = -7.857361509e-7
+ ags = 1.631988120e-01 lags = 6.468605781e-7
+ a1 = 0.0
+ a2 = 5.883765817e-01 la2 = 4.355569708e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.074975873e-02 lketa = -3.116565955e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.490103892e-01 lpclm = 3.778587940e-7
+ pdiblc1 = 7.614176700e-01 lpdiblc1 = -7.644407059e-7
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 9.440520000e-02 ldrout = 9.582732495e-7
+ pscbe1 = 7.985241057e+08 lpscbe1 = -1.293279044e+1
+ pscbe2 = 9.536577846e-09 lpscbe2 = -3.807531059e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.831389756e+00 lbeta0 = 1.943688500e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.694326460e-10 lagidl = 8.227161552e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.581851405e-01 lkt1 = -2.209416583e-8
+ kt2 = -5.638602898e-02 lkt2 = 8.282135728e-9
+ at = 9.763617505e+04 lat = -3.796124776e-2
+ ute = 9.699104623e-01 lute = -2.135461409e-06 pute = -6.661338148e-28
+ ua1 = 6.248983323e-09 lua1 = -7.067927273e-15 pua1 = -6.617444900e-36
+ ub1 = -4.359386902e-18 lub1 = 5.559913481e-24 pub1 = 6.162975822e-45
+ uc1 = -1.319123403e-10 luc1 = 2.103971287e-16 wuc1 = -1.033975766e-31 puc1 = -1.033975766e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.95 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 8.6e-07 wmax = 9.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.247665622e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.363172925e-07 wvth0 = 7.230985761e-08 pvth0 = -7.651612203e-14
+ k1 = 4.481980183e-01 lk1 = 7.194463086e-08 wk1 = 5.840886778e-08 pk1 = -6.180651162e-14
+ k2 = -2.453605667e-01 lk2 = 2.479452061e-07 wk2 = 1.783663756e-07 pk2 = -1.887419477e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.970730402e+00 ldsub = -1.263404116e-06 wdsub = -5.312029420e-07 pdsub = 5.621030171e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-6.808742382e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.181047173e-07 wvoff = 3.947971450e-07 pvoff = -4.177624950e-13
+ nfactor = {1.973684900e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.920403158e-05 wnfactor = -1.452544976e-05 pnfactor = 1.537039517e-11
+ eta0 = -4.864342334e-01 leta0 = 7.475275127e-07 weta0 = 3.470726336e-07 peta0 = -3.672618487e-13
+ etab = -1.747468907e+00 letab = 9.751934795e-07 wetab = 2.701294789e-10 petab = -2.858429106e-16
+ u0 = 4.918215320e-02 lu0 = -4.132804963e-08 wu0 = -2.708495895e-08 pu0 = 2.866049101e-14
+ ua = 6.558027621e-09 lua = -7.869991380e-15 wua = -5.499603017e-15 pua = 5.819514925e-21
+ ub = 1.323403901e-18 lub = 2.485023878e-25 wub = 4.617932673e-25 pub = -4.886557817e-31
+ uc = -1.194399028e-10 luc = 5.789284870e-17 wuc = 1.340047268e-17 puc = -1.417997818e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -3.735723379e+06 lvsat = 4.003166503e+00 wvsat = 2.851697252e+00 pvsat = -3.017580481e-6
+ a0 = 1.023395018e+00 la0 = -3.385033115e-07 wa0 = -2.865515246e-07 pa0 = 3.032202268e-13
+ ags = 2.436803294e-01 lags = 5.616974509e-07 wags = 5.487734711e-16 pags = -5.806946035e-22
+ a1 = 0.0
+ a2 = 5.924824229e-01 la2 = 4.312122929e-07 wa2 = 3.586729199e-07 pa2 = -3.795369236e-13
+ b0 = 9.508678650e-16 lb0 = -1.006179849e-21 wb0 = -8.148195926e-22 pb0 = 8.622176483e-28
+ b1 = 3.953193012e-19 lb1 = -4.183150249e-25 wb1 = -3.387578062e-25 pb1 = 3.584633478e-31
+ keta = 8.236469144e-03 lketa = -2.320722270e-08 wketa = 4.187235104e-09 pketa = -4.430806570e-15
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.015045473e+00 lpclm = -1.279272551e-06 wpclm = -2.914860920e-07 ppclm = 3.084418379e-13
+ pdiblc1 = 1.197445943e-01 lpdiblc1 = -8.544150736e-08 wpdiblc1 = -4.240683724e-08 ppdiblc1 = 4.487364296e-14
+ pdiblc2 = 1.507009810e-03 lpdiblc2 = -1.139659471e-09 wpdiblc2 = -5.499626122e-10 ppdiblc2 = 5.819539373e-16
+ pdiblcb = -2.038246775e-01 lpdiblcb = 1.892269089e-07 wpdiblcb = 1.480052940e-07 ppdiblcb = -1.566147620e-13
+ drout = 5.897696755e-01 ldrout = 4.340934225e-07 wdrout = 3.515353902e-07 pdrout = -3.719842038e-13
+ pscbe1 = 2.147777701e+08 lpscbe1 = 6.047700694e+02 wpscbe1 = 4.766484275e+02 ppscbe1 = -5.043750665e-4
+ pscbe2 = 6.687980330e-08 lpscbe2 = -6.105963399e-14 wpscbe2 = -4.959183740e-14 ppscbe2 = 5.247659458e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.198724385e+00 lbeta0 = 1.554986016e-06 wbeta0 = 2.229060778e-07 pbeta0 = -2.358725244e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.227472365e-09 lagidl = 1.836485045e-15 wagidl = 1.789013309e-15 pagidl = -1.893080213e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.676430767e-01 lkt1 = -1.179030615e-07 wkt1 = -3.903428073e-08 pkt1 = 4.130490484e-14
+ kt2 = -8.889678767e-02 lkt2 = 4.268404525e-08 wkt2 = 1.936154988e-08 pkt2 = -2.048781124e-14
+ at = 1.292855489e+05 lat = -7.145166574e-02 wat = -3.234896720e-02 pat = 3.423070663e-8
+ ute = -2.030278943e+00 lute = 1.039249013e-06 wute = 2.884891202e-08 pute = -3.052705323e-14
+ ua1 = -4.533257979e-09 lua1 = 4.341517005e-15 wua1 = 6.489386230e-16 pua1 = -6.866873827e-22
+ ub1 = 5.937735397e-18 lub1 = -5.336192422e-24 wub1 = -1.132462345e-24 pub1 = 1.198337680e-30
+ uc1 = 4.672575110e-10 luc1 = -4.236264329e-16 wuc1 = -9.218760338e-17 puc1 = 9.755015627e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.96 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 8.6e-07 wmax = 9.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-8.908044207e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -6.287192448e-08 wvth0 = -1.611894670e-07 pvth0 = 5.381619598e-14
+ k1 = 1.124209172e+00 lk1 = -3.053845150e-07 wk1 = -5.426247336e-07 pk1 = 2.736724137e-13
+ k2 = 1.418437008e-01 lk2 = 3.181940005e-08 wk2 = -8.547734764e-08 pk2 = -4.147229666e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.009869217e+00 ldsub = 9.584471735e-07 wdsub = 1.364716845e-06 pdsub = -4.961425302e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {8.279012174e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -3.240484789e-07 wvoff = -8.361407187e-07 pvoff = 2.693100925e-13
+ nfactor = {-3.493576818e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.131258315e-05 wnfactor = 2.943420863e-05 pnfactor = -9.166567353e-12
+ eta0 = 1.300044873e+00 leta0 = -2.496315302e-07 weta0 = -6.941452728e-07 peta0 = 2.139147501e-13
+ etab = -1.542022699e-03 letab = 6.694707014e-10 wetab = 1.322247343e-10 petab = -2.088686194e-16
+ u0 = -6.592633025e-02 lu0 = 2.292205258e-08 wu0 = 5.714658411e-08 pu0 = -1.835502938e-14
+ ua = -1.722047064e-08 lua = 5.402452994e-15 wua = 1.186299674e-14 pua = -3.871767382e-21
+ ub = 4.702772645e-18 lub = -1.637759864e-24 wub = -1.609574398e-24 pub = 6.675195083e-31
+ uc = -4.757769023e-11 luc = 1.778151753e-17 wuc = -1.615858291e-17 puc = 2.318999881e-24
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.953115006e+06 lvsat = -3.079362419e+00 wvsat = -6.864246731e+00 pvsat = 2.405567972e-6
+ a0 = 4.567634909e-01 la0 = -2.222659183e-08 wa0 = 3.529035259e-07 pa0 = -5.370439875e-14
+ ags = 6.566598032e-01 lags = 3.311846979e-07 wags = 2.152144425e-07 pags = -1.201262456e-13
+ a1 = 0.0
+ a2 = 2.013906680e+00 la2 = -3.621840847e-07 wa2 = -6.765373739e-07 pa2 = 1.982864061e-13
+ b0 = 1.234351656e-14 lb0 = -7.365214571e-21 wb0 = -1.057743090e-20 pb0 = 6.311414400e-27
+ b1 = -3.828899432e-17 lb1 = 2.117410831e-23 wb1 = 3.281068159e-23 pb1 = -1.814455924e-29
+ keta = -1.459823775e-02 lketa = -1.046157436e-08 wketa = -2.446593746e-08 pketa = 1.156253476e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.421837156e+00 lpclm = 6.390922263e-07 wpclm = 5.971381945e-07 ppclm = -1.875615800e-13
+ pdiblc1 = -6.281934495e-01 lpdiblc1 = 3.320350705e-07 wpdiblc1 = 1.275441663e-07 ppdiblc1 = -4.998790869e-14
+ pdiblc2 = -1.991148667e-02 lpdiblc2 = 1.081550271e-08 wpdiblc2 = 7.428285008e-09 ppdiblc2 = -3.871264537e-15
+ pdiblcb = -2.876384900e-01 lpdiblcb = 2.360092647e-07 wpdiblcb = 4.377978006e-07 ppdiblcb = -3.183682454e-13
+ drout = 2.924526594e+00 ldrout = -8.690978465e-07 wdrout = -1.109463665e-06 pdrout = 4.435016388e-13
+ pscbe1 = 1.912528878e+09 lpscbe1 = -3.428636663e+02 wpscbe1 = -9.533198908e+02 ppscbe1 = 2.937903497e-4
+ pscbe2 = -1.099154682e-07 lpscbe2 = 3.762218270e-14 wpscbe2 = 1.023654995e-13 ppscbe2 = -3.234143218e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.459537072e+00 lbeta0 = 2.930681987e-07 wbeta0 = 3.359715877e-08 pbeta0 = -1.302059650e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 3.263034153e-09 lagidl = -6.699809782e-16 wagidl = -2.533365839e-15 pagidl = 5.195421558e-22
+ bgidl = 4.434916209e+08 lbgidl = 3.106262820e+02 wbgidl = 2.018548977e+02 pbgidl = -1.126693483e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.00081386752815302
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207367379934e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -7.173284075e-01 lkt1 = 7.728079965e-08 wkt1 = 1.317825326e-07 pkt1 = -5.403991586e-14
+ kt2 = 3.960963984e-02 lkt2 = -2.904438739e-08 wkt2 = -4.047100361e-08 pkt2 = 1.290892515e-14
+ at = -1.358929867e+05 lat = 7.656303749e-02 wat = 1.074719794e-01 pat = -4.381315114e-8
+ ute = 1.042737061e+00 lute = -6.760163298e-07 wute = -3.606380872e-07 pute = 1.868729051e-13
+ ua1 = 6.942046448e-09 lua1 = -2.063653667e-15 wua1 = -1.345252456e-15 pua1 = 4.264102517e-22
+ ub1 = -7.817446288e-18 lub1 = 2.341537339e-24 wub1 = 2.217112002e-24 pub1 = -6.712942336e-31
+ uc1 = -4.544898362e-10 luc1 = 9.086528389e-17 wuc1 = 1.252380322e-16 puc1 = -2.381031076e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.97 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 8.6e-07 wmax = 9.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-3.016248679e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.921262325e-07 wvth0 = 1.518451741e-06 pvth0 = -4.637988352e-13
+ k1 = 2.880591799e+00 lk1 = -8.466489491e-07 wk1 = -3.197590255e-06 pk1 = 1.091853138e-12
+ k2 = -1.105556427e+00 lk2 = 4.162306973e-07 wk2 = 1.336442815e-06 pk2 = -4.796654333e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.136633748e+01 ldsub = 6.923529998e-06 wdsub = 1.846474280e-05 pdsub = -5.765857529e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.410178643e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 6.738305918e-07 wvoff = 1.808577362e-06 pvoff = -5.457126784e-13
+ nfactor = {-2.218820869e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.230201496e-06 wnfactor = 1.522660814e-06 pnfactor = -5.650656616e-13
+ eta0 = -5.449783762e+00 leta0 = 1.830463160e-06 weta0 = 5.329844089e-06 peta0 = -1.642498052e-12
+ etab = -9.013276580e-01 letab = 2.779564099e-07 wetab = 7.723621436e-07 petab = -2.381869627e-13
+ u0 = 1.667369527e-01 lu0 = -4.877779134e-08 wu0 = -1.278412258e-07 pu0 = 3.865266399e-14
+ ua = 5.324395453e-08 lua = -1.631256891e-14 wua = -4.098521625e-14 pua = 1.241446642e-20
+ ub = -4.222368766e-17 lub = 1.282356741e-23 wub = 3.146620700e-23 pub = -9.525444045e-30
+ uc = 4.056687881e-10 luc = -1.218954497e-16 wuc = -3.187853634e-16 puc = 9.557949483e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -6.819829584e+06 lvsat = 1.781385916e+00 wvsat = 5.657474775e+00 pvsat = -1.453250945e-6
+ a0 = 5.771857206e+00 la0 = -1.660179022e-06 wa0 = -5.378047953e-06 pa0 = 1.712402918e-12
+ ags = 3.369072419e+00 lags = -5.046994979e-07 wags = -7.686232554e-07 pags = 1.830630177e-13
+ a1 = 0.0
+ a2 = 4.254890783e+00 la2 = -1.052788156e-06 wa2 = -2.288602635e-06 pa2 = 6.950765576e-13
+ b0 = -1.934555114e-06 lb0 = 5.961718459e-13 wb0 = 1.657762837e-12 pb0 = -5.108727705e-19
+ b1 = 1.623342727e-13 lb1 = -5.001717824e-20 wb1 = -1.391078097e-19 pb1 = 4.286082041e-26
+ keta = 1.666884925e+00 lketa = -5.286442407e-07 wketa = -1.405659213e-06 pketa = 4.372048665e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.489653964e+00 lpclm = 6.599913319e-07 wpclm = 1.692380531e-06 ppclm = -5.250824108e-13
+ pdiblc1 = -6.995892739e+00 lpdiblc1 = 2.294368961e-06 wpdiblc1 = 6.375853807e-06 ppdiblc1 = -1.975529491e-12
+ pdiblc2 = -1.678382620e-01 lpdiblc2 = 5.640209707e-08 wpdiblc2 = 1.495307479e-07 ppdiblc2 = -4.766298053e-14
+ pdiblcb = -5.569933789e+00 lpdiblcb = 1.863854207e-06 wpdiblcb = 4.345951682e-06 ppdiblcb = -1.522744027e-12
+ drout = 1.565973586e+01 ldrout = -4.793707285e-06 wdrout = -1.300154399e-05 pdrout = 4.108284032e-12
+ pscbe1 = 7.997765439e+08 lpscbe1 = 5.322040342e-02 wpscbe1 = 8.226946134e-02 ppscbe1 = -1.959400463e-8
+ pscbe2 = 5.475163447e-08 lpscbe2 = -1.312327832e-14 wpscbe2 = -3.178948879e-14 ppscbe2 = 9.001110573e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -1.996281420e+01 lbeta0 = 9.051984191e-06 wbeta0 = 2.390820550e-05 pbeta0 = -7.487644017e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 4.182598126e-09 lagidl = -9.533630079e-16 wagidl = -3.861956906e-15 pagidl = 9.289740651e-22
+ bgidl = 2.987531367e+09 lbgidl = -4.733704466e+02 wbgidl = -7.209115844e+02 pbgidl = 1.716995985e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.00081386752815302
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207367379934e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.524560080e-01 lkt1 = -9.679592770e-08 wkt1 = -2.515803420e-07 pkt1 = 6.410102121e-14
+ kt2 = -1.853879540e+00 lkt2 = 5.544721731e-07 wkt2 = 1.514133684e-06 pkt2 = -4.661736014e-13
+ at = -6.673738997e+03 lat = 3.674154193e-02 wat = 1.283192874e-01 pat = -5.023766603e-8
+ ute = 2.308535144e+00 lute = -1.066097325e-06 wute = -4.515959981e-06 pute = 1.467418453e-12
+ ua1 = 1.855843567e-08 lua1 = -5.643476333e-15 wua1 = -1.537492687e-14 pua1 = 4.749935017e-21
+ ub1 = -3.000691454e-17 lub1 = 9.179665769e-24 wub1 = 2.398317585e-23 pub1 = -7.378942130e-30
+ uc1 = -1.465508807e-10 luc1 = -4.032264020e-18 wuc1 = -1.629511762e-16 puc1 = 6.500095759e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.98 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 8.6e-07 wmax = 9.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -3.7585e-8
+ vth0 = {2.683109888e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -8.199145511e-07 wvth0 = -2.939136478e-06 pvth0 = 6.405391089e-13
+ k1 = -1.266881946e+01 lk1 = 3.060662562e-06 wk1 = 1.073342358e-05 pk1 = -2.384989818e-12
+ k2 = 6.333017879e+00 lk2 = -1.452160765e-06 wk2 = -5.006548666e-06 pk2 = 1.104638342e-12
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 6.350585798e+01 ldsub = -1.423912325e-05 wdsub = -4.909233128e-05 pdsub = 1.106112806e-11
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {5.558802475e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.311517918e-06 wvoff = -4.466374268e-06 pvoff = 1.016515075e-12
+ nfactor = {4.640493227e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.108931278e-05 wnfactor = -3.390879545e-05 pnfactor = 8.435646011e-12
+ eta0 = 1.812578947e+01 leta0 = -4.054661816e-06 weta0 = -1.389667234e-05 peta0 = 3.146294598e-12
+ etab = 1.787942674e+00 letab = -3.884248427e-07 wetab = -1.423787198e-06 petab = 3.052032539e-13
+ u0 = -2.359718134e-01 lu0 = 5.049976344e-08 wu0 = 1.954866664e-07 pu0 = -4.109198034e-14
+ ua = -6.948096770e-08 lua = 1.383879768e-14 wua = 5.434204655e-14 pua = -1.102407657e-20
+ ub = 4.851141506e-17 lub = -9.413993450e-24 wub = -3.810102691e-23 pub = 7.546123817e-30
+ uc = -9.003804298e-10 luc = 2.026685261e-16 wuc = 6.996511701e-16 puc = -1.574727217e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.951694611e+06 lvsat = -3.296928845e-01 wvsat = -3.142042224e+00 pvsat = 6.883922614e-7
+ a0 = -9.390038959e+00 la0 = 2.090182449e-06 wa0 = 8.362051947e-06 pa0 = -1.671431184e-12
+ ags = 1.249999290e+00 lags = 1.599978567e-13 wags = 6.065636029e-13 pags = -1.365799278e-19
+ a1 = 0.0
+ a2 = -1.316854408e+01 la2 = 3.318004240e-06 wa2 = 1.059506508e-05 pa2 = -2.542836046e-12
+ b0 = 6.388770759e-06 lb0 = -1.485137909e-12 wb0 = -4.332845930e-12 pb0 = 9.812860027e-19
+ b1 = -2.311818848e-13 lb1 = 4.682623416e-20 wb1 = 1.876469122e-19 pb1 = -3.745788002e-26
+ keta = -4.651323511e+00 lketa = 1.045839656e-06 wketa = 3.615432584e-06 pketa = -8.128204987e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.223951270e+00 lpclm = -1.261180727e-06 wpclm = -4.352347274e-06 ppclm = 9.798716674e-13
+ pdiblc1 = 2.180100999e+01 lpdiblc1 = -4.889970188e-06 wpdiblc1 = -1.679494625e-05 ppdiblc1 = 3.795955031e-12
+ pdiblc2 = 6.016733293e-01 lpdiblc2 = -1.359283301e-07 wpdiblc2 = -4.635839144e-07 ppdiblc2 = 1.053834193e-13
+ pdiblcb = 2.022731196e+01 lpdiblcb = -4.585791575e-06 wpdiblcb = -1.604590048e-05 ppdiblcb = 3.571955095e-12
+ drout = -4.550485825e+01 ldrout = 1.047149893e-05 wdrout = 3.613064855e-05 pdrout = -8.135538134e-12
+ pscbe1 = 7.999999957e+08 lpscbe1 = 9.653663635e-07 wpscbe1 = 4.034484863e-06 ppscbe1 = -9.084453583e-13
+ pscbe2 = -9.950073780e-08 lpscbe2 = 2.530059156e-14 wpscbe2 = 8.222083106e-14 ppscbe2 = -1.944842519e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.602233588e+01 lbeta0 = -1.989783776e-05 wbeta0 = -6.800971202e-05 pbeta0 = 1.543260103e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.491828662e-09 lagidl = -3.348081153e-16 wagidl = 3.531301069e-16 pagidl = -8.028176051e-23
+ bgidl = 9.999963961e+08 lbgidl = 8.114767914e-04 wbgidl = 3.088467194e-03 pbgidl = -6.954301548e-10
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -2.8385e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 5.656543700e-01 lkt1 = -2.869452126e-07 wkt1 = -8.306027999e-07 pkt1 = 2.164255580e-13
+ kt2 = 4.755641863e+00 lkt2 = -1.092502517e-06 wkt2 = -3.769548540e-06 pkt2 = 8.487892447e-13
+ at = 1.760662207e+06 lat = -4.116070489e-01 wat = -1.319688053e+00 pat = 3.156645235e-7
+ ute = -1.999236540e+01 lute = 4.548328013e-06 wute = 1.545540238e-05 pute = -3.523933292e-12
+ ua1 = -4.927233127e-08 lua1 = 1.126208274e-14 wua1 = 3.885846099e-14 pua1 = -8.749759662e-21
+ ub1 = 7.614797079e-17 lub1 = -1.725265392e-23 wub1 = -5.952820787e-23 pub1 = 1.340396657e-29
+ uc1 = -1.225848697e-09 luc1 = 2.710843464e-16 wuc1 = 9.353439166e-16 puc1 = -2.106113897e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.99 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 8.4e-07 wmax = 8.6e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.143603+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43165561
+ k2 = 0.046387026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
+ voff = {-0.16725342+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.5720692+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.00827017
+ ua = -7.4124916e-10
+ ub = 6.3364395e-19
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = 5.7286e-9
+ b1 = 3.5674e-8
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.100 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 8.4e-07 wmax = 8.6e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.159803279e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.249479557e-7
+ k1 = 4.210039986e-01 lk1 = 2.136518329e-7
+ k2 = 6.434930204e-02 lk2 = -3.602903863e-7
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.172472591e-06 lcit = 1.303205335e-10 wcit = -1.355252716e-26 pcit = 8.131516294e-32
+ voff = {-1.497245500e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -3.515970554e-7
+ nfactor = {1.532188847e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.999269080e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 7.555725933e-03 lu0 = 1.433044056e-8
+ ua = -7.522405845e-10 lua = 2.204678604e-16
+ ub = 3.410671347e-19 lub = 5.868555500e-24
+ uc = -1.284179734e-10 luc = 4.564233263e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.633145348e+04 lvsat = 1.079621904e+0
+ a0 = 1.655334532e+00 la0 = -3.837820560e-6
+ ags = -2.111356046e-02 lags = 2.695889464e-6
+ a1 = 0.0
+ a2 = 1.084157408e+00 la2 = -2.289788703e-6
+ b0 = 9.575436055e-09 lb0 = -7.716049156e-14
+ b1 = 5.962959638e-08 lb1 = -4.805054247e-13
+ keta = 4.030454116e-02 lketa = -3.398512340e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.958323949e-02 lpclm = 1.696584997e-06 ppclm = -3.552713679e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 1.920375883e-03 lpdiblc2 = -1.290175761e-8
+ pdiblcb = -2.719257256e-01 lpdiblcb = 9.412441810e-7
+ drout = 0.56
+ pscbe1 = 8.000327363e+08 lpscbe1 = -6.566305840e-1
+ pscbe2 = 1.317320208e-08 lpscbe2 = -6.243260025e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.715141667e-11 lalpha0 = 1.346934531e-15
+ alpha1 = -6.715141667e-11 lalpha1 = 1.346934531e-15
+ beta0 = 4.592926334e+01 lbeta0 = -3.195118720e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.877417733e-09 lagidl = -1.960004808e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -4.274405672e-01 legidl = 1.057949256e-05 wegidl = -8.881784197e-22 pegidl = 2.842170943e-26
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.365567770e-01 lkt1 = -3.396295421e-8
+ kt2 = -6.270101271e-02 lkt2 = 8.334195126e-8
+ at = 1.186607907e+05 lat = -9.561888237e-1
+ ute = -4.988367220e-02 lute = -6.638517694e-7
+ ua1 = 2.269813722e-09 lua1 = -3.602722566e-15
+ ub1 = -1.573394235e-18 lub1 = 6.909923924e-24
+ uc1 = -4.390941745e-11 luc1 = 2.832297336e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.101 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 8.4e-07 wmax = 8.6e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.119308571e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.365284442e-9
+ k1 = 4.557431136e-01 lk1 = -6.628186177e-8
+ k2 = 1.736465621e-02 lk2 = 1.831987716e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.866729821e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.386030771e-8
+ nfactor = {1.917980732e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.308849687e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 9.209108364e-03 lu0 = 1.007203851e-9
+ ua = -7.714556020e-10 lua = 3.753057380e-16
+ ub = 1.139159733e-18 lub = -5.626103368e-25
+ uc = -7.082993503e-11 luc = -7.630877232e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.687361861e+05 lvsat = -8.737166397e-1
+ a0 = 1.298282802e+00 la0 = -9.606370240e-7
+ ags = 3.007947423e-01 lags = 1.018976364e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.275546728e-04 lketa = -8.401813297e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.415723457e-01 lpclm = -8.107596053e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -1.412456511e-03 lpdiblc2 = 1.395477241e-08 wpdiblc2 = 3.469446952e-24 ppdiblc2 = 2.775557562e-29
+ pdiblcb = -2.502133320e-01 lpdiblcb = 7.662820228e-7
+ drout = 0.56
+ pscbe1 = 1.230892076e+09 lpscbe1 = -3.472594437e+3
+ pscbe2 = -1.731012336e-08 lpscbe2 = 1.832072184e-13 ppscbe2 = 2.117582368e-34
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.405041024e+00 lbeta0 = 2.315554051e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.940678393e-10 lagidl = -2.006243465e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 1.682321702e+00 legidl = -6.421330460e-6
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.058118873e-01 lkt1 = -2.817105026e-7
+ kt2 = -4.835860979e-02 lkt2 = -3.223156969e-8
+ at = -9.199465573e+04 lat = 7.413085750e-1
+ ute = -1.650014701e-01 lute = 2.637870157e-7
+ ua1 = 5.595420866e-10 lua1 = 1.017893702e-14
+ ub1 = 8.371840607e-19 lub1 = -1.251492578e-23 pub1 = -2.465190329e-44
+ uc1 = -1.167338578e-11 luc1 = 2.346631032e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.102 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 8.4e-07 wmax = 8.6e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.116324143e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.347660345e-8
+ k1 = 4.428654258e-01 lk1 = -1.402201541e-8
+ k2 = 2.164134381e-02 lk2 = 9.643518320e-10
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.673887289e-01 ldsub = -1.247435718e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.076298863e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.118637217e-8
+ nfactor = {8.205595117e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.144672185e-6
+ eta0 = 1.618122575e-01 leta0 = -3.320080490e-7
+ etab = -1.415226926e-01 letab = 2.902512456e-7
+ u0 = 8.961795572e-03 lu0 = 2.010841203e-9
+ ua = -8.686534836e-10 lua = 7.697512652e-16
+ ub = 1.145979433e-18 lub = -5.902858386e-25
+ uc = -7.565336861e-11 luc = 1.194343622e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 53438.0
+ a0 = 1.058775121e+00 la0 = 1.132585948e-8
+ ags = 1.699111794e-01 lags = 6.330453849e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.740613019e-03 lketa = -3.911472438e-08 pketa = 5.551115123e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.662082328e-01 lpclm = 2.467351305e-06 wpclm = 1.332267630e-21 ppclm = 8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 3.668885335e-03 lpdiblc2 = -6.666176630e-09 wpdiblc2 = 1.387778781e-23
+ pdiblcb = -9.883598245e-02 lpdiblcb = 1.519670040e-7
+ drout = 0.56
+ pscbe1 = -5.399535418e+07 lpscbe1 = 1.741697186e+3
+ pscbe2 = 4.685632485e-08 lpscbe2 = -7.719113680e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.151404795e+01 lbeta0 = -9.752188105e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.711119258e-10 lagidl = -2.898164661e-16 wagidl = 1.654361225e-30
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.817235264e-01 lkt1 = 2.635183383e-8
+ kt2 = -6.035456581e-02 lkt2 = 1.645005918e-8
+ at = 1.024940121e+05 lat = -4.795950233e-2
+ ute = -1.332981033e-01 lute = 1.351293641e-7
+ ua1 = 3.328055596e-09 lua1 = -1.056161454e-15
+ ub1 = -2.852522339e-18 lub1 = 2.458530043e-24
+ uc1 = 1.859730957e-11 luc1 = -9.937731742e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.103 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 8.4e-07 wmax = 8.6e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.127136425e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.776911808e-9
+ k1 = 3.512559901e-01 lk1 = 1.745257769e-7
+ k2 = 5.719390124e-02 lk2 = -7.220885529e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.841659314e-01 ldsub = 1.122659537e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.937752555e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.671186683e-9
+ nfactor = {2.152613232e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.969208211e-7
+ eta0 = -2.317683150e-01 leta0 = 4.780476779e-07 weta0 = 1.873501354e-22 peta0 = 5.065392550e-28
+ etab = 8.728991787e-01 letab = -1.797601417e-06 wetab = 1.231653668e-21 petab = 2.567390744e-27
+ u0 = 9.740710576e-03 lu0 = 4.077017098e-10
+ ua = -8.760198240e-11 lua = -8.377855030e-16
+ ub = 1.194459582e-19 lub = 1.522494564e-24
+ uc = -7.526918424e-11 luc = 1.115271947e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.984839386e+04 lvsat = -1.319368033e-2
+ a0 = 1.446042456e+00 la0 = -7.857361509e-7
+ ags = 1.631988120e-01 lags = 6.468605781e-7
+ a1 = 0.0
+ a2 = 5.883765817e-01 la2 = 4.355569708e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.074975873e-02 lketa = -3.116565955e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.490103892e-01 lpclm = 3.778587940e-7
+ pdiblc1 = 7.614176700e-01 lpdiblc1 = -7.644407059e-7
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 9.440520000e-02 ldrout = 9.582732495e-7
+ pscbe1 = 7.985241057e+08 lpscbe1 = -1.293279044e+1
+ pscbe2 = 9.536577846e-09 lpscbe2 = -3.807531059e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.831389756e+00 lbeta0 = 1.943688500e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.694326460e-10 lagidl = 8.227161552e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.581851405e-01 lkt1 = -2.209416583e-8
+ kt2 = -5.638602898e-02 lkt2 = 8.282135728e-9
+ at = 9.763617505e+04 lat = -3.796124776e-2
+ ute = 9.699104623e-01 lute = -2.135461409e-06 pute = 2.664535259e-27
+ ua1 = 6.248983323e-09 lua1 = -7.067927273e-15
+ ub1 = -4.359386902e-18 lub1 = 5.559913481e-24 wub1 = -1.232595164e-38 pub1 = 1.232595164e-44
+ uc1 = -1.319123403e-10 luc1 = 2.103971287e-16 wuc1 = -2.067951531e-31 puc1 = -4.135903063e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.104 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 8.4e-07 wmax = 8.6e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.154593399e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.783105829e-8
+ k1 = 5.233778534e-01 lk1 = -7.608415156e-9
+ k2 = -1.577976505e-02 lk2 = 5.009689160e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.287002896e+00 ldsub = -5.399041805e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.727187927e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.961013053e-8
+ nfactor = {1.040699630e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.796727960e-7
+ eta0 = -3.970646192e-02 leta0 = 2.748135868e-7
+ etab = -1.747121215e+00 letab = 9.748255624e-7
+ u0 = 1.432027652e-02 lu0 = -4.438257587e-9
+ ua = -5.206791442e-10 lua = -3.795162426e-16
+ ub = 1.917792099e-18 lub = -3.804613713e-25
+ uc = -1.021917457e-10 luc = 3.964136635e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -6.521687765e+04 lvsat = 1.191466380e-01 pvsat = 2.328306437e-22
+ a0 = 6.545658119e-01 la0 = 5.178068979e-8
+ ags = 2.436803301e-01 lags = 5.616974501e-7
+ a1 = 0.0
+ a2 = 1.054141277e+00 la2 = -5.730125626e-8
+ b0 = -9.791128221e-17 lb0 = 1.036067815e-22
+ b1 = -4.070620229e-20 lb1 = 4.307408208e-26
+ keta = 1.362598715e-02 lketa = -2.891024897e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.639864835e+00 lpclm = -8.822676549e-7
+ pdiblc1 = 6.516146082e-02 lpdiblc1 = -2.768327299e-8
+ pdiblc2 = 7.991361598e-04 lpdiblc2 = -3.906088102e-10
+ pdiblcb = -1.332254979e-02 lpdiblcb = -1.235672748e-8
+ drout = 1.042241597e+00 ldrout = -4.469879061e-8
+ pscbe1 = 8.282864975e+08 lpscbe1 = -4.442646058e+1
+ pscbe2 = 3.048636988e-09 lpscbe2 = 6.484591271e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.485633595e+00 lbeta0 = 1.251387297e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.075221224e-09 lagidl = -6.001562308e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.178852899e-01 lkt1 = -6.473825875e-8
+ kt2 = -6.397594635e-02 lkt2 = 1.631355860e-8
+ at = 8.764820671e+04 lat = -2.739227930e-2
+ ute = -1.993146628e+00 lute = 9.999567120e-7
+ ua1 = -3.697989286e-09 lua1 = 3.457660733e-15 pua1 = -6.617444900e-36
+ ub1 = 4.480108576e-18 lub1 = -3.793775449e-24
+ uc1 = 3.486000352e-10 luc1 = -2.980666517e-16 puc1 = 4.135903063e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.105 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 8.4e-07 wmax = 8.6e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.098276299e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.396542597e-9
+ k1 = 4.257803294e-01 lk1 = 4.686759479e-8
+ k2 = 3.182319986e-02 lk2 = -2.156085776e-08 wk2 = 5.551115123e-23 pk2 = -2.775557562e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.533005469e-01 ldsub = 3.198469920e-07 pdsub = 8.881784197e-28
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.483210014e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.258875430e-8
+ nfactor = {2.949899408e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.859852442e-7
+ eta0 = 4.065893232e-01 leta0 = 2.570466844e-8
+ etab = -1.371832211e-03 letab = 4.006295315e-10
+ u0 = 7.628780961e-03 lu0 = -7.032655101e-10
+ ua = -1.951245750e-09 lua = 4.189831196e-16
+ ub = 2.631040349e-18 lub = -7.785751474e-25
+ uc = -6.837589508e-11 luc = 2.076637300e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.179337001e+05 lvsat = 1.691748002e-2
+ a0 = 9.109963816e-01 la0 = -9.135116129e-8
+ ags = 9.336688756e-01 lags = 1.765665437e-7
+ a1 = 0.0
+ a2 = 1.143114794e+00 la2 = -1.069636043e-7
+ b0 = -1.271017328e-15 lb0 = 7.583993833e-22 wb0 = 1.577721810e-36
+ b1 = 3.942634583e-18 lb1 = -2.180307244e-24 wb1 = 1.194076566e-38 pb1 = 2.792598419e-45
+ keta = -4.608909199e-02 lketa = 4.420916754e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.532423753e-01 lpclm = 3.976759966e-07 wpclm = 8.881784197e-22 ppclm = 8.881784197e-28
+ pdiblc1 = -4.640274633e-01 lpdiblc1 = 2.676941088e-07 wpdiblc1 = -8.881784197e-22 ppdiblc1 = -3.885780586e-28
+ pdiblc2 = -1.035031450e-02 lpdiblc2 = 5.832680064e-09 wpdiblc2 = 2.688821388e-23 ppdiblc2 = 6.071532166e-30
+ pdiblcb = 2.758644106e-01 lpdiblcb = -1.737722132e-07 ppdiblcb = -4.440892099e-28
+ drout = 1.496502075e+00 ldrout = -2.982533618e-7
+ pscbe1 = 6.854817729e+08 lpscbe1 = 3.528285254e+1
+ pscbe2 = 2.184228811e-08 lpscbe2 = -4.005460978e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.502780999e+00 lbeta0 = 1.254761302e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.261721264e-12 lagidl = -1.262424958e-18
+ bgidl = 7.033052157e+08 lbgidl = 1.656061277e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.00081386752815302
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207367379934e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.477070908e-01 lkt1 = 7.724375894e-9
+ kt2 = -1.248182315e-02 lkt2 = -1.242891616e-8
+ at = 2.437475586e+03 lat = 2.016979449e-2
+ ute = 5.785487810e-01 lute = -4.354865146e-07 pute = 8.881784197e-28
+ ua1 = 5.210530986e-09 lua1 = -1.514808027e-15
+ ub1 = -4.963733815e-18 lub1 = 1.477494058e-24
+ uc1 = -2.932921455e-10 luc1 = 6.021830677e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.106 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 8.4e-07 wmax = 8.6e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.061803134e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.843392784e-9
+ k1 = -1.235124135e+00 lk1 = 5.587085235e-7
+ k2 = 6.146198786e-01 lk2 = -2.011613102e-07 wk2 = 1.776356839e-21 pk2 = -2.220446049e-28
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.400196095e+00 ldsub = -4.978810681e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-8.230356455e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.857283922e-8
+ nfactor = {-2.589576988e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.028882504e-7
+ eta0 = 1.410421109e+00 leta0 = -2.836461730e-7
+ etab = 9.280321174e-02 letab = -2.862129376e-08 wetab = -1.890848589e-22 petab = 5.637851297e-30
+ u0 = 2.188612260e-03 lu0 = 9.732312786e-10
+ ua = 4.906327663e-10 lua = -3.335305827e-16
+ ub = -1.722573007e-18 lub = 5.630778806e-25 pub = 7.703719778e-46
+ uc = -4.649575163e-12 luc = 1.127832989e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.620787347e+05 lvsat = -8.913769527e-2
+ a0 = -1.150392329e+00 la0 = 5.439069975e-7
+ ags = 2.379753986e+00 lags = -2.690735049e-7
+ a1 = 0.0
+ a2 = 1.309160536e+00 la2 = -1.581339208e-7
+ b0 = 1.992019908e-07 lb0 = -6.138807714e-14 wb0 = -5.323208145e-29 pb0 = 7.629039736e-35
+ b1 = -1.671563145e-14 lb1 = 5.150290839e-21 wb1 = -3.328006944e-35 pb1 = -1.182058763e-41
+ keta = -1.423819160e-01 lketa = 3.409547632e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.886606297e-01 lpclm = -1.585825243e-8
+ pdiblc1 = 1.210663141e+00 lpdiblc1 = -2.483952947e-7
+ pdiblc2 = 2.462732385e-02 lpdiblc2 = -4.946378746e-9
+ pdiblcb = 2.387315920e-02 lpdiblcb = -9.611606923e-8
+ drout = -1.074947920e+00 ldrout = 4.941903832e-7
+ pscbe1 = 7.998824354e+08 lpscbe1 = 2.800036250e-2
+ pscbe2 = 1.383441396e-08 lpscbe2 = -1.537674398e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.081016622e+01 lbeta0 = -5.855907746e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -7.882443863e-10 lagidl = 2.423478422e-16 wagidl = 7.237830360e-31 pagidl = -4.006656092e-37
+ bgidl = 2.059624081e+09 lbgidl = -2.523706570e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.00081386752815302
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207367379934e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.762727387e-01 lkt1 = -1.428954841e-8
+ kt2 = 9.500810120e-02 lkt2 = -4.555408614e-8
+ at = 1.584899291e+05 lat = -2.792089011e-2
+ ute = -3.504094670e+00 lute = 8.226617178e-7
+ ua1 = -1.231101597e-09 lua1 = 4.703098857e-16
+ ub1 = 8.625625182e-19 lub1 = -3.179956828e-25
+ uc1 = -3.562903090e-10 luc1 = 7.963245083e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.107 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 8.4e-07 wmax = 8.6e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -3.7585e-8
+ vth0 = {-1.773728647e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.764729308e-07 wvth0 = 5.234794304e-07 pvth0 = -1.335762463e-13
+ k1 = 2.500725974e+00 lk1 = -3.546890823e-07 wk1 = -1.052130001e-06 pk1 = 2.684720124e-13
+ k2 = 4.389924596e+00 lk2 = -1.178864224e-06 wk2 = -3.496916746e-06 pk2 = 8.923082462e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 6.155372620e-01 ldsub = -7.802722317e-08 wdsub = -2.314575264e-07 pdsub = 5.906101702e-14
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {2.742883855e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.216038674e-07 wvoff = -3.607190127e-07 pvoff = 9.204467048e-14
+ nfactor = {3.710063192e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -8.994263282e-06 wnfactor = -2.668007982e-05 pnfactor = 6.807955967e-12
+ eta0 = 9.760944361e-01 leta0 = -1.930650154e-07 weta0 = -5.726969806e-07 peta0 = 1.461350885e-13
+ etab = -6.989563216e-01 letab = 1.713690675e-07 wetab = 5.083393439e-07 petab = -1.297129504e-13
+ u0 = 3.702679942e-01 lu0 = -9.288011772e-08 wu0 = -2.755143774e-07 pu0 = 7.030300369e-14
+ ua = 5.246991730e-08 lua = -1.362089123e-14 wua = -4.040427892e-14 pua = 1.030995985e-20
+ ub = -4.485452068e-17 lub = 1.160924811e-23 wub = 3.443702262e-23 pub = -8.787295062e-30
+ uc = 3.041376388e-12 luc = -7.541651208e-19 wuc = -2.237106428e-18 puc = 5.708424473e-25
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -8.460994898e+07 lvsat = 2.161232918e+01 wvsat = 6.410960304e+01 pvsat = -1.635884741e-5
+ a0 = 1.044522570e+01 la0 = -2.376124087e-06 wa0 = -7.048401546e-06 pa0 = 1.798540622e-12
+ ags = 1.249999979e+00 lags = 7.421803616e-15 wags = 7.069888852e-14 pags = -1.804023952e-20
+ a1 = 0.0
+ a2 = -6.211877916e+00 la2 = 1.749722243e-06 wa2 = 5.190278091e-06 pa2 = -1.324403261e-12
+ b0 = 3.375230690e-05 lb0 = -8.627515589e-12 wb0 = -2.559217915e-11 pb0 = 6.530356355e-18
+ b1 = 2.160520618e-13 lb1 = -5.387742611e-20 wb1 = -1.598189800e-19 pb1 = 4.078100913e-26
+ keta = 5.654630095e-02 lketa = -1.423138395e-08 wketa = -4.221504654e-08 pketa = 1.077201343e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.156898003e-01 lpclm = 1.629790326e-09 wpclm = 4.834443994e-09 ppclm = -1.233605074e-15
+ pdiblc1 = 7.889652504e-01 lpdiblc1 = -1.585205008e-07 wpdiblc1 = -4.702264283e-07 ppdiblc1 = 1.199876777e-13
+ pdiblc2 = 4.741710782e-02 lpdiblc2 = -1.111470850e-08 wpdiblc2 = -3.297006227e-08 ppdiblc2 = 8.412970790e-15
+ pdiblcb = -2.173113372e+00 lpdiblcb = 4.576284509e-07 wpdiblcb = 1.357482767e-06 ppdiblcb = -3.463888778e-13
+ drout = 1.000002905e+00 ldrout = -7.015411541e-13 wdrout = -1.195128249e-12 pdrout = 3.049608779e-19
+ pscbe1 = 8.000000149e+08 lpscbe1 = -3.790267944e-06 wpscbe1 = -1.091946411e-05 ppscbe1 = 2.786315918e-12
+ pscbe2 = -3.341037846e-08 lpscbe2 = 1.040802379e-14 wpscbe2 = 3.087377690e-14 ppscbe2 = -7.878061651e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.353769600e+01 lbeta0 = -1.323372603e-06 wbeta0 = -3.925580628e-06 pbeta0 = 1.001690409e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.693023107e-08 lagidl = -1.702007734e-14 wagidl = -5.048740437e-14 pagidl = 1.288287097e-20
+ bgidl = 1.000000381e+09 lbgidl = -8.618704224e-05 wbgidl = -7.777648926e-06 pbgidl = 1.984626770e-12
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -2.8385e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 7.390551914e-01 lkt1 = -3.254247298e-07 wkt1 = -9.653217130e-07 pkt1 = 2.463211415e-13
+ kt2 = -9.625899412e-02 lkt2 = -2.194799897e-15 wkt2 = -2.199544014e-14 pkt2 = 5.612577070e-21
+ at = 8.489649324e+05 lat = -2.061023225e-01 wat = -6.113703824e-01 pat = 1.560033805e-7
+ ute = -1.962988343e+00 lute = 4.881372249e-07 wute = 1.447982697e-06 pute = -3.694817449e-13
+ ua1 = 7.435795145e-10 lua1 = 9.157036950e-23 wua1 = -4.480532446e-22 pua1 = 1.143297477e-28
+ ub1 = -4.726034449e-19 lub1 = 8.513161447e-31 wub1 = 1.908134943e-30 pub1 = -4.868987897e-37
+ uc1 = -2.193904752e-11 luc1 = 1.165633720e-23 wuc1 = 2.411704716e-23 puc1 = -6.153947065e-30
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.108 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 8.2e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.143603+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43165561
+ k2 = 0.046387026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
+ voff = {-0.16725342+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.5720692+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.00827017
+ ua = -7.4124916e-10
+ ub = 6.3364395e-19
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = 5.7286e-9
+ b1 = 3.5674e-8
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.109 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 8.2e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.159803279e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.249479557e-7
+ k1 = 4.210039986e-01 lk1 = 2.136518329e-7
+ k2 = 6.434930204e-02 lk2 = -3.602903863e-7
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.172472591e-06 lcit = 1.303205335e-10 wcit = -3.388131789e-27 pcit = 1.355252716e-31
+ voff = {-1.497245500e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -3.515970554e-07 wvoff = -8.881784197e-22
+ nfactor = {1.532188847e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.999269080e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 7.555725933e-03 lu0 = 1.433044056e-8
+ ua = -7.522405845e-10 lua = 2.204678604e-16
+ ub = 3.410671347e-19 lub = 5.868555500e-24
+ uc = -1.284179734e-10 luc = 4.564233263e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.633145348e+04 lvsat = 1.079621904e+0
+ a0 = 1.655334532e+00 la0 = -3.837820560e-6
+ ags = -2.111356046e-02 lags = 2.695889464e-06 pags = -7.105427358e-27
+ a1 = 0.0
+ a2 = 1.084157408e+00 la2 = -2.289788703e-6
+ b0 = 9.575436055e-09 lb0 = -7.716049156e-14
+ b1 = 5.962959638e-08 lb1 = -4.805054247e-13
+ keta = 4.030454116e-02 lketa = -3.398512340e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.958323949e-02 lpclm = 1.696584997e-06 ppclm = 1.776356839e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 1.920375883e-03 lpdiblc2 = -1.290175761e-8
+ pdiblcb = -2.719257256e-01 lpdiblcb = 9.412441810e-7
+ drout = 0.56
+ pscbe1 = 8.000327363e+08 lpscbe1 = -6.566305839e-1
+ pscbe2 = 1.317320208e-08 lpscbe2 = -6.243260025e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.715141667e-11 lalpha0 = 1.346934531e-15
+ alpha1 = -6.715141667e-11 lalpha1 = 1.346934531e-15
+ beta0 = 4.592926334e+01 lbeta0 = -3.195118720e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.877417733e-09 lagidl = -1.960004808e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -4.274405672e-01 legidl = 1.057949256e-05 pegidl = 2.131628207e-26
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.365567770e-01 lkt1 = -3.396295421e-8
+ kt2 = -6.270101271e-02 lkt2 = 8.334195126e-8
+ at = 1.186607907e+05 lat = -9.561888237e-1
+ ute = -4.988367220e-02 lute = -6.638517694e-7
+ ua1 = 2.269813722e-09 lua1 = -3.602722566e-15
+ ub1 = -1.573394235e-18 lub1 = 6.909923924e-24
+ uc1 = -4.390941745e-11 luc1 = 2.832297336e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.110 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 8.2e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.119308571e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.365284442e-9
+ k1 = 4.557431136e-01 lk1 = -6.628186177e-8
+ k2 = 1.736465621e-02 lk2 = 1.831987716e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.866729821e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.386030771e-8
+ nfactor = {1.917980732e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.308849687e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 9.209108364e-03 lu0 = 1.007203851e-9
+ ua = -7.714556020e-10 lua = 3.753057380e-16
+ ub = 1.139159733e-18 lub = -5.626103368e-25
+ uc = -7.082993503e-11 luc = -7.630877232e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.687361861e+05 lvsat = -8.737166397e-1
+ a0 = 1.298282802e+00 la0 = -9.606370240e-7
+ ags = 3.007947423e-01 lags = 1.018976364e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.275546728e-04 lketa = -8.401813297e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.415723457e-01 lpclm = -8.107596053e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -1.412456511e-03 lpdiblc2 = 1.395477241e-08 wpdiblc2 = -3.469446952e-24 ppdiblc2 = -1.387778781e-29
+ pdiblcb = -2.502133320e-01 lpdiblcb = 7.662820228e-7
+ drout = 0.56
+ pscbe1 = 1.230892076e+09 lpscbe1 = -3.472594437e+3
+ pscbe2 = -1.731012336e-08 lpscbe2 = 1.832072184e-13 ppscbe2 = 2.117582368e-34
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.405041024e+00 lbeta0 = 2.315554051e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.940678393e-10 lagidl = -2.006243465e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 1.682321702e+00 legidl = -6.421330460e-6
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.058118873e-01 lkt1 = -2.817105026e-7
+ kt2 = -4.835860979e-02 lkt2 = -3.223156969e-8
+ at = -9.199465573e+04 lat = 7.413085750e-1
+ ute = -1.650014701e-01 lute = 2.637870157e-7
+ ua1 = 5.595420866e-10 lua1 = 1.017893702e-14
+ ub1 = 8.371840607e-19 lub1 = -1.251492578e-23
+ uc1 = -1.167338578e-11 luc1 = 2.346631032e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.111 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 8.2e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.116324143e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.347660345e-8
+ k1 = 4.428654258e-01 lk1 = -1.402201541e-8
+ k2 = 2.164134381e-02 lk2 = 9.643518320e-10
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.673887289e-01 ldsub = -1.247435718e-06 wdsub = -3.552713679e-21
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.076298863e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.118637217e-8
+ nfactor = {8.205595117e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.144672185e-6
+ eta0 = 1.618122575e-01 leta0 = -3.320080490e-7
+ etab = -1.415226926e-01 letab = 2.902512456e-7
+ u0 = 8.961795572e-03 lu0 = 2.010841203e-9
+ ua = -8.686534836e-10 lua = 7.697512652e-16
+ ub = 1.145979433e-18 lub = -5.902858386e-25
+ uc = -7.565336861e-11 luc = 1.194343622e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 53438.0
+ a0 = 1.058775121e+00 la0 = 1.132585948e-8
+ ags = 1.699111794e-01 lags = 6.330453849e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.740613019e-03 lketa = -3.911472438e-08 pketa = 5.551115123e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.662082328e-01 lpclm = 2.467351305e-06 wpclm = -4.440892099e-22 ppclm = -6.217248938e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 3.668885335e-03 lpdiblc2 = -6.666176630e-9
+ pdiblcb = -9.883598245e-02 lpdiblcb = 1.519670040e-7
+ drout = 0.56
+ pscbe1 = -5.399535418e+07 lpscbe1 = 1.741697186e+3
+ pscbe2 = 4.685632485e-08 lpscbe2 = -7.719113680e-14 ppscbe2 = -4.235164736e-34
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.151404795e+01 lbeta0 = -9.752188105e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.711119258e-10 lagidl = -2.898164661e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.817235263e-01 lkt1 = 2.635183383e-8
+ kt2 = -6.035456581e-02 lkt2 = 1.645005918e-8
+ at = 1.024940121e+05 lat = -4.795950233e-2
+ ute = -1.332981033e-01 lute = 1.351293641e-7
+ ua1 = 3.328055596e-09 lua1 = -1.056161454e-15
+ ub1 = -2.852522340e-18 lub1 = 2.458530043e-24
+ uc1 = 1.859730957e-11 luc1 = -9.937731742e-17 puc1 = -1.033975766e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.112 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 8.2e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.127136425e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.776911808e-9
+ k1 = 3.512559901e-01 lk1 = 1.745257769e-7
+ k2 = 5.719390124e-02 lk2 = -7.220885529e-08 pk2 = 2.220446049e-28
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.841659314e-01 ldsub = 1.122659537e-06 pdsub = -1.776356839e-27
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.937752555e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.671186683e-9
+ nfactor = {2.152613232e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.969208211e-7
+ eta0 = -2.317683150e-01 leta0 = 4.780476779e-07 weta0 = 3.608224830e-22 peta0 = 7.042977312e-28
+ etab = 8.728991787e-01 letab = -1.797601417e-06 wetab = -7.702172233e-22 petab = -9.887923813e-28
+ u0 = 9.740710576e-03 lu0 = 4.077017098e-10
+ ua = -8.760198240e-11 lua = -8.377855030e-16
+ ub = 1.194459582e-19 lub = 1.522494564e-24
+ uc = -7.526918424e-11 luc = 1.115271947e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.984839386e+04 lvsat = -1.319368033e-2
+ a0 = 1.446042456e+00 la0 = -7.857361509e-7
+ ags = 1.631988120e-01 lags = 6.468605781e-7
+ a1 = 0.0
+ a2 = 5.883765817e-01 la2 = 4.355569708e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.074975873e-02 lketa = -3.116565955e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.490103892e-01 lpclm = 3.778587940e-7
+ pdiblc1 = 7.614176700e-01 lpdiblc1 = -7.644407059e-07 ppdiblc1 = 3.552713679e-27
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 9.440520000e-02 ldrout = 9.582732495e-7
+ pscbe1 = 7.985241057e+08 lpscbe1 = -1.293279044e+1
+ pscbe2 = 9.536577846e-09 lpscbe2 = -3.807531059e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.831389756e+00 lbeta0 = 1.943688500e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.694326460e-10 lagidl = 8.227161552e-16 pagidl = -1.654361225e-36
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.581851405e-01 lkt1 = -2.209416583e-8
+ kt2 = -5.638602898e-02 lkt2 = 8.282135728e-9
+ at = 9.763617505e+04 lat = -3.796124776e-2
+ ute = 9.699104623e-01 lute = -2.135461409e-06 wute = -4.440892099e-22 pute = -1.776356839e-27
+ ua1 = 6.248983323e-09 lua1 = -7.067927273e-15
+ ub1 = -4.359386902e-18 lub1 = 5.559913481e-24
+ uc1 = -1.319123403e-10 luc1 = 2.103971287e-16 puc1 = 4.135903063e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.113 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 8.2e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.154593399e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.783105829e-8
+ k1 = 5.233778534e-01 lk1 = -7.608415156e-9
+ k2 = -1.577976505e-02 lk2 = 5.009689160e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.287002896e+00 ldsub = -5.399041805e-07 wdsub = 7.105427358e-21
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.727187927e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.961013053e-8
+ nfactor = {1.040699630e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.796727960e-7
+ eta0 = -3.970646192e-02 leta0 = 2.748135868e-7
+ etab = -1.747121215e+00 letab = 9.748255624e-7
+ u0 = 1.432027652e-02 lu0 = -4.438257587e-9
+ ua = -5.206791442e-10 lua = -3.795162426e-16
+ ub = 1.917792099e-18 lub = -3.804613713e-25
+ uc = -1.021917457e-10 luc = 3.964136635e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -6.521687765e+04 lvsat = 1.191466380e-1
+ a0 = 6.545658119e-01 la0 = 5.178068979e-8
+ ags = 2.436803301e-01 lags = 5.616974501e-7
+ a1 = 0.0
+ a2 = 1.054141277e+00 la2 = -5.730125626e-8
+ b0 = -9.791128221e-17 lb0 = 1.036067815e-22
+ b1 = -4.070620229e-20 lb1 = 4.307408208e-26
+ keta = 1.362598715e-02 lketa = -2.891024897e-08 pketa = 5.551115123e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.639864835e+00 lpclm = -8.822676549e-07 wpclm = 7.105427358e-21
+ pdiblc1 = 6.516146082e-02 lpdiblc1 = -2.768327299e-8
+ pdiblc2 = 7.991361598e-04 lpdiblc2 = -3.906088102e-10 ppdiblc2 = -1.734723476e-30
+ pdiblcb = -1.332254979e-02 lpdiblcb = -1.235672748e-8
+ drout = 1.042241597e+00 ldrout = -4.469879061e-8
+ pscbe1 = 8.282864975e+08 lpscbe1 = -4.442646058e+1
+ pscbe2 = 3.048636988e-09 lpscbe2 = 6.484591271e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.485633595e+00 lbeta0 = 1.251387297e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.075221224e-09 lagidl = -6.001562308e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.178852899e-01 lkt1 = -6.473825875e-8
+ kt2 = -6.397594635e-02 lkt2 = 1.631355860e-8
+ at = 8.764820671e+04 lat = -2.739227930e-2
+ ute = -1.993146628e+00 lute = 9.999567120e-7
+ ua1 = -3.697989286e-09 lua1 = 3.457660733e-15 pua1 = 6.617444900e-36
+ ub1 = 4.480108576e-18 lub1 = -3.793775449e-24 wub1 = 6.162975822e-39
+ uc1 = 3.486000352e-10 luc1 = -2.980666517e-16 puc1 = -4.135903063e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.114 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 8.2e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.098276299e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.396542597e-9
+ k1 = 4.257803294e-01 lk1 = 4.686759479e-8
+ k2 = 3.182319986e-02 lk2 = -2.156085776e-08 pk2 = -2.775557562e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.533005469e-01 ldsub = 3.198469920e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.483210014e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.258875430e-8
+ nfactor = {2.949899408e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.859852442e-7
+ eta0 = 4.065893232e-01 leta0 = 2.570466844e-8
+ etab = -1.371832211e-03 letab = 4.006295315e-10
+ u0 = 7.628780961e-03 lu0 = -7.032655101e-10
+ ua = -1.951245750e-09 lua = 4.189831196e-16
+ ub = 2.631040349e-18 lub = -7.785751474e-25
+ uc = -6.837589508e-11 luc = 2.076637300e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.179337001e+05 lvsat = 1.691748002e-2
+ a0 = 9.109963816e-01 la0 = -9.135116129e-8
+ ags = 9.336688756e-01 lags = 1.765665437e-7
+ a1 = 0.0
+ a2 = 1.143114794e+00 la2 = -1.069636043e-7
+ b0 = -1.271017328e-15 lb0 = 7.583993833e-22 wb0 = -7.888609052e-37 pb0 = 1.183291358e-42
+ b1 = 3.942634583e-18 lb1 = -2.180307244e-24 wb1 = 3.081487911e-39 pb1 = 3.274080905e-45
+ keta = -4.608909199e-02 lketa = 4.420916754e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.532423753e-01 lpclm = 3.976759966e-07 wpclm = 4.440892099e-22 ppclm = -4.440892099e-28
+ pdiblc1 = -4.640274633e-01 lpdiblc1 = 2.676941088e-07 wpdiblc1 = -7.771561172e-22 ppdiblc1 = -1.110223025e-28
+ pdiblc2 = -1.035031450e-02 lpdiblc2 = 5.832680064e-09 wpdiblc2 = -5.204170428e-24 ppdiblc2 = -1.322726650e-29
+ pdiblcb = 2.758644106e-01 lpdiblcb = -1.737722132e-07 wpdiblcb = 4.440892099e-22 ppdiblcb = 4.440892099e-28
+ drout = 1.496502075e+00 ldrout = -2.982533618e-07 wdrout = -7.105427358e-21
+ pscbe1 = 6.854817729e+08 lpscbe1 = 3.528285254e+1
+ pscbe2 = 2.184228811e-08 lpscbe2 = -4.005460978e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.502780999e+00 lbeta0 = 1.254761302e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.261721264e-12 lagidl = -1.262424958e-18
+ bgidl = 7.033052157e+08 lbgidl = 1.656061277e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.00081386752815302
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207367379934e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.477070908e-01 lkt1 = 7.724375894e-9
+ kt2 = -1.248182315e-02 lkt2 = -1.242891616e-8
+ at = 2.437475586e+03 lat = 2.016979449e-2
+ ute = 5.785487810e-01 lute = -4.354865146e-07 pute = -4.440892099e-28
+ ua1 = 5.210530986e-09 lua1 = -1.514808027e-15
+ ub1 = -4.963733815e-18 lub1 = 1.477494058e-24
+ uc1 = -2.932921455e-10 luc1 = 6.021830677e-17 wuc1 = 1.654361225e-30
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.115 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 8.2e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.425443662e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.072197087e-07 wvth0 = 2.752475156e-07 pvth0 = -8.482302689e-14
+ k1 = -1.614380478e+00 lk1 = 6.755839509e-07 wk1 = 2.870674700e-07 pk1 = -8.846558223e-14
+ k2 = -1.527986494e-01 lk2 = 3.533405753e-08 wk2 = 5.808759670e-07 pk2 = -1.790085468e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 3.607758708e+00 ldsub = -8.700156386e-07 wdsub = -9.140307082e-07 pdsub = 2.816768434e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {7.017265876e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.701874112e-07 wvoff = -5.934496709e-07 pvoff = 1.828833851e-13
+ nfactor = {-9.133380099e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.237719001e-06 wnfactor = 6.717245552e-06 pnfactor = -2.070053562e-12
+ eta0 = 3.973435074e+00 leta0 = -1.073490187e-06 weta0 = -1.940001657e-06 peta0 = 5.978503106e-13
+ etab = 3.505557030e-01 letab = -1.080528790e-07 wetab = -1.950985312e-07 petab = 6.012351435e-14
+ u0 = -1.127474389e-01 lu0 = 3.639307418e-08 wu0 = 8.699762574e-08 pu0 = -2.681005833e-14
+ ua = -6.254698954e-09 lua = 1.745178294e-15 wua = 5.105689976e-15 pua = -1.573420480e-21
+ ub = 9.403636789e-19 lub = -2.575593179e-25 wub = -2.015635362e-24 pub = 6.211583495e-31
+ uc = -1.350796830e-10 luc = 4.132247933e-17 wuc = 9.872541811e-17 puc = -3.042421210e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.243370564e+07 lvsat = -9.941833959e+00 wvsat = -2.420002778e+01 pvsat = 7.457722562e-6
+ a0 = -3.577457238e+00 la0 = 1.291855591e-06 wa0 = 1.837098826e-06 pa0 = -5.661387451e-13
+ ags = 2.379754019e+00 lags = -2.690735150e-07 wags = -2.482957484e-14 pags = 7.651728140e-21
+ a1 = 0.0
+ a2 = 2.315094335e+00 la2 = -4.681325395e-07 wa2 = -7.614134227e-07 pa2 = 2.346447745e-13
+ b0 = -1.102019744e-05 lb0 = 3.396094245e-12 wb0 = 8.492210255e-12 pb0 = -2.617044434e-18
+ b1 = -6.322399300e-14 lb1 = 1.948277262e-20 wb1 = 3.520320204e-20 pb1 = -1.084857077e-26
+ keta = -2.686774101e-01 lketa = 7.301595873e-08 wketa = 9.559583797e-08 pketa = -2.945976939e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.759765930e-01 lpclm = -1.194941282e-08 wpclm = 9.600826471e-09 ppclm = -2.958686693e-15
+ pdiblc1 = 3.031697176e+00 lpdiblc1 = -8.095833533e-07 wpdiblc1 = -1.378380724e-06 ppdiblc1 = 4.247755877e-13
+ pdiblc2 = -8.587854913e-04 lpdiblc2 = 2.907675570e-09 wpdiblc2 = 1.929099685e-08 ppdiblc2 = -5.944906500e-15
+ pdiblcb = -7.357524250e+00 lpdiblcb = 2.178609170e-06 wpdiblcb = 5.587142090e-06 ppdiblcb = -1.721789578e-12
+ drout = -1.074949400e+00 ldrout = 4.941908394e-07 wdrout = 1.120598256e-12 pdrout = -3.453347688e-19
+ pscbe1 = 7.998824399e+08 lpscbe1 = 2.799899600e-02 wpscbe1 = -3.356353760e-06 ppscbe1 = 1.034328461e-12
+ pscbe2 = -7.780222608e-09 lpscbe2 = 5.123308152e-15 wpscbe2 = 1.636059394e-14 ppscbe2 = -5.041844234e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.083435857e+01 lbeta0 = -5.930461286e-07 wbeta0 = -1.831171567e-08 pbeta0 = 5.643121418e-15
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.973257276e-08 lagidl = 9.162121516e-15 wagidl = 2.190859892e-14 pagidl = -6.751572928e-21
+ bgidl = 2.059624098e+09 lbgidl = -2.523706621e+02 wbgidl = -1.245748901e-05 pbgidl = 3.839019775e-12
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.00081386752815302
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207367379934e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -9.539742204e-01 lkt1 = 1.329237172e-07 wkt1 = 3.615827610e-07 pkt1 = -1.114289594e-13
+ kt2 = 5.370217045e-01 lkt2 = -1.817694183e-07 wkt2 = -3.345698207e-07 pkt2 = 1.031043816e-13
+ at = -6.487415677e+04 lat = 4.091322023e-02 wat = 1.690691906e-01 pat = -5.210205247e-8
+ ute = -7.715440743e+00 lute = 2.120472237e-06 wute = 3.187660492e-06 pute = -9.823413338e-13
+ ua1 = -5.057032436e-09 lua1 = 1.649346992e-15 wua1 = 2.895931223e-15 pua1 = -8.924391249e-22
+ ub1 = 4.349547267e-18 lub1 = -1.392579773e-24 wub1 = -2.639375470e-24 pub1 = 8.133763386e-31
+ uc1 = -4.278515557e-10 luc1 = 1.016854802e-16 wuc1 = 5.416628198e-17 puc1 = -1.669242312e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.116 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 8.2e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -3.7585e-8
+ vth0 = {-9.877019919e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.174250880e-09 wvth0 = -7.148143777e-08 pvth0 = -2.402662870e-15
+ k1 = 1.222183289e+00 lk1 = -4.730905516e-13 wk1 = -8.437291471e-08 pk1 = 4.009047245e-19
+ k2 = -3.108482717e+00 lk2 = 7.920580207e-07 wk2 = 2.178792714e-06 pk2 = -5.995261612e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -4.516858891e-02 ldsub = 2.202478967e-12 wdsub = 2.686452677e-07 pdsub = -1.171902426e-18
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-4.327045731e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 6.249814888e-14 wvoff = 1.744195115e-07 pvoff = -1.938775185e-20
+ nfactor = {4.460766989e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.060078631e-12 wnfactor = -1.974247975e-06 pnfactor = -5.876839708e-19
+ eta0 = -5.338071192e-01 leta0 = -3.358259075e-13 weta0 = 5.701807245e-07 peta0 = 1.851715101e-19
+ etab = -1.031250668e-01 letab = 2.892096040e-13 wetab = 5.734155881e-08 petab = -1.520053525e-19
+ u0 = 2.053075635e-02 lu0 = 4.982126918e-09 wu0 = -1.079056785e-08 pu0 = -3.771082247e-15
+ ua = 1.074011371e-09 lua = -3.221038047e-19 wua = -1.501587012e-15 pua = 2.514312319e-25
+ ub = -1.410500722e-19 lub = 1.066259793e-30 wub = 5.924130195e-25 pub = -5.715911522e-37
+ uc = 3.842025846e-11 luc = -1.858469419e-24 wuc = -2.901616060e-17 puc = -3.175161975e-31
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.872837417e+06 lvsat = -3.618751337e+00 wvsat = -3.621886607e+00 pvsat = 2.739112522e-6
+ a0 = 1.846628526e+00 la0 = 1.161647546e-12 wa0 = -5.399341727e-07 pa0 = -8.526774025e-19
+ ags = 1.249999994e+00 lags = 1.290217710e-15 wags = 5.980808737e-14 pags = -1.339910227e-20
+ a1 = 0.0
+ a2 = 3.495549234e-01 la2 = -1.918162695e-14 wa2 = 2.237852231e-07 pa2 = 1.392614024e-20
+ b0 = -4.598634766e-06 lb0 = 1.999909112e-12 wb0 = 3.436492312e-12 pb0 = -1.513775205e-18
+ b1 = 1.857796618e-14 wb1 = -1.034649260e-20
+ keta = 3.789399842e-02 lketa = -1.645887490e-13 wketa = -2.809670840e-08 pketa = 9.040532479e-20
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.258043778e-01 lpclm = 1.110664201e-13 wpclm = -2.821502260e-09 ppclm = -6.498945737e-20
+ pdiblc1 = -3.674873658e-01 lpdiblc1 = 4.596202796e-13 wpdiblc1 = 4.051179988e-07 ppdiblc1 = -3.247182949e-19
+ pdiblc2 = 1.134957933e-02 lpdiblc2 = 9.984561733e-15 wpdiblc2 = -5.669756477e-09 ppdiblc2 = -4.156634426e-21
+ pdiblcb = 1.789758797e+00 lpdiblcb = 8.218082463e-13 wpdiblcb = -1.642102361e-06 ppdiblcb = -4.575190609e-19
+ drout = 1.000004908e+00 ldrout = -1.101582583e-12 wdrout = -2.711141263e-12 pdrout = 6.077610379e-19
+ pscbe1 = 7.999999842e+08 lpscbe1 = 3.725318909e-06 wpscbe1 = 1.236087036e-05 ppscbe1 = -2.902404785e-12
+ pscbe2 = 1.373091736e-08 lpscbe2 = -5.974726888e-23 wpscbe2 = -4.808507019e-15 ppscbe2 = 5.797315837e-28
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.344338710e+00 lbeta0 = 2.036374212e-12 wbeta0 = 5.385755724e-09 pbeta0 = -9.699650150e-19
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 8.736259242e-09 lagidl = -2.154858998e-22 wagidl = -6.439106825e-15 pagidl = 1.587963007e-28
+ bgidl = 1.000000406e+09 lbgidl = -9.371633911e-05 wbgidl = -2.645077515e-05 pbgidl = 7.683715820e-12
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -2.8385e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.958690043e-01 lkt1 = -2.165353550e-13 wkt1 = -1.062726209e-07 pkt1 = 1.680465687e-19
+ kt2 = -2.261694949e-01 lkt2 = -1.824726681e-13 wkt2 = 9.833209406e-08 pkt2 = 1.420688616e-19
+ at = 1.069072837e+05 lat = 3.702746658e-08 wat = -4.969062283e-02 pat = -2.968154708e-14
+ ute = 1.187746727e+00 lute = 8.293636933e-14 wute = -9.368779927e-07 pute = -3.112410329e-21
+ ua1 = 1.868043066e-09 lua1 = 1.885774775e-21 wua1 = -8.511316484e-16 pua1 = -1.243743032e-27
+ ub1 = -1.497452469e-18 lub1 = 1.652608869e-31 wub1 = 7.757326811e-25 pub1 = 3.239153164e-38
+ uc1 = -9.067130942e-13 luc1 = 2.898996504e-23 wuc1 = -1.591981252e-17 puc1 = -1.927415096e-29
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.117 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 7.9e-07 wmax = 8.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.143603+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43165561
+ k2 = 0.046387026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
+ voff = {-0.16725342+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.5720692+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.00827017
+ ua = -7.4124916e-10
+ ub = 6.3364395e-19
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = 5.7286e-9
+ b1 = 3.5674e-8
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.118 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 7.9e-07 wmax = 8.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.159803279e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.249479557e-7
+ k1 = 4.210039986e-01 lk1 = 2.136518329e-7
+ k2 = 6.434930204e-02 lk2 = -3.602903863e-7
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.172472591e-06 lcit = 1.303205335e-10 pcit = 1.355252716e-32
+ voff = {-1.497245500e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -3.515970554e-7
+ nfactor = {1.532188847e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.999269080e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 7.555725933e-03 lu0 = 1.433044056e-8
+ ua = -7.522405845e-10 lua = 2.204678604e-16
+ ub = 3.410671347e-19 lub = 5.868555500e-24
+ uc = -1.284179734e-10 luc = 4.564233263e-16 wuc = 4.135903063e-31
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.633145348e+04 lvsat = 1.079621904e+0
+ a0 = 1.655334532e+00 la0 = -3.837820560e-6
+ ags = -2.111356046e-02 lags = 2.695889464e-06 pags = -3.552713679e-27
+ a1 = 0.0
+ a2 = 1.084157408e+00 la2 = -2.289788703e-6
+ b0 = 9.575436055e-09 lb0 = -7.716049156e-14
+ b1 = 5.962959638e-08 lb1 = -4.805054247e-13
+ keta = 4.030454116e-02 lketa = -3.398512340e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.958323949e-02 lpclm = 1.696584997e-06 wpclm = 1.110223025e-22 ppclm = 8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 1.920375883e-03 lpdiblc2 = -1.290175761e-8
+ pdiblcb = -2.719257256e-01 lpdiblcb = 9.412441810e-7
+ drout = 0.56
+ pscbe1 = 8.000327363e+08 lpscbe1 = -6.566305840e-1
+ pscbe2 = 1.317320208e-08 lpscbe2 = -6.243260025e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.715141667e-11 lalpha0 = 1.346934531e-15
+ alpha1 = -6.715141667e-11 lalpha1 = 1.346934531e-15
+ beta0 = 4.592926334e+01 lbeta0 = -3.195118720e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.877417733e-09 lagidl = -1.960004808e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -4.274405672e-01 legidl = 1.057949256e-05 pegidl = 3.552713679e-27
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.365567770e-01 lkt1 = -3.396295421e-8
+ kt2 = -6.270101271e-02 lkt2 = 8.334195126e-8
+ at = 1.186607907e+05 lat = -9.561888237e-1
+ ute = -4.988367220e-02 lute = -6.638517694e-7
+ ua1 = 2.269813722e-09 lua1 = -3.602722566e-15
+ ub1 = -1.573394235e-18 lub1 = 6.909923924e-24
+ uc1 = -4.390941745e-11 luc1 = 2.832297336e-16 puc1 = -8.271806126e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.119 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 7.9e-07 wmax = 8.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.119308571e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.365284442e-9
+ k1 = 4.557431136e-01 lk1 = -6.628186177e-8
+ k2 = 1.736465621e-02 lk2 = 1.831987716e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.866729821e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.386030771e-8
+ nfactor = {1.917980732e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.308849687e-06 wnfactor = -7.105427358e-21
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 9.209108364e-03 lu0 = 1.007203851e-9
+ ua = -7.714556020e-10 lua = 3.753057380e-16
+ ub = 1.139159733e-18 lub = -5.626103368e-25
+ uc = -7.082993503e-11 luc = -7.630877232e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.687361861e+05 lvsat = -8.737166397e-1
+ a0 = 1.298282802e+00 la0 = -9.606370240e-7
+ ags = 3.007947423e-01 lags = 1.018976364e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.275546727e-04 lketa = -8.401813297e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.415723457e-01 lpclm = -8.107596053e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -1.412456511e-03 lpdiblc2 = 1.395477241e-08 ppdiblc2 = 1.387778781e-29
+ pdiblcb = -2.502133320e-01 lpdiblcb = 7.662820228e-7
+ drout = 0.56
+ pscbe1 = 1.230892076e+09 lpscbe1 = -3.472594437e+3
+ pscbe2 = -1.731012336e-08 lpscbe2 = 1.832072184e-13 wpscbe2 = 2.646977960e-29
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.405041024e+00 lbeta0 = 2.315554051e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.940678393e-10 lagidl = -2.006243465e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 1.682321702e+00 legidl = -6.421330460e-6
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.058118873e-01 lkt1 = -2.817105026e-7
+ kt2 = -4.835860979e-02 lkt2 = -3.223156969e-8
+ at = -9.199465573e+04 lat = 7.413085750e-1
+ ute = -1.650014701e-01 lute = 2.637870157e-7
+ ua1 = 5.595420866e-10 lua1 = 1.017893702e-14
+ ub1 = 8.371840607e-19 lub1 = -1.251492578e-23 pub1 = 1.232595164e-44
+ uc1 = -1.167338578e-11 luc1 = 2.346631032e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.120 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 7.9e-07 wmax = 8.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.116324143e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.347660345e-8
+ k1 = 4.428654258e-01 lk1 = -1.402201541e-8
+ k2 = 2.164134381e-02 lk2 = 9.643518320e-10
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.673887289e-01 ldsub = -1.247435718e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.076298863e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.118637217e-8
+ nfactor = {8.205595117e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.144672185e-6
+ eta0 = 1.618122575e-01 leta0 = -3.320080490e-7
+ etab = -1.415226926e-01 letab = 2.902512456e-7
+ u0 = 8.961795573e-03 lu0 = 2.010841203e-9
+ ua = -8.686534836e-10 lua = 7.697512652e-16
+ ub = 1.145979433e-18 lub = -5.902858386e-25
+ uc = -7.565336861e-11 luc = 1.194343622e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 53438.0
+ a0 = 1.058775121e+00 la0 = 1.132585948e-8
+ ags = 1.699111794e-01 lags = 6.330453849e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.740613018e-03 lketa = -3.911472438e-08 pketa = -2.775557562e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.662082328e-01 lpclm = 2.467351305e-06 wpclm = -6.661338148e-22 ppclm = -1.776356839e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 3.668885335e-03 lpdiblc2 = -6.666176630e-9
+ pdiblcb = -9.883598245e-02 lpdiblcb = 1.519670040e-7
+ drout = 0.56
+ pscbe1 = -5.399535418e+07 lpscbe1 = 1.741697186e+3
+ pscbe2 = 4.685632485e-08 lpscbe2 = -7.719113680e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.151404795e+01 lbeta0 = -9.752188105e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.711119258e-10 lagidl = -2.898164661e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.817235264e-01 lkt1 = 2.635183383e-8
+ kt2 = -6.035456581e-02 lkt2 = 1.645005918e-8
+ at = 1.024940121e+05 lat = -4.795950233e-2
+ ute = -1.332981033e-01 lute = 1.351293641e-7
+ ua1 = 3.328055597e-09 lua1 = -1.056161454e-15
+ ub1 = -2.852522340e-18 lub1 = 2.458530043e-24
+ uc1 = 1.859730957e-11 luc1 = -9.937731742e-17 wuc1 = 2.584939414e-32 puc1 = -5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.121 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 7.9e-07 wmax = 8.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.127136425e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.776911808e-9
+ k1 = 3.512559901e-01 lk1 = 1.745257769e-7
+ k2 = 5.719390124e-02 lk2 = -7.220885529e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.841659314e-01 ldsub = 1.122659537e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.937752555e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.671186683e-9
+ nfactor = {2.152613232e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.969208211e-7
+ eta0 = -2.317683150e-01 leta0 = 4.780476779e-07 weta0 = 4.232725281e-22 peta0 = -3.295974604e-28
+ etab = 8.728991787e-01 letab = -1.797601417e-06 wetab = -5.898059818e-22 petab = 1.144917494e-28
+ u0 = 9.740710576e-03 lu0 = 4.077017098e-10
+ ua = -8.760198240e-11 lua = -8.377855030e-16
+ ub = 1.194459582e-19 lub = 1.522494564e-24
+ uc = -7.526918424e-11 luc = 1.115271947e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.984839386e+04 lvsat = -1.319368033e-2
+ a0 = 1.446042456e+00 la0 = -7.857361509e-7
+ ags = 1.631988120e-01 lags = 6.468605781e-7
+ a1 = 0.0
+ a2 = 5.883765817e-01 la2 = 4.355569708e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.074975873e-02 lketa = -3.116565955e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.490103892e-01 lpclm = 3.778587940e-7
+ pdiblc1 = 7.614176700e-01 lpdiblc1 = -7.644407059e-07 ppdiblc1 = -1.776356839e-27
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 9.440520000e-02 ldrout = 9.582732495e-7
+ pscbe1 = 7.985241057e+08 lpscbe1 = -1.293279044e+1
+ pscbe2 = 9.536577846e-09 lpscbe2 = -3.807531059e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.831389756e+00 lbeta0 = 1.943688500e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.694326460e-10 lagidl = 8.227161552e-16 pagidl = 8.271806126e-37
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.581851405e-01 lkt1 = -2.209416583e-8
+ kt2 = -5.638602898e-02 lkt2 = 8.282135728e-9
+ at = 9.763617505e+04 lat = -3.796124776e-2
+ ute = 9.699104623e-01 lute = -2.135461409e-06 wute = 8.881784197e-22 pute = 8.881784197e-28
+ ua1 = 6.248983323e-09 lua1 = -7.067927273e-15
+ ub1 = -4.359386902e-18 lub1 = 5.559913481e-24
+ uc1 = -1.319123403e-10 luc1 = 2.103971287e-16 wuc1 = -2.067951531e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.122 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 7.9e-07 wmax = 8.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.154593399e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.783105829e-8
+ k1 = 5.233778534e-01 lk1 = -7.608415156e-9
+ k2 = -1.577976505e-02 lk2 = 5.009689160e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.287002896e+00 ldsub = -5.399041805e-07 wdsub = 3.552713679e-21
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.727187927e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.961013053e-8
+ nfactor = {1.040699630e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.796727960e-7
+ eta0 = -3.970646192e-02 leta0 = 2.748135868e-7
+ etab = -1.747121215e+00 letab = 9.748255624e-7
+ u0 = 1.432027652e-02 lu0 = -4.438257587e-9
+ ua = -5.206791442e-10 lua = -3.795162426e-16
+ ub = 1.917792099e-18 lub = -3.804613713e-25
+ uc = -1.021917457e-10 luc = 3.964136635e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -6.521687765e+04 lvsat = 1.191466380e-01 pvsat = -1.164153218e-22
+ a0 = 6.545658119e-01 la0 = 5.178068979e-8
+ ags = 2.436803301e-01 lags = 5.616974501e-7
+ a1 = 0.0
+ a2 = 1.054141277e+00 la2 = -5.730125626e-8
+ b0 = -9.791128221e-17 lb0 = 1.036067815e-22
+ b1 = -4.070620229e-20 lb1 = 4.307408208e-26
+ keta = 1.362598715e-02 lketa = -2.891024897e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.639864835e+00 lpclm = -8.822676549e-7
+ pdiblc1 = 6.516146082e-02 lpdiblc1 = -2.768327299e-08 wpdiblc1 = -2.220446049e-22
+ pdiblc2 = 7.991361598e-04 lpdiblc2 = -3.906088102e-10
+ pdiblcb = -1.332254979e-02 lpdiblcb = -1.235672748e-8
+ drout = 1.042241597e+00 ldrout = -4.469879061e-8
+ pscbe1 = 8.282864975e+08 lpscbe1 = -4.442646058e+1
+ pscbe2 = 3.048636988e-09 lpscbe2 = 6.484591271e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.485633595e+00 lbeta0 = 1.251387297e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.075221224e-09 lagidl = -6.001562308e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.178852899e-01 lkt1 = -6.473825875e-8
+ kt2 = -6.397594635e-02 lkt2 = 1.631355860e-08 wkt2 = 2.220446049e-22
+ at = 8.764820671e+04 lat = -2.739227930e-2
+ ute = -1.993146628e+00 lute = 9.999567120e-07 pute = -3.552713679e-27
+ ua1 = -3.697989286e-09 lua1 = 3.457660733e-15 pua1 = -1.654361225e-36
+ ub1 = 4.480108576e-18 lub1 = -3.793775449e-24 wub1 = -6.162975822e-39 pub1 = 3.081487911e-45
+ uc1 = 3.486000352e-10 luc1 = -2.980666517e-16 puc1 = -4.135903063e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.123 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 7.9e-07 wmax = 8.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.098276299e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.396542597e-9
+ k1 = 4.257803294e-01 lk1 = 4.686759479e-8
+ k2 = 3.182319986e-02 lk2 = -2.156085776e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.533005469e-01 ldsub = 3.198469920e-07 pdsub = 4.440892099e-28
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.483210014e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.258875430e-8
+ nfactor = {2.949899408e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.859852442e-7
+ eta0 = 4.065893232e-01 leta0 = 2.570466844e-8
+ etab = -1.371832211e-03 letab = 4.006295315e-10
+ u0 = 7.628780961e-03 lu0 = -7.032655101e-10 wu0 = -2.775557562e-23
+ ua = -1.951245750e-09 lua = 4.189831196e-16
+ ub = 2.631040349e-18 lub = -7.785751474e-25
+ uc = -6.837589508e-11 luc = 2.076637300e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.179337001e+05 lvsat = 1.691748002e-2
+ a0 = 9.109963816e-01 la0 = -9.135116129e-8
+ ags = 9.336688756e-01 lags = 1.765665437e-7
+ a1 = 0.0
+ a2 = 1.143114794e+00 la2 = -1.069636043e-7
+ b0 = -1.271017328e-15 lb0 = 7.583993833e-22 wb0 = 1.183291358e-36 pb0 = -5.916456789e-43
+ b1 = 3.942634583e-18 lb1 = -2.180307244e-24 wb1 = -2.118522939e-39 pb1 = 1.444447458e-45
+ keta = -4.608909199e-02 lketa = 4.420916754e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.532423753e-01 lpclm = 3.976759966e-07 ppclm = 3.330669074e-28
+ pdiblc1 = -4.640274633e-01 lpdiblc1 = 2.676941088e-07 wpdiblc1 = -3.330669074e-22 ppdiblc1 = -3.608224830e-28
+ pdiblc2 = -1.035031450e-02 lpdiblc2 = 5.832680064e-09 wpdiblc2 = 4.336808690e-24 ppdiblc2 = -2.385244779e-30
+ pdiblcb = 2.758644106e-01 lpdiblcb = -1.737722132e-07 wpdiblcb = -2.220446049e-22
+ drout = 1.496502075e+00 ldrout = -2.982533618e-7
+ pscbe1 = 6.854817729e+08 lpscbe1 = 3.528285254e+1
+ pscbe2 = 2.184228811e-08 lpscbe2 = -4.005460978e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.502780999e+00 lbeta0 = 1.254761302e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.261721264e-12 lagidl = -1.262424958e-18
+ bgidl = 7.033052157e+08 lbgidl = 1.656061277e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.00081386752815302
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207367379934e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.477070908e-01 lkt1 = 7.724375894e-9
+ kt2 = -1.248182315e-02 lkt2 = -1.242891616e-8
+ at = 2.437475586e+03 lat = 2.016979449e-2
+ ute = 5.785487810e-01 lute = -4.354865146e-07 wute = 8.881784197e-22
+ ua1 = 5.210530986e-09 lua1 = -1.514808027e-15
+ ub1 = -4.963733815e-18 lub1 = 1.477494058e-24
+ uc1 = -2.932921455e-10 luc1 = 6.021830677e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.124 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7.9e-07 wmax = 8.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.051933961e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.884775766e-9
+ k1 = -1.224831150e+00 lk1 = 5.555365344e-7
+ k2 = 6.354475517e-01 lk2 = -2.075797743e-07 wk2 = 4.440892099e-22
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.367422949e+00 ldsub = -4.877813677e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.035820758e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.201544042e-8
+ nfactor = {-1.810663453e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.286651779e-7
+ eta0 = 1.340861129e+00 leta0 = -2.622098740e-7
+ etab = 8.580783120e-02 letab = -2.646552734e-08 wetab = 2.081668171e-23 petab = -1.778091563e-29
+ u0 = 5.307966851e-03 lu0 = 1.193977425e-11
+ ua = 6.737004918e-10 lua = -3.899465637e-16
+ ub = -1.794844881e-18 lub = 5.853499039e-25 wub = -1.540743956e-39 pub = -3.851859889e-46
+ uc = -1.109713200e-12 luc = 3.695372767e-20
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -4.056284828e+05 lvsat = 1.782636380e-1
+ a0 = -1.084521995e+00 la0 = 5.236077367e-7
+ ags = 2.379753985e+00 lags = -2.690735046e-7
+ a1 = 0.0
+ a2 = 1.281859579e+00 la2 = -1.497205848e-7
+ b0 = 5.036955310e-07 lb0 = -1.552238514e-13 wb0 = 5.529275022e-28 pb0 = 1.240793165e-34
+ b1 = -1.545339850e-14 lb1 = 4.761308510e-21 wb1 = -8.036520472e-36 pb1 = 5.706915611e-42
+ keta = -1.389542671e-01 lketa = 3.303917776e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.890048734e-01 lpclm = -1.596433800e-8
+ pdiblc1 = 1.161240433e+00 lpdiblc1 = -2.331646988e-07 ppdiblc1 = 8.881784197e-28
+ pdiblc2 = 2.531901467e-02 lpdiblc2 = -5.159537107e-9
+ pdiblcb = 2.242036531e-01 lpdiblcb = -1.578519175e-7
+ drout = -1.074947880e+00 ldrout = 4.941903708e-7
+ pscbe1 = 7.998824353e+08 lpscbe1 = 2.800039958e-2
+ pscbe2 = 1.442103334e-08 lpscbe2 = -1.718452894e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.080950965e+01 lbeta0 = -5.853884369e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.697791983e-12 lagidl = 2.659482394e-19
+ bgidl = 2.059624081e+09 lbgidl = -2.523706569e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.00081386752815302
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207367379934e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.633079613e-01 lkt1 = -1.828490384e-8
+ kt2 = 8.301188984e-02 lkt2 = -4.185721369e-8
+ at = 1.645520113e+05 lat = -2.978904198e-2
+ ute = -3.389799098e+00 lute = 7.874392514e-7
+ ua1 = -1.127266161e-09 lua1 = 4.383109196e-16
+ ub1 = 7.679260506e-19 lub1 = -2.888315626e-25
+ uc1 = -3.543481429e-10 luc1 = 7.903393350e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.125 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7.9e-07 wmax = 8.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -3.7585e-8
+ vth0 = {-1.803182576e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.832485370e-07 wvth0 = 5.294641452e-07 pvth0 = -1.351033659e-13
+ k1 = 2.530924127e-01 lk1 = 2.180676365e-07 wk1 = 6.297714720e-07 pk1 = -1.606987865e-13
+ k2 = -6.736204000e-02 lk2 = -4.306039424e-08 wk2 = -6.227601752e-08 pk2 = 1.589097139e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 3.040443347e+00 ldsub = -6.943326399e-07 wdsub = -2.005210051e-06 pdsub = 5.116694488e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {1.580472589e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.533070783e-07 wvoff = -1.309135029e-06 pvoff = 3.340519854e-13
+ nfactor = {-1.832633365e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.130972551e-06 wnfactor = 1.481806780e-05 pnfactor = -3.781126361e-12
+ eta0 = 6.047313612e+00 leta0 = -1.481871262e-06 weta0 = -4.279591927e-06 peta0 = 1.092023472e-12
+ etab = 5.554943358e-01 letab = -1.482044782e-07 wetab = -4.280095686e-07 petab = 1.092152016e-13
+ u0 = -5.112236642e-02 lu0 = 1.441212015e-08 wu0 = 4.201219468e-08 pu0 = -1.072025172e-14
+ ua = -1.624581782e-08 lua = 3.899573479e-15 wua = 1.126177616e-14 pua = -2.873667422e-21
+ ub = 6.695056422e-18 lub = -1.539237348e-24 wub = -4.445264251e-24 pub = 1.134298079e-30
+ uc = -2.948599301e-10 luc = 7.499583424e-17 wuc = 2.165853425e-16 puc = -5.526608185e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -5.043338314e+05 lvsat = 2.161743101e-01 wvsat = 3.406691839e-01 pvsat = -8.692855566e-8
+ a0 = -4.385411395e+00 la0 = 1.403269542e-06 wa0 = 4.052593150e-06 pa0 = -1.034100194e-12
+ ags = 1.250000075e+00 lags = -1.689230800e-14
+ a1 = 0.0
+ a2 = 2.919956882e+00 la2 = -5.784005676e-07 wa2 = -1.670400529e-06 pa2 = 4.262361029e-13
+ b0 = 1.649372300e-06 lb0 = -4.586456965e-13 wb0 = -1.167801551e-12 pb0 = 2.979879217e-19
+ b1 = -1.008413062e-13 lb1 = 2.688959163e-20 wb1 = 7.765619642e-20 pb1 = -1.981553164e-26
+ keta = -2.863984327e-01 lketa = 7.302076231e-08 wketa = 2.108815185e-07 pketa = -5.381063709e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.933936123e-01 lpclm = 7.293291559e-09 wpclm = 2.106270386e-08 ppclm = -5.374570145e-15
+ pdiblc1 = 4.285691073e+00 lpdiblc1 = -1.047073502e-06 wpdiblc1 = -3.023911563e-06 ppdiblc1 = 7.716115134e-13
+ pdiblc2 = -5.377353945e-02 lpdiblc2 = 1.465423462e-08 wpdiblc2 = 4.232090247e-08 ppdiblc2 = -1.079902468e-14
+ pdiblcb = -1.707148083e+01 lpdiblcb = 4.244220802e-06 wpdiblcb = 1.225716007e-05 ppdiblcb = -3.127659534e-12
+ drout = 1.000001229e+00 ldrout = -2.768534628e-13
+ pscbe1 = 8.000000009e+08 lpscbe1 = -2.132339478e-7
+ pscbe2 = -4.149965967e-08 lpscbe2 = 1.242817132e-14 wpscbe2 = 3.589212027e-14 ppscbe2 = -9.158592330e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.406156022e+00 lbeta0 = -1.390830688e-08 wbeta0 = -4.016878163e-08 pbeta0 = 1.024986801e-14
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -3.528826449e-10 lagidl = 8.964159991e-17 wagidl = 2.588817929e-16 pagidl = -6.605886709e-23
+ bgidl = 1.000000370e+09 lbgidl = -8.328957367e-5
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -2.8385e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.622476916e+00 lkt1 = 2.761951060e-07 wkt1 = 7.976417347e-07 pkt1 = -2.035342415e-13
+ kt2 = 9.032812045e-01 lkt2 = -2.541530016e-07 wkt2 = -7.339849742e-07 pkt2 = 1.872909459e-13
+ at = -4.638414938e+05 lat = 1.284318588e-01 wat = 3.709067078e-01 pat = -9.464426463e-8
+ ute = -9.573251807e+00 lute = 2.421476393e-06 wute = 6.993138569e-06 pute = -1.784439169e-12
+ ua1 = -7.908127221e-09 lua1 = 2.199868812e-15 wua1 = 6.353143312e-15 pua1 = -1.621131579e-21
+ ub1 = 7.412629296e-18 lub1 = -2.004976590e-24 wub1 = -5.790302593e-24 pub1 = 1.477511513e-30
+ uc1 = -1.837628492e-10 luc1 = 4.114693562e-17 wuc1 = 1.188308970e-16 puc1 = -3.032208000e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.126 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 7.5e-07 wmax = 7.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.143603+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43165561
+ k2 = 0.046387026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
+ voff = {-0.16725342+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.5720692+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.00827017
+ ua = -7.4124916e-10
+ ub = 6.3364395e-19
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = 5.7286e-9
+ b1 = 3.5674e-8
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.127 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 7.5e-07 wmax = 7.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.159803279e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.249479557e-7
+ k1 = 4.210039986e-01 lk1 = 2.136518329e-7
+ k2 = 6.434930204e-02 lk2 = -3.602903863e-7
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.172472591e-06 lcit = 1.303205335e-10 wcit = -2.541098842e-27 pcit = 1.355252716e-32
+ voff = {-1.497245500e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -3.515970554e-7
+ nfactor = {1.532188847e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 7.999269080e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 7.555725933e-03 lu0 = 1.433044056e-8
+ ua = -7.522405845e-10 lua = 2.204678604e-16
+ ub = 3.410671347e-19 lub = 5.868555500e-24
+ uc = -1.284179734e-10 luc = 4.564233263e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.633145348e+04 lvsat = 1.079621904e+0
+ a0 = 1.655334532e+00 la0 = -3.837820560e-06 wa0 = 3.552713679e-21
+ ags = -2.111356046e-02 lags = 2.695889464e-6
+ a1 = 0.0
+ a2 = 1.084157408e+00 la2 = -2.289788703e-6
+ b0 = 9.575436055e-09 lb0 = -7.716049156e-14
+ b1 = 5.962959638e-08 lb1 = -4.805054247e-13
+ keta = 4.030454116e-02 lketa = -3.398512340e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.958323949e-02 lpclm = 1.696584997e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 1.920375883e-03 lpdiblc2 = -1.290175761e-8
+ pdiblcb = -2.719257256e-01 lpdiblcb = 9.412441810e-7
+ drout = 0.56
+ pscbe1 = 8.000327363e+08 lpscbe1 = -6.566305840e-1
+ pscbe2 = 1.317320208e-08 lpscbe2 = -6.243260025e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.715141667e-11 lalpha0 = 1.346934531e-15
+ alpha1 = -6.715141667e-11 lalpha1 = 1.346934531e-15
+ beta0 = 4.592926334e+01 lbeta0 = -3.195118720e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.877417733e-09 lagidl = -1.960004808e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -4.274405672e-01 legidl = 1.057949256e-05 wegidl = -2.220446049e-22 pegidl = -1.776356839e-27
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.365567770e-01 lkt1 = -3.396295421e-8
+ kt2 = -6.270101271e-02 lkt2 = 8.334195126e-8
+ at = 1.186607907e+05 lat = -9.561888237e-1
+ ute = -4.988367220e-02 lute = -6.638517694e-7
+ ua1 = 2.269813722e-09 lua1 = -3.602722566e-15
+ ub1 = -1.573394235e-18 lub1 = 6.909923924e-24
+ uc1 = -4.390941745e-11 luc1 = 2.832297336e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.128 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 7.5e-07 wmax = 7.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.119308571e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.365284442e-9
+ k1 = 4.557431136e-01 lk1 = -6.628186177e-8
+ k2 = 1.736465621e-02 lk2 = 1.831987716e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.866729821e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.386030771e-8
+ nfactor = {1.917980732e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.308849687e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 9.209108364e-03 lu0 = 1.007203851e-9
+ ua = -7.714556020e-10 lua = 3.753057380e-16
+ ub = 1.139159733e-18 lub = -5.626103368e-25
+ uc = -7.082993503e-11 luc = -7.630877232e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.687361861e+05 lvsat = -8.737166397e-1
+ a0 = 1.298282802e+00 la0 = -9.606370240e-7
+ ags = 3.007947423e-01 lags = 1.018976364e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.275546727e-04 lketa = -8.401813297e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.415723457e-01 lpclm = -8.107596053e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -1.412456511e-03 lpdiblc2 = 1.395477241e-08 ppdiblc2 = 6.938893904e-30
+ pdiblcb = -2.502133320e-01 lpdiblcb = 7.662820228e-07 wpdiblcb = -4.440892099e-22
+ drout = 0.56
+ pscbe1 = 1.230892076e+09 lpscbe1 = -3.472594437e+3
+ pscbe2 = -1.731012336e-08 lpscbe2 = 1.832072184e-13
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.405041024e+00 lbeta0 = 2.315554051e-5
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.940678393e-10 lagidl = -2.006243465e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 1.682321702e+00 legidl = -6.421330460e-6
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.058118873e-01 lkt1 = -2.817105026e-7
+ kt2 = -4.835860979e-02 lkt2 = -3.223156969e-8
+ at = -9.199465573e+04 lat = 7.413085750e-1
+ ute = -1.650014701e-01 lute = 2.637870157e-7
+ ua1 = 5.595420866e-10 lua1 = 1.017893702e-14
+ ub1 = 8.371840607e-19 lub1 = -1.251492578e-23
+ uc1 = -1.167338578e-11 luc1 = 2.346631032e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.129 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 7.5e-07 wmax = 7.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.116324143e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.347660345e-8
+ k1 = 4.428654258e-01 lk1 = -1.402201541e-8
+ k2 = 2.164134381e-02 lk2 = 9.643518320e-10
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.673887289e-01 ldsub = -1.247435718e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.076298863e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.118637217e-8
+ nfactor = {8.205595117e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.144672185e-6
+ eta0 = 1.618122575e-01 leta0 = -3.320080490e-7
+ etab = -1.415226926e-01 letab = 2.902512456e-7
+ u0 = 8.961795572e-03 lu0 = 2.010841203e-9
+ ua = -8.686534836e-10 lua = 7.697512652e-16
+ ub = 1.145979433e-18 lub = -5.902858386e-25
+ uc = -7.565336861e-11 luc = 1.194343622e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 53438.0
+ a0 = 1.058775121e+00 la0 = 1.132585948e-8
+ ags = 1.699111794e-01 lags = 6.330453849e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.740613018e-03 lketa = -3.911472438e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.662082328e-01 lpclm = 2.467351305e-06 wpclm = 1.110223025e-22 ppclm = -1.332267630e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 3.668885335e-03 lpdiblc2 = -6.666176630e-9
+ pdiblcb = -9.883598245e-02 lpdiblcb = 1.519670040e-7
+ drout = 0.56
+ pscbe1 = -5.399535418e+07 lpscbe1 = 1.741697186e+3
+ pscbe2 = 4.685632485e-08 lpscbe2 = -7.719113680e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.151404795e+01 lbeta0 = -9.752188105e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.711119258e-10 lagidl = -2.898164661e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.817235263e-01 lkt1 = 2.635183383e-8
+ kt2 = -6.035456582e-02 lkt2 = 1.645005918e-8
+ at = 1.024940121e+05 lat = -4.795950233e-2
+ ute = -1.332981033e-01 lute = 1.351293641e-7
+ ua1 = 3.328055597e-09 lua1 = -1.056161454e-15
+ ub1 = -2.852522340e-18 lub1 = 2.458530043e-24
+ uc1 = 1.859730957e-11 luc1 = -9.937731742e-17 puc1 = 5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.130 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 7.5e-07 wmax = 7.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.127136425e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.776911808e-9
+ k1 = 3.512559901e-01 lk1 = 1.745257769e-7
+ k2 = 5.719390124e-02 lk2 = -7.220885529e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.841659314e-01 ldsub = 1.122659537e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.937752555e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.671186683e-9
+ nfactor = {2.152613232e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.969208211e-7
+ eta0 = -2.317683150e-01 leta0 = 4.780476779e-07 weta0 = -1.058181320e-22 peta0 = -3.920475056e-28
+ etab = 8.728991787e-01 letab = -1.797601417e-06 wetab = 8.847089727e-22 petab = 1.335737077e-28
+ u0 = 9.740710576e-03 lu0 = 4.077017098e-10
+ ua = -8.760198240e-11 lua = -8.377855030e-16
+ ub = 1.194459582e-19 lub = 1.522494564e-24
+ uc = -7.526918424e-11 luc = 1.115271947e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.984839386e+04 lvsat = -1.319368033e-2
+ a0 = 1.446042456e+00 la0 = -7.857361509e-7
+ ags = 1.631988120e-01 lags = 6.468605781e-7
+ a1 = 0.0
+ a2 = 5.883765817e-01 la2 = 4.355569708e-7
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.074975873e-02 lketa = -3.116565955e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.490103892e-01 lpclm = 3.778587940e-7
+ pdiblc1 = 7.614176700e-01 lpdiblc1 = -7.644407059e-7
+ pdiblc2 = 0.00043
+ pdiblcb = -0.025
+ drout = 9.440520000e-02 ldrout = 9.582732495e-7
+ pscbe1 = 7.985241057e+08 lpscbe1 = -1.293279044e+1
+ pscbe2 = 9.536577846e-09 lpscbe2 = -3.807531059e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 5.831389756e+00 lbeta0 = 1.943688500e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.694326460e-10 lagidl = 8.227161552e-16 pagidl = 4.135903063e-37
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.581851405e-01 lkt1 = -2.209416583e-8
+ kt2 = -5.638602898e-02 lkt2 = 8.282135728e-9
+ at = 9.763617505e+04 lat = -3.796124776e-2
+ ute = 9.699104623e-01 lute = -2.135461409e-06 wute = 4.440892099e-22 pute = -2.220446049e-28
+ ua1 = 6.248983323e-09 lua1 = -7.067927273e-15 pua1 = 1.323488980e-35
+ ub1 = -4.359386902e-18 lub1 = 5.559913481e-24 pub1 = 6.162975822e-45
+ uc1 = -1.319123403e-10 luc1 = 2.103971287e-16 puc1 = 2.067951531e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.131 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 7.5e-07 wmax = 7.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.154593399e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.783105829e-8
+ k1 = 5.233778534e-01 lk1 = -7.608415156e-9
+ k2 = -1.577976505e-02 lk2 = 5.009689160e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.287002896e+00 ldsub = -5.399041805e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.727187927e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.961013053e-8
+ nfactor = {1.040699630e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.796727960e-7
+ eta0 = -3.970646192e-02 leta0 = 2.748135868e-7
+ etab = -1.747121215e+00 letab = 9.748255624e-7
+ u0 = 1.432027652e-02 lu0 = -4.438257587e-9
+ ua = -5.206791442e-10 lua = -3.795162426e-16
+ ub = 1.917792099e-18 lub = -3.804613713e-25
+ uc = -1.021917457e-10 luc = 3.964136635e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -6.521687765e+04 lvsat = 1.191466380e-01 pvsat = 1.164153218e-22
+ a0 = 6.545658119e-01 la0 = 5.178068979e-8
+ ags = 2.436803301e-01 lags = 5.616974501e-7
+ a1 = 0.0
+ a2 = 1.054141277e+00 la2 = -5.730125626e-8
+ b0 = -9.791128221e-17 lb0 = 1.036067815e-22
+ b1 = -4.070620229e-20 lb1 = 4.307408208e-26
+ keta = 1.362598715e-02 lketa = -2.891024897e-08 pketa = -2.775557562e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.639864835e+00 lpclm = -8.822676549e-7
+ pdiblc1 = 6.516146082e-02 lpdiblc1 = -2.768327299e-8
+ pdiblc2 = 7.991361598e-04 lpdiblc2 = -3.906088102e-10
+ pdiblcb = -1.332254979e-02 lpdiblcb = -1.235672748e-8
+ drout = 1.042241597e+00 ldrout = -4.469879061e-8
+ pscbe1 = 8.282864975e+08 lpscbe1 = -4.442646058e+1
+ pscbe2 = 3.048636988e-09 lpscbe2 = 6.484591271e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 6.485633595e+00 lbeta0 = 1.251387297e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.075221224e-09 lagidl = -6.001562308e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.178852899e-01 lkt1 = -6.473825875e-8
+ kt2 = -6.397594635e-02 lkt2 = 1.631355860e-8
+ at = 8.764820671e+04 lat = -2.739227930e-2
+ ute = -1.993146628e+00 lute = 9.999567120e-7
+ ua1 = -3.697989286e-09 lua1 = 3.457660733e-15 wua1 = 3.308722450e-30 pua1 = 3.308722450e-36
+ ub1 = 4.480108576e-18 lub1 = -3.793775449e-24 wub1 = -3.081487911e-39 pub1 = 1.540743956e-45
+ uc1 = 3.486000352e-10 luc1 = -2.980666517e-16 wuc1 = -2.067951531e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.132 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 7.5e-07 wmax = 7.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.098276299e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.396542597e-9
+ k1 = 4.257803294e-01 lk1 = 4.686759479e-8
+ k2 = 3.182319986e-02 lk2 = -2.156085776e-08 pk2 = 2.081668171e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.533005469e-01 ldsub = 3.198469920e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.483210014e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.258875430e-8
+ nfactor = {2.949899408e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.859852442e-07 wnfactor = -7.105427358e-21
+ eta0 = 4.065893232e-01 leta0 = 2.570466844e-8
+ etab = -1.371832211e-03 letab = 4.006295315e-10 wetab = -3.469446952e-24
+ u0 = 7.628780961e-03 lu0 = -7.032655101e-10
+ ua = -1.951245750e-09 lua = 4.189831196e-16
+ ub = 2.631040349e-18 lub = -7.785751474e-25
+ uc = -6.837589508e-11 luc = 2.076637300e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.179337001e+05 lvsat = 1.691748002e-2
+ a0 = 9.109963816e-01 la0 = -9.135116129e-8
+ ags = 9.336688756e-01 lags = 1.765665437e-7
+ a1 = 0.0
+ a2 = 1.143114794e+00 la2 = -1.069636043e-7
+ b0 = -1.271017328e-15 lb0 = 7.583993833e-22 wb0 = 7.888609052e-37 pb0 = -2.958228395e-43
+ b1 = 3.942634583e-18 lb1 = -2.180307244e-24 wb1 = -1.925929944e-39 pb1 = 8.185202264e-46
+ keta = -4.608909199e-02 lketa = 4.420916754e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.532423753e-01 lpclm = 3.976759966e-07 wpclm = 2.220446049e-22 ppclm = 3.885780586e-28
+ pdiblc1 = -4.640274633e-01 lpdiblc1 = 2.676941088e-07 wpdiblc1 = -2.775557562e-22 ppdiblc1 = -1.387778781e-28
+ pdiblc2 = -1.035031450e-02 lpdiblc2 = 5.832680064e-09 wpdiblc2 = -6.071532166e-24 ppdiblc2 = -3.035766083e-30
+ pdiblcb = 2.758644106e-01 lpdiblcb = -1.737722132e-07 wpdiblcb = -1.110223025e-22 ppdiblcb = 1.665334537e-28
+ drout = 1.496502075e+00 ldrout = -2.982533618e-7
+ pscbe1 = 6.854817729e+08 lpscbe1 = 3.528285254e+1
+ pscbe2 = 2.184228811e-08 lpscbe2 = -4.005460978e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.502780999e+00 lbeta0 = 1.254761302e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.261721264e-12 lagidl = -1.262424958e-18
+ bgidl = 7.033052157e+08 lbgidl = 1.656061277e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.00081386752815302
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207367379934e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.477070908e-01 lkt1 = 7.724375894e-9
+ kt2 = -1.248182315e-02 lkt2 = -1.242891616e-8
+ at = 2.437475586e+03 lat = 2.016979449e-2
+ ute = 5.785487810e-01 lute = -4.354865146e-07 pute = 4.440892099e-28
+ ua1 = 5.210530986e-09 lua1 = -1.514808027e-15
+ ub1 = -4.963733815e-18 lub1 = 1.477494058e-24
+ uc1 = -2.932921455e-10 luc1 = 6.021830677e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.133 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7.5e-07 wmax = 7.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.051933961e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.884775766e-9
+ k1 = -1.224831150e+00 lk1 = 5.555365344e-7
+ k2 = 6.354475517e-01 lk2 = -2.075797743e-07 wk2 = -2.220446049e-22 pk2 = -5.551115123e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.367422949e+00 ldsub = -4.877813677e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.035820758e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.201544042e-8
+ nfactor = {-1.810663453e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.286651779e-7
+ eta0 = 1.340861129e+00 leta0 = -2.622098740e-7
+ etab = 8.580783120e-02 letab = -2.646552734e-08 wetab = -6.201636427e-23 petab = -1.637145280e-29
+ u0 = 5.307966851e-03 lu0 = 1.193977425e-11
+ ua = 6.737004918e-10 lua = -3.899465637e-16
+ ub = -1.794844881e-18 lub = 5.853499039e-25 wub = -7.703719778e-40 pub = -1.925929944e-46
+ uc = -1.109713200e-12 luc = 3.695372767e-20
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -4.056284828e+05 lvsat = 1.782636380e-1
+ a0 = -1.084521995e+00 la0 = 5.236077367e-7
+ ags = 2.379753985e+00 lags = -2.690735046e-7
+ a1 = 0.0
+ a2 = 1.281859579e+00 la2 = -1.497205848e-7
+ b0 = 5.036955310e-07 lb0 = -1.552238514e-13 wb0 = 3.989876326e-28 pb0 = 8.147784885e-35
+ b1 = -1.545339850e-14 lb1 = 4.761308510e-21 wb1 = 2.465190329e-38 pb1 = -3.112302790e-42
+ keta = -1.389542671e-01 lketa = 3.303917776e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.890048734e-01 lpclm = -1.596433800e-8
+ pdiblc1 = 1.161240433e+00 lpdiblc1 = -2.331646988e-7
+ pdiblc2 = 2.531901467e-02 lpdiblc2 = -5.159537107e-9
+ pdiblcb = 2.242036531e-01 lpdiblcb = -1.578519175e-7
+ drout = -1.074947880e+00 ldrout = 4.941903708e-7
+ pscbe1 = 7.998824353e+08 lpscbe1 = 2.800039958e-2
+ pscbe2 = 1.442103334e-08 lpscbe2 = -1.718452894e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.080950965e+01 lbeta0 = -5.853884369e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.697791983e-12 lagidl = 2.659482394e-19
+ bgidl = 2.059624081e+09 lbgidl = -2.523706569e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.00081386752815302
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207367379934e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.633079613e-01 lkt1 = -1.828490384e-8
+ kt2 = 8.301188984e-02 lkt2 = -4.185721369e-8
+ at = 1.645520113e+05 lat = -2.978904198e-2
+ ute = -3.389799098e+00 lute = 7.874392514e-7
+ ua1 = -1.127266161e-09 lua1 = 4.383109196e-16
+ ub1 = 7.679260506e-19 lub1 = -2.888315626e-25
+ uc1 = -3.543481429e-10 luc1 = 7.903393350e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.134 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7.5e-07 wmax = 7.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -3.7585e-8
+ vth0 = {-8.731429556e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -5.406967295e-08 wvth0 = -1.280013233e-07 pvth0 = 3.266209767e-14
+ k1 = 2.605390056e-01 lk1 = 2.161674894e-07 wk1 = 6.245073117e-07 pk1 = -1.593555307e-13
+ k2 = 5.406176255e-02 lk2 = -7.404410594e-08 wk2 = -1.481131749e-07 pk2 = 3.779403883e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 3.016733186e+00 ldsub = -6.882825181e-07 wdsub = -1.988448817e-06 pdsub = 5.073924846e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {1.580472458e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -4.533070449e-07 wvoff = -1.309134937e-06 pvoff = 3.340519618e-13
+ nfactor = {-1.832633458e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.130972790e-06 wnfactor = 1.481806846e-05 pnfactor = -3.781126529e-12
+ eta0 = 6.047314715e+00 leta0 = -1.481871544e-06 weta0 = -4.279592707e-06 peta0 = 1.092023671e-12
+ etab = 5.504334317e-01 letab = -1.469130873e-07 wetab = -4.244319042e-07 petab = 1.083022890e-13
+ u0 = -3.977912834e-02 lu0 = 1.151766609e-08 wu0 = 3.399341013e-08 pu0 = -8.674098463e-15
+ ua = -1.624724534e-08 lua = 3.899937740e-15 wua = 1.126278530e-14 pua = -2.873924926e-21
+ ub = 6.695224152e-18 lub = -1.539280147e-24 wub = -4.445382822e-24 pub = 1.134328335e-30
+ uc = -2.922989648e-10 luc = 7.434235273e-17 wuc = 2.147749398e-16 puc = -5.480412139e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -6.122296385e+06 lvsat = 1.649709815e+00 wvsat = 4.312130508e+00 pvsat = -1.100326342e-6
+ a0 = -4.385412326e+00 la0 = 1.403269780e-06 wa0 = 4.052593808e-06 pa0 = -1.034100362e-12
+ ags = 1.250000075e+00 lags = -1.689230800e-14
+ a1 = 0.0
+ a2 = 2.900205602e+00 la2 = -5.733606335e-07 wa2 = -1.656437914e-06 pa2 = 4.226732626e-13
+ b0 = 4.386162231e-06 lb0 = -1.156992383e-12 wb0 = -3.102498563e-12 pb0 = 7.916645583e-19
+ b1 = -1.008426163e-13 lb1 = 2.688992593e-20 wb1 = 7.765712257e-20 pb1 = -1.981576797e-26
+ keta = -2.863984220e-01 lketa = 7.302075956e-08 wketa = 2.108815109e-07 pketa = -5.381063514e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.936426636e-01 lpclm = 7.229741149e-09 wpclm = 2.088664405e-08 ppclm = -5.329644961e-15
+ pdiblc1 = 4.249935502e+00 lpdiblc1 = -1.037949753e-06 wpdiblc1 = -2.998635163e-06 ppdiblc1 = 7.651617346e-13
+ pdiblc2 = -5.327312534e-02 lpdiblc2 = 1.452654395e-08 wpdiblc2 = 4.196714872e-08 ppdiblc2 = -1.070875734e-14
+ pdiblcb = -1.692654876e+01 lpdiblcb = 4.207238487e-06 wpdiblcb = 1.215470440e-05 ppdiblcb = -3.101515922e-12
+ drout = 1.000001229e+00 ldrout = -2.768534912e-13 wdrout = -8.526512829e-20 pdrout = 2.131628207e-26
+ pscbe1 = 8.000000009e+08 lpscbe1 = -2.132301331e-7
+ pscbe2 = -4.107526127e-08 lpscbe2 = 1.231987758e-14 wpscbe2 = 3.559210371e-14 ppscbe2 = -9.082037103e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.405681055e+00 lbeta0 = -1.378710959e-08 wbeta0 = -3.983301712e-08 pbeta0 = 1.016419098e-14
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.990456390e-10 lagidl = 5.038701111e-17 wagidl = 1.501310290e-16 pagidl = -3.830893466e-23
+ bgidl = 1.000000370e+09 lbgidl = -8.328956985e-5
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -2.8385e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.622475620e+00 lkt1 = 2.761947753e-07 wkt1 = 7.976408186e-07 pkt1 = -2.035340077e-13
+ kt2 = 8.946023622e-01 lkt2 = -2.519384215e-07 wkt2 = -7.278497097e-07 pkt2 = 1.857254104e-13
+ at = -4.594557899e+05 lat = 1.273127587e-01 wat = 3.678063572e-01 pat = -9.385314816e-8
+ ute = -9.490562993e+00 lute = 2.400376689e-06 wute = 6.934684027e-06 pute = -1.769523323e-12
+ ua1 = -7.833005889e-09 lua1 = 2.180700102e-15 wua1 = 6.300038390e-15 pua1 = -1.607580796e-21
+ ub1 = 7.344163149e-18 lub1 = -1.987506083e-24 wub1 = -5.741902368e-24 pub1 = 1.465161227e-30
+ uc1 = -1.823577597e-10 luc1 = 4.078839892e-17 wuc1 = 1.178376083e-16 puc1 = -3.006862252e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.135 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 7.0e-07 wmax = 7.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.143603+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43165561
+ k2 = 0.046387026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
+ voff = {-0.16725342+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.5720692+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.00827017
+ ua = -7.4124916e-10
+ ub = 6.3364395e-19
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = 5.7286e-9
+ b1 = 3.5674e-8
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.136 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 7.0e-07 wmax = 7.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.452847595e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.202880665e-06 wvth0 = 1.954377014e-07 pvth0 = -3.920122638e-12
+ k1 = 4.706663295e-01 lk1 = -7.824836434e-07 wk1 = -3.312090106e-08 pk1 = 6.643446641e-13
+ k2 = 4.866593871e-02 lk2 = -4.571081856e-08 wk2 = 1.045958004e-08 pk2 = -2.098000345e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.172472591e-06 lcit = 1.303205335e-10 pcit = -3.388131789e-32
+ voff = {-3.363084542e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.390934615e-06 wvoff = 1.244369106e-07 pvoff = -2.495976707e-12
+ nfactor = {4.298984170e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.290985573e-05 wnfactor = 7.351417379e-07 pnfactor = -1.474559795e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.475904365e-02 lu0 = -1.301549309e-07 wu0 = -4.804051062e-09 pu0 = 9.636047289e-14
+ ua = -1.115353601e-09 lua = 7.503850467e-15 wua = 2.421680589e-16 pua = -4.857448095e-21
+ ub = 1.482786469e-18 lub = -1.703224500e-23 wub = -7.614377418e-25 pub = 1.527304767e-29
+ uc = -4.216885731e-10 luc = 6.338894870e-15 wuc = 1.955886149e-16 puc = -3.923149687e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -7.959650191e+05 lvsat = 1.757338434e+01 wvsat = 5.484076081e-01 pvsat = -1.100005303e-5
+ a0 = 2.002085880e+00 la0 = -1.079301806e-05 wa0 = -2.312561031e-07 pa0 = 4.638574230e-12
+ ags = -1.672674376e+00 lags = 3.582317707e-05 wags = 1.101462242e-06 pags = -2.209331691e-11
+ a1 = 0.0
+ a2 = 1.084157408e+00 la2 = -2.289788703e-06 wa2 = 1.776356839e-21
+ b0 = -1.199766986e-06 lb0 = 2.418003539e-11 wb0 = 8.065370665e-13 pb0 = -1.617765759e-17
+ b1 = 9.274897472e-08 lb1 = -1.144819546e-12 wb1 = -2.208804204e-14 pb1 = 4.430457022e-19
+ keta = 1.148779199e-01 lketa = -1.835656743e-06 wketa = -4.973462692e-08 pketa = 9.975856016e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.958323949e-02 lpclm = 1.696584997e-06 ppclm = -6.661338148e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 2.019180054e-03 lpdiblc2 = -1.488358846e-08 wpdiblc2 = -6.589467512e-11 ppdiblc2 = 1.321726596e-15
+ pdiblcb = -8.509159751e-01 lpdiblcb = 1.255472903e-05 wpdiblcb = 3.861413352e-07 ppdiblcb = -7.745288545e-12
+ drout = 0.56
+ pscbe1 = 8.004366514e+08 lpscbe1 = -8.758427647e+00 wpscbe1 = -2.693798438e-01 ppscbe1 = 5.403266701e-6
+ pscbe2 = 6.644581452e-08 lpscbe2 = -1.130983717e-12 wpscbe2 = -3.552867723e-14 ppscbe2 = 7.126402478e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.715141667e-11 lalpha0 = 1.346934531e-15
+ alpha1 = -6.715141667e-11 lalpha1 = 1.346934531e-15
+ beta0 = 1.876471741e+01 lbeta0 = 2.253592082e-04 wbeta0 = 1.811663330e-05 pbeta0 = -3.633865106e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 3.636609780e-09 lagidl = -3.482805122e-14 wagidl = -5.063218785e-16 pagidl = 1.015589031e-20
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = -6.935234359e+00 legidl = 1.411139268e-04 wegidl = 4.340190851e-06 pegidl = -8.705628592e-11
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.395611516e-01 lkt1 = -1.979517698e-06 wkt1 = -6.468851651e-08 pkt1 = 1.297533261e-12
+ kt2 = -3.122222552e-02 lkt2 = -5.480649136e-07 wkt2 = -2.099389571e-08 pkt2 = 4.210991292e-13
+ at = 6.303838371e+05 lat = -1.122041668e+01 wat = -3.412793575e-01 pat = 6.845439371e-6
+ ute = -7.638463290e+00 lute = 1.515491683e-04 wute = 5.060990696e-06 pute = -1.015142117e-10
+ ua1 = -1.639833935e-08 lua1 = 3.708462654e-13 wua1 = 1.245020198e-14 pua1 = -2.497282679e-19
+ ub1 = 1.177257624e-17 lub1 = -2.607858206e-22 wub1 = -8.900721318e-24 pub1 = 1.785321813e-28
+ uc1 = 5.831329189e-10 luc1 = -1.229409205e-14 wuc1 = -4.181883290e-16 puc1 = 8.388092596e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.137 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 7.0e-07 wmax = 7.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-7.323783409e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.972169331e-07 wvth0 = -2.580522832e-07 pvth0 = -2.658232497e-13
+ k1 = 3.974239423e-01 lk1 = -1.922840360e-07 wk1 = 3.889433838e-08 pk1 = 8.403362203e-14
+ k2 = 5.514245814e-02 lk2 = -9.789971315e-08 wk2 = -2.519484722e-08 pk2 = 7.750940161e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {3.752401916e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.342845335e-06 wvoff = -3.747522576e-07 pvoff = 1.526574473e-12
+ nfactor = {1.527342211e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -9.670178160e-05 wnfactor = -8.907037677e-06 pnfactor = 6.295272294e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 7.878270188e-03 lu0 = -7.470848854e-08 wu0 = 8.875652582e-10 pu0 = 5.049646100e-14
+ ua = 1.346836232e-09 lua = -1.233689378e-14 wua = -1.412735427e-15 pua = 8.478045525e-21
+ ub = -6.211156914e-19 lub = -7.864372655e-26 wub = 1.173966407e-24 pub = -3.227679797e-31
+ uc = 3.755222512e-10 luc = -8.516547800e-17 wuc = -2.976820928e-16 puc = 5.170953101e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.801505774e+06 lvsat = -1.141564687e+01 wvsat = -1.689159759e+00 pvsat = 7.030645196e-6
+ a0 = 2.896423090e+00 la0 = -1.799973934e-05 wa0 = -1.065834917e-06 pa0 = 1.136375219e-11
+ ags = 3.467134723e+00 lags = -5.594278418e-06 wags = -2.111701793e-06 pags = 3.798905127e-12
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 1.407607172e-06 lb0 = 3.169371178e-12 wb0 = -9.387641901e-13 pb0 = -2.113723365e-18
+ b1 = -1.117269189e-07 lb1 = 5.028819662e-13 wb1 = 7.451314022e-14 pb1 = -3.353830467e-19
+ keta = -1.041186394e-01 lketa = -7.094523796e-08 wketa = 6.888709684e-08 pketa = 4.171158586e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 8.351120709e+00 lpclm = -6.615887894e-05 wpclm = -5.408436214e-06 ppclm = 4.358209844e-11
+ pdiblc1 = 0.39
+ pdiblc2 = -2.169026521e-02 lpdiblc2 = 1.761711521e-07 wpdiblc2 = 1.352371673e-08 ppdiblc2 = -1.081856724e-13
+ pdiblcb = -5.613065166e-01 lpdiblcb = 1.022100678e-05 wpdiblcb = 2.074748888e-07 ppdiblcb = -6.305563947e-12
+ drout = 0.56
+ pscbe1 = 6.547428104e+09 lpscbe1 = -4.631899254e+04 wpscbe1 = -3.545714841e+03 ppscbe1 = 2.857520551e-2
+ pscbe2 = -4.117572346e-07 lpscbe2 = 2.722457748e-12 wpscbe2 = 2.630654563e-13 ppscbe2 = -1.693482041e-18
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.151787176e-09 lalpha0 = 1.008711387e-14 walpha0 = 8.348444072e-16 palpha0 = -6.727318157e-21
+ alpha1 = -1.151787176e-09 lalpha1 = 1.008711387e-14 walpha1 = 8.348444072e-16 palpha1 = -6.727318157e-21
+ beta0 = 3.463851530e+02 lbeta0 = -2.414661957e-03 wbeta0 = -2.287409822e-04 pbeta0 = 1.625834121e-9
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.702958287e-10 lagidl = -1.092498913e-14 wagidl = 1.585407687e-17 pagidl = 5.948107695e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 2.120570308e+01 legidl = -8.565053105e-05 wegidl = -1.302057255e-05 pegidl = 5.283969692e-11
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.089950963e-01 lkt1 = -2.225824168e-06 wkt1 = -6.456924785e-08 pkt1 = 1.296572174e-12
+ kt2 = -1.708975935e-01 lkt2 = 5.774629462e-07 wkt2 = 8.172394408e-08 pkt2 = -4.066186859e-13
+ at = -1.498054465e+06 lat = 5.930900995e+00 wat = 9.377322204e-01 pat = -3.461053356e-6
+ ute = 2.156200438e+01 lute = -8.375316433e-05 wute = -1.449021820e-05 pute = 5.603275323e-11
+ ua1 = 4.432652987e-08 lua1 = -1.184850541e-13 wua1 = -2.918916703e-14 pua1 = 8.580884625e-20
+ ub1 = -2.520825029e-17 lub1 = 3.721196633e-23 wub1 = 1.737027317e-23 pub1 = -3.316395834e-29
+ uc1 = -7.053281763e-09 luc1 = 4.924143565e-14 wuc1 = 4.696203542e-15 puc1 = -3.282454655e-20
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.138 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 7.0e-07 wmax = 7.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-6.307830655e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.507396575e-08 wvth0 = -3.238180263e-07 pvth0 = 1.065316062e-15
+ k1 = 1.165578175e+00 lk1 = -3.309584499e-06 wk1 = -4.819930321e-07 pk1 = 2.197883122e-12
+ k2 = -2.582624379e-01 lk2 = 1.173950634e-06 wk2 = 1.866739899e-07 pk2 = -7.822903571e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.508951855e-01 ldsub = -1.180502115e-06 wdsub = 1.099990691e-08 pdsub = -4.463949222e-14
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.553313680e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.161212505e-07 wvoff = 3.181316759e-08 pvoff = -1.233371390e-13
+ nfactor = {-1.673578421e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.319701922e-05 wnfactor = 1.170871187e-05 pnfactor = -2.070949339e-11
+ eta0 = 1.618122575e-01 leta0 = -3.320080490e-7
+ etab = -1.415385492e-01 letab = 2.903155940e-07 wetab = 1.057506178e-11 petab = -4.291539845e-17
+ u0 = -3.059207770e-02 lu0 = 8.141072313e-08 wu0 = 2.637934827e-08 pu0 = -5.295352806e-14
+ ua = -8.165784812e-09 lua = 2.626693956e-14 wua = 4.866617420e-15 pua = -1.700463582e-20
+ ub = 5.127087384e-18 lub = -2.340582900e-23 wub = -2.655088477e-24 pub = 1.521618768e-29
+ uc = 6.474875467e-10 luc = -1.188846881e-15 wuc = -4.822785855e-16 puc = 8.008334801e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -3.276084994e+05 lvsat = 1.282830794e+00 wvsat = 2.541282935e-01 pvsat = -8.555480787e-7
+ a0 = -3.187982892e+00 la0 = 6.691814487e-06 wa0 = 2.832256348e-06 pa0 = -4.455364836e-12
+ ags = 2.861238532e+00 lags = -3.135448671e-06 wags = -1.794905420e-06 pags = 2.513291593e-12
+ a1 = 0.0
+ a2 = 0.8
+ b0 = 2.724418696e-06 lb0 = -2.174473846e-12 wb0 = -1.816974766e-12 pb0 = 1.450204446e-18
+ b1 = 2.005556412e-08 lb1 = -3.191375300e-14 wb1 = -1.337549693e-14 pb1 = 2.128398398e-20
+ keta = -1.949412298e-01 lketa = 2.976282734e-07 wketa = 1.345060579e-07 pketa = -2.245813135e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -1.501163856e+01 lpclm = 2.865116986e-05 wpclm = 9.633975288e-06 ppclm = -1.746256464e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 4.377545778e-02 lpdiblc2 = -8.949988100e-08 wpdiblc2 = -2.674795551e-08 ppdiblc2 = 5.524361978e-14
+ pdiblcb = 3.997291884e+00 lpdiblcb = -8.278560486e-06 wpdiblcb = -2.731797789e-06 ppdiblcb = 5.622504255e-12
+ drout = 0.56
+ pscbe1 = -1.059096579e+10 lpscbe1 = 2.323152342e+04 wpscbe1 = 7.027337398e+03 ppscbe1 = -1.433203789e-2
+ pscbe2 = 5.175719873e-07 lpscbe2 = -1.048918221e-12 wpscbe2 = -3.139306311e-13 ppscbe2 = 6.480661705e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.603574353e-09 lalpha0 = -5.152781626e-15 walpha0 = -1.669688814e-15 palpha0 = 3.436503427e-21
+ alpha1 = 2.603574353e-09 lalpha1 = -5.152781626e-15 walpha1 = -1.669688814e-15 palpha1 = 3.436503427e-21
+ beta0 = -5.267956115e+02 lbeta0 = 1.128854026e-03 wbeta0 = 3.590105547e-04 pbeta0 = -7.593615334e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 4.618749036e-09 lagidl = -2.694848348e-14 wagidl = -2.899534837e-15 pagidl = 1.777925152e-20
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.053539139e+00 lkt1 = 7.956621305e-07 wkt1 = 3.813564122e-07 pkt1 = -5.130699617e-13
+ kt2 = -2.412218004e-02 lkt2 = -1.817663334e-08 wkt2 = -2.416417518e-08 pkt2 = 2.309330303e-14
+ at = -6.528240797e+05 lat = 2.500812401e+00 wat = 5.037382524e-01 pat = -1.699832055e-6
+ ute = -6.677563222e-01 lute = 6.458983670e-06 wute = 3.564419442e-07 pute = -4.217517561e-12
+ ua1 = 8.602136075e-09 lua1 = 2.649060912e-14 wua1 = -3.517400301e-15 pua1 = -1.837154732e-20
+ ub1 = -1.438177108e-17 lub1 = -6.723726813e-24 wub1 = 7.689109630e-24 pub1 = 6.123849107e-30
+ uc1 = 1.116758930e-08 luc1 = -2.470195668e-14 wuc1 = -7.435508037e-15 puc1 = 1.640800143e-20
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.139 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 7.0e-07 wmax = 7.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-6.368486973e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.589864392e-09 wvth0 = -3.269836720e-07 pvth0 = 7.580753117e-15
+ k1 = -1.563455235e+00 lk1 = 2.307230194e-06 wk1 = 1.276963039e-06 pk1 = -1.422347495e-12
+ k2 = 7.820085420e-01 lk2 = -9.671038889e-07 wk2 = -4.833948298e-07 pk2 = 5.968251856e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -6.998324879e+00 ldsub = 1.497452715e-05 wdsub = 4.477820314e-06 pdsub = -9.238115249e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.063693748e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -9.046785504e-08 wvoff = -5.829290477e-08 pvoff = 6.211647598e-14
+ nfactor = {-3.154547172e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.244524586e-06 wnfactor = 3.539462032e-06 pnfactor = -3.895788454e-12
+ eta0 = 3.293396790e+00 leta0 = -6.777341386e-06 weta0 = -2.351010162e-06 peta0 = 4.838778585e-12
+ etab = 1.163952993e+01 letab = -2.395712612e-05 wetab = -7.180502916e-06 petab = 1.477867454e-11
+ u0 = -3.040990412e-02 lu0 = 8.103577894e-08 wu0 = 2.677732825e-08 pu0 = -5.377263852e-14
+ ua = 1.712862072e-09 lua = 5.935004908e-15 wua = -1.200769088e-15 pua = -4.516922926e-21
+ ub = -1.198176999e-17 lub = 1.180710799e-23 wub = 8.070567145e-24 pub = -6.859034954e-30
+ uc = 4.883536647e-10 luc = -8.613222993e-16 wuc = -3.758924777e-16 puc = 5.818727845e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.162923705e+05 lvsat = -6.598776594e-01 wvsat = -3.711047298e-01 pvsat = 4.312877727e-7
+ a0 = 6.615588193e+00 la0 = -1.348560141e-05 wa0 = -3.447683782e-06 pa0 = 8.469819541e-12
+ ags = -8.108816771e-01 lags = 4.422398979e-06 wags = 6.496357080e-07 pags = -2.517989621e-12
+ a1 = 0.0
+ a2 = -2.022726268e+00 la2 = 5.809650522e-06 wa2 = 1.741401934e-06 pa2 = -3.584101219e-12
+ b0 = 4.406306160e-07 lb0 = 2.525950267e-12 wb0 = -2.938662517e-13 pb0 = -1.684611804e-18
+ b1 = 1.105321430e-08 lb1 = -1.338538667e-14 wb1 = -7.371631787e-15 pb1 = 8.927008848e-21
+ keta = 7.616438446e-02 lketa = -2.603531687e-07 wketa = -5.796495421e-08 pketa = 1.715567495e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -5.422912625e+00 lpclm = 8.915941795e-06 wpclm = 3.916114641e-06 ppclm = -5.694235391e-12
+ pdiblc1 = 5.270223172e+00 lpdiblc1 = -1.004432893e-05 wpdiblc1 = -3.007021583e-06 ppdiblc1 = 6.188961612e-12
+ pdiblc2 = 1.424398499e-04 lpdiblc2 = 3.042875240e-10 wpdiblc2 = 1.917801904e-10 ppdiblc2 = -2.029360441e-16
+ pdiblcb = -2.636233411e+00 lpdiblcb = 5.374362269e-06 wpdiblcb = 1.741489009e-06 ppdiblcb = -3.584280433e-12
+ drout = -3.347651265e+00 ldrout = 8.042610604e-06 wdrout = 2.295583182e-06 pdrout = -4.724700437e-12
+ pscbe1 = 7.803138721e+08 lpscbe1 = -1.725032493e+02 wpscbe1 = 1.214480539e+01 ppscbe1 = 1.064210496e-4
+ pscbe2 = 6.535715718e-09 lpscbe2 = 2.881302063e-15 wpscbe2 = 2.001340972e-15 ppscbe2 = -2.175536358e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 2.087752126e+01 lbeta0 = 1.649614145e-06 wbeta0 = -1.003459611e-05 pbeta0 = 1.961246568e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -8.500506878e-09 lagidl = 5.317546391e-17 wagidl = 5.489484489e-15 pagidl = 5.132236169e-22
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -8.657685837e-01 lkt1 = 4.091984063e-07 wkt1 = 2.718263651e-07 pkt1 = -2.876385048e-13
+ kt2 = -1.644031208e-02 lkt2 = -3.398722352e-08 wkt2 = -2.664067740e-08 pkt2 = 2.819036561e-14
+ at = 9.612733707e+05 lat = -8.212745485e-01 wat = -5.759786458e-01 pat = 5.224088732e-7
+ ute = 6.193758896e+00 lute = -7.663181106e-06 wute = -3.483899445e-06 pute = 3.686557876e-12
+ ua1 = 4.465070811e-08 lua1 = -4.770348039e-14 wua1 = -2.561095510e-14 pua1 = 2.710074436e-20
+ ub1 = -3.779304433e-17 lub1 = 4.146065344e-23 wub1 = 2.229764168e-23 pub1 = -2.394299330e-29
+ uc1 = -1.787970850e-09 luc1 = 1.962788562e-15 wuc1 = 1.104461854e-15 puc1 = -1.168708400e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.140 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 7.0e-07 wmax = 7.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.397114219e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -5.286456151e-07 wvth0 = -6.768471182e-07 pvth0 = 3.777957560e-13
+ k1 = 7.366067346e-01 lk1 = -1.266263798e-07 wk1 = -1.422070319e-07 pk1 = 7.937569902e-14
+ k2 = -2.716156154e-01 lk2 = 1.478095858e-07 wk2 = 1.706225570e-07 pk2 = -9.523639265e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.478129496e+01 ldsub = -8.072013185e-06 wdsub = -8.999640255e-06 pdsub = 5.023329201e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.740163146e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.888589274e-08 wvoff = 8.653458885e-10 pvoff = -4.830101146e-16
+ nfactor = {1.491834592e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 3.278627939e-07 wnfactor = -3.008718316e-07 pnfactor = 1.679376302e-13
+ eta0 = -7.090036672e+00 leta0 = 4.210096400e-06 weta0 = 4.702020324e-06 peta0 = -2.624526684e-12
+ etab = -2.328031930e+01 letab = 1.299401074e-05 wetab = 1.436096353e-05 petab = -8.015859014e-12
+ u0 = 9.060407908e-02 lu0 = -4.701758766e-08 wu0 = -5.087534617e-08 pu0 = 2.839709197e-14
+ ua = 1.683529577e-08 lua = -1.006710076e-14 wua = -1.157508150e-14 pua = 6.460863243e-21
+ ub = -3.123268421e-18 lub = 2.433307379e-24 wub = 3.361994164e-24 pub = -1.876564283e-30
+ uc = -6.543242032e-10 luc = 3.478251401e-16 wuc = 3.682292828e-16 puc = -2.055345388e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.809601903e+05 lvsat = 1.837510828e-01 wvsat = 7.719176154e-02 pvsat = -4.308612554e-8
+ a0 = -1.380464829e+01 la0 = 8.122480225e-06 wa0 = 9.643167987e-06 pa0 = -5.382527075e-12
+ ags = 5.733271630e+00 lags = -2.502427726e-06 wags = -3.661129209e-06 pags = 2.043532490e-12
+ a1 = 0.0
+ a2 = 6.276346975e+00 la2 = -2.972179811e-06 wa2 = -3.482803869e-06 pa2 = 1.943996636e-12
+ b0 = 5.984424731e-06 lb0 = -3.340326352e-12 wb0 = -3.991144511e-12 pb0 = 2.227737131e-18
+ b1 = -3.378413787e-09 lb1 = 1.885729224e-15 wb1 = 2.253138480e-15 pb1 = -1.257634305e-21
+ keta = -3.169073405e-01 lketa = 1.555835385e-07 wketa = 2.204399479e-07 pketa = -1.230429657e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.289045284e+00 lpclm = -3.477300706e-06 wpclm = -3.100640724e-06 ppclm = 1.730684633e-12
+ pdiblc1 = -8.952449544e+00 lpdiblc1 = 5.005676662e-06 wpdiblc1 = 6.014043167e-06 ppdiblc1 = -3.356858474e-12
+ pdiblc2 = 7.991361598e-04 lpdiblc2 = -3.906088102e-10
+ pdiblcb = 5.209144272e+00 lpdiblcb = -2.927381033e-06 wpdiblcb = -3.482978018e-06 ppdiblcb = 1.944093840e-12
+ drout = 7.926354527e+00 ldrout = -3.887204105e-06 wdrout = -4.591166364e-06 pdrout = 2.562651329e-12
+ pscbe1 = 4.706065341e+08 lpscbe1 = 1.552197646e+02 wpscbe1 = 2.385446366e+02 ppscbe1 = -1.331484598e-4
+ pscbe2 = 3.221902770e-09 lpscbe2 = 6.387879510e-15 wpscbe2 = -1.155547617e-16 ppscbe2 = 6.449920134e-23
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 3.774021483e+01 lbeta0 = -1.619398231e-05 wbeta0 = -2.084436782e-05 pbeta0 = 1.163470079e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.788361180e-08 lagidl = 9.982095598e-15 wagidl = 1.264406284e-14 pagidl = -7.057536554e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.178852899e-01 lkt1 = -6.473825875e-8
+ kt2 = -6.397594635e-02 lkt2 = 1.631355860e-8
+ at = 3.487715478e+05 lat = -1.731434946e-01 wat = -1.741489009e-01 pat = 9.720469201e-8
+ ute = -1.993146628e+00 lute = 9.999567120e-7
+ ua1 = -3.697989286e-09 lua1 = 3.457660733e-15 wua1 = -1.654361225e-30 pua1 = 8.271806126e-37
+ ub1 = 5.524601940e-18 lub1 = -4.376780310e-24 wub1 = -6.965956036e-25 pub1 = 3.888187680e-31
+ uc1 = 3.486000352e-10 luc1 = -2.980666517e-16 wuc1 = -2.067951531e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.141 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 7.0e-07 wmax = 7.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.098276299e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.396542597e-9
+ k1 = 4.257803294e-01 lk1 = 4.686759479e-8
+ k2 = 3.182319986e-02 lk2 = -2.156085776e-08 wk2 = 2.775557562e-23 pk2 = 1.387778781e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.533005469e-01 ldsub = 3.198469920e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.483210014e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.258875430e-8
+ nfactor = {2.949899408e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.859852442e-7
+ eta0 = 4.065893232e-01 leta0 = 2.570466844e-8
+ etab = -1.371832211e-03 letab = 4.006295315e-10
+ u0 = 7.628780961e-03 lu0 = -7.032655101e-10 wu0 = 1.387778781e-23
+ ua = -1.951245750e-09 lua = 4.189831196e-16
+ ub = 2.631040349e-18 lub = -7.785751474e-25
+ uc = -6.837589508e-11 luc = 2.076637300e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.179337001e+05 lvsat = 1.691748002e-2
+ a0 = 9.109963816e-01 la0 = -9.135116129e-8
+ ags = 9.336688756e-01 lags = 1.765665437e-7
+ a1 = 0.0
+ a2 = 1.143114794e+00 la2 = -1.069636043e-7
+ b0 = -1.271017328e-15 lb0 = 7.583993833e-22 wb0 = -3.944304526e-37 pb0 = -9.860761315e-44
+ b1 = 3.942634583e-18 lb1 = -2.180307244e-24 wb1 = -3.851859889e-40 pb1 = -2.648153674e-46
+ keta = -4.608909199e-02 lketa = 4.420916754e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.532423753e-01 lpclm = 3.976759966e-07 wpclm = 2.220446049e-22 ppclm = -2.220446049e-28
+ pdiblc1 = -4.640274633e-01 lpdiblc1 = 2.676941088e-07 wpdiblc1 = 1.110223025e-22 ppdiblc1 = -1.804112415e-28
+ pdiblc2 = -1.035031450e-02 lpdiblc2 = 5.832680064e-09 wpdiblc2 = -2.168404345e-25 ppdiblc2 = 5.421010862e-31
+ pdiblcb = 2.758644106e-01 lpdiblcb = -1.737722132e-07 wpdiblcb = -2.220446049e-22 ppdiblcb = -1.110223025e-28
+ drout = 1.496502075e+00 ldrout = -2.982533618e-7
+ pscbe1 = 6.854817729e+08 lpscbe1 = 3.528285254e+1
+ pscbe2 = 2.184228811e-08 lpscbe2 = -4.005460978e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.502780999e+00 lbeta0 = 1.254761302e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.261721264e-12 lagidl = -1.262424958e-18
+ bgidl = 7.033052157e+08 lbgidl = 1.656061277e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.00081386752815302
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207367379934e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.477070908e-01 lkt1 = 7.724375894e-9
+ kt2 = -1.248182315e-02 lkt2 = -1.242891616e-8
+ at = 2.437475586e+03 lat = 2.016979449e-2
+ ute = 5.785487810e-01 lute = -4.354865146e-07 pute = 2.220446049e-28
+ ua1 = 5.210530986e-09 lua1 = -1.514808027e-15
+ ub1 = -4.963733815e-18 lub1 = 1.477494058e-24
+ uc1 = -2.932921455e-10 luc1 = 6.021830677e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.142 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7.0e-07 wmax = 7.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {1.268406560e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -7.229441142e-07 wvth0 = -1.547486141e-06 pvth0 = 4.768888041e-13
+ k1 = -2.735775594e+00 lk1 = 1.021164284e-06 wk1 = 1.007682090e-06 pk1 = -3.105373898e-13
+ k2 = 2.494241474e+00 lk2 = -7.804042973e-07 wk2 = -1.239670560e-06 pk2 = 3.820292766e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 7.178321780e+00 ldsub = -1.970356061e-06 wdsub = -3.208494270e-06 pdsub = 9.887616793e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {3.107867034e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.011687712e-06 wvoff = -2.141786063e-06 pvoff = 6.600342110e-13
+ nfactor = {-3.636841564e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.163073990e-05 wnfactor = 2.424282078e-05 pnfactor = -7.470910080e-12
+ eta0 = 1.183916011e+01 leta0 = -3.497470671e-06 weta0 = -7.001546553e-06 peta0 = 2.157666601e-12
+ etab = 1.112686979e+00 letab = -3.429188742e-07 wetab = -6.848482947e-07 petab = 2.110496990e-13
+ u0 = -8.843026746e-02 lu0 = 2.889925144e-08 wu0 = 6.251609070e-08 pu0 = -1.926558367e-14
+ ua = -2.695314968e-08 lua = 8.123819854e-15 wua = 1.842495417e-14 pua = -5.678018127e-21
+ ub = 9.110366980e-18 lub = -2.775309235e-24 wub = -7.272925705e-24 pub = 2.241297514e-30
+ uc = -5.207398385e-10 luc = 1.601713694e-16 wuc = 3.465527624e-16 puc = -1.067971648e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.171198063e+07 lvsat = 3.662542178e+00 wvsat = 7.540454985e+00 pvsat = -2.323742013e-6
+ a0 = -1.102596120e+01 la0 = 3.587261058e-06 wa0 = 6.630164520e-06 pa0 = -2.043217800e-12
+ ags = 2.379753974e+00 lags = -2.690735012e-07 wags = 7.325915874e-15 pags = -2.257626974e-21
+ a1 = 0.0
+ a2 = 5.289473919e+00 la2 = -1.384747096e-06 wa2 = -2.672766171e-06 pa2 = 8.236663509e-13
+ b0 = 6.718513157e-06 lb0 = -2.070444199e-12 wb0 = -4.144798601e-12 pb0 = 1.277302585e-18
+ b1 = -2.059540609e-13 lb1 = 6.346789763e-20 wb1 = 1.270490828e-19 pb1 = -3.915271583e-26
+ keta = -6.562700810e-01 lketa = 1.924603921e-07 wketa = 3.450092973e-07 pketa = -1.063215151e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.384720155e-01 lpclm = -3.916271915e-10 wpclm = 3.370147463e-08 ppclm = -1.038578344e-14
+ pdiblc1 = 8.416192265e+00 lpdiblc1 = -2.468923205e-06 wpdiblc1 = -4.838486986e-06 ppdiblc1 = 1.491076534e-12
+ pdiblc2 = -7.621696804e-02 lpdiblc2 = 2.613080669e-08 wpdiblc2 = 6.771658067e-08 ppdiblc2 = -2.086821866e-14
+ pdiblcb = -2.918309026e+01 lpdiblcb = 8.904593847e-06 wpdiblcb = 1.961237127e-05 ppdiblcb = -6.043944454e-12
+ drout = -1.074952843e+00 ldrout = 4.941919004e-07 wdrout = 3.310101523e-12 pdrout = -1.020073984e-18
+ pscbe1 = 7.998824338e+08 lpscbe1 = 2.800085717e-02 wpscbe1 = 9.902839661e-07 ppscbe1 = -3.051767349e-13
+ pscbe2 = -7.169111669e-08 lpscbe2 = 2.481872838e-14 wpscbe2 = 5.743008732e-14 ppscbe2 = -1.769823001e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.090589208e+01 lbeta0 = -6.150906110e-07 wbeta0 = -6.427956436e-08 pbeta0 = 1.980903335e-14
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 4.352779938e-08 lagidl = -1.341452737e-14 wagidl = -2.903144623e-14 pagidl = 8.946620786e-21
+ bgidl = 2.059624075e+09 lbgidl = -2.523706552e+02 wbgidl = 3.675559998e-06 pbgidl = -1.132696152e-12
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.00081386752815302
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207367379934e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.420009438e+00 lkt1 = 5.847117903e-07 wkt1 = 1.304967262e-06 pkt1 = -4.021517613e-13
+ kt2 = 1.843982654e+00 lkt2 = -5.845355742e-07 wkt2 = -1.174430144e-06 pkt2 = 3.619241375e-13
+ at = -7.253247705e+05 lat = 2.444442859e-01 wat = 5.934784031e-01 pat = -1.828922395e-7
+ ute = -2.016769134e+01 lute = 5.957882304e-06 wute = 1.118954545e-05 pute = -3.448282222e-12
+ ua1 = -1.636967365e-08 lua1 = 5.135563635e-15 wua1 = 1.016549689e-14 pua1 = -3.132701176e-21
+ ub1 = 1.465998202e-17 lub1 = -4.569946451e-24 wub1 = -9.264917751e-24 pub1 = 2.855169703e-30
+ uc1 = -6.394463681e-10 luc1 = 1.668926536e-16 wuc1 = 1.901382786e-16 puc1 = -5.859491330e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.143 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7.0e-07 wmax = 7.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -3.7585e-8
+ vth0 = {-6.407328415e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.184071173e-06 wvth0 = 3.562868712e-06 pvth0 = -7.930812714e-13
+ k1 = 4.048980968e+00 lk1 = -6.372138054e-07 wk1 = -1.902087979e-06 pk1 = 4.097832291e-13
+ k2 = -4.400987363e+00 lk2 = 9.233478689e-07 wk2 = 2.823057098e-06 pk2 = -6.273886118e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -9.045795639e+00 ldsub = 2.028912719e-06 wdsub = 6.056317032e-06 pdsub = -1.304764798e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-6.447769205e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.354412159e-06 wvoff = 4.045076050e-06 pvoff = -8.715557448e-13
+ nfactor = {7.254511478e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.533055150e-05 wnfactor = -4.578610029e-05 pnfactor = 9.865114172e-12
+ eta0 = -2.019718424e+01 leta0 = 4.427602298e-06 weta0 = 1.322344103e-05 peta0 = -2.849134443e-12
+ etab = -2.024295281e+00 letab = 4.330681672e-07 wetab = 1.292711319e-06 petab = -2.784999692e-13
+ u0 = 1.751832401e-01 lu0 = -3.630424844e-08 wu0 = -1.093697226e-07 pu0 = 2.321938842e-14
+ ua = 5.281805625e-08 lua = -1.165154010e-14 wua = -3.479838377e-14 pua = 7.497697780e-21
+ ub = -2.056670330e-17 lub = 4.599293910e-24 wub = 1.373619636e-23 pub = -2.959621753e-30
+ uc = 1.010587176e-09 luc = -2.191446989e-16 wuc = -6.541484909e-16 puc = 1.409288501e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.481328213e+07 lvsat = -5.396185694e+00 wvsat = -1.631948738e+01 pvsat = 3.598736383e-6
+ a0 = 2.046700378e+01 la0 = -4.192748777e-06 wa0 = -1.252202924e-05 pa0 = 2.698007526e-12
+ ags = 1.250000102e+00 lags = -2.307554681e-14 wags = -1.831389795e-14 pags = 4.123741348e-21
+ a1 = 0.0
+ a2 = -7.148221011e+00 la2 = 1.690139612e-06 wa2 = 5.045078859e-06 pa2 = -1.086904848e-12
+ b0 = -1.354524638e-05 lb0 = 2.952476009e-12 wb0 = 8.856352328e-12 pb0 = -1.949030321e-18
+ b1 = 3.753865214e-13 lb1 = -8.034259334e-20 wb1 = -2.399505664e-19 pb1 = 5.169995825e-26
+ keta = 1.006829561e+00 lketa = -2.181753849e-07 wketa = -6.516006816e-07 pketa = 1.403944799e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 7.203454074e-01 lpclm = -2.131121400e-08 wpclm = -6.361420327e-08 ppclm = 1.370494593e-14
+ pdiblc1 = -1.394064992e+01 lpdiblc1 = 3.059646433e-06 wpdiblc1 = 9.133066448e-06 ppdiblc1 = -1.967615309e-12
+ pdiblc2 = 2.013114694e-01 lpdiblc2 = -4.282097075e-08 wpdiblc2 = -1.278209184e-07 ppdiblc2 = 2.753756186e-14
+ pdiblcb = 5.680735122e+01 lpdiblcb = -1.240199868e-05 wpdiblcb = -3.702005564e-05 ppdiblcb = 7.975549748e-12
+ drout = 1.000013637e+00 ldrout = -3.070658778e-12 wdrout = -8.274860022e-12 pdrout = 1.863250231e-18
+ pscbe1 = 8.000000046e+08 lpscbe1 = -1.049053192e-06 wpscbe1 = -2.475601196e-06 ppscbe1 = 5.574302673e-13
+ pscbe2 = 1.748366370e-07 lpscbe2 = -3.631625759e-14 wpscbe2 = -1.084042913e-13 ppscbe2 = 2.335447143e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.164018205e+00 lbeta0 = 4.064966148e-08 wbeta0 = 1.213372543e-07 pbeta0 = -2.614088926e-14
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.087874781e-07 lagidl = 2.449426539e-14 wagidl = 7.257014558e-14 pagidl = -1.634046919e-20
+ bgidl = 1.000000384e+09 lbgidl = -8.639182663e-05 wbgidl = -9.188446045e-06 pbgidl = 2.068965912e-12
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -2.8385e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 3.269044674e+00 lkt1 = -8.252288306e-07 wkt1 = -2.464621679e-06 pkt1 = 5.310296265e-13
+ kt2 = -3.520739043e+00 lkt2 = 7.426577223e-07 wkt2 = 2.216838611e-06 pkt2 = -4.775926390e-13
+ at = 1.771762283e+06 lat = -3.752895741e-01 wat = -1.120242062e+00 pat = 2.413434048e-7
+ ute = 3.257721216e+01 lute = -7.075775458e-06 wute = -2.112124071e-05 pute = 4.550331018e-12
+ ua1 = 3.038479664e-08 lua1 = -6.428210405e-15 wua1 = -1.918825491e-14 pua1 = 4.133891018e-21
+ ub1 = -2.748785737e-17 lub1 = 5.858725975e-24 wub1 = 1.748833842e-23 pub1 = -3.767663550e-30
+ uc1 = 5.324786376e-10 luc1 = -1.202350552e-16 wuc1 = -3.589025114e-16 puc1 = 7.732146153e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.144 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 6.4e-07 wmax = 7.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.143603+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43165561
+ k2 = 0.046387026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
+ voff = {-0.16725342+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.5720692+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.00827017
+ ua = -7.4124916e-10
+ ub = 6.3364395e-19
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = 5.7286e-9
+ b1 = 3.5674e-8
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.145 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 6.4e-07 wmax = 7.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.136052763e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.514439310e-7
+ k1 = 4.169789897e-01 lk1 = 2.943861458e-7
+ k2 = 6.562039979e-02 lk2 = -3.857862811e-7
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.172472591e-06 lcit = 1.303205335e-10 wcit = 1.270549421e-27 pcit = 5.421010862e-32
+ voff = {-1.346023867e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.549199771e-7
+ nfactor = {1.621526756e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -9.920280577e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 6.971914874e-03 lu0 = 2.604062203e-8
+ ua = -7.228111739e-10 lua = -3.698322591e-16
+ ub = 2.485336107e-19 lub = 7.724608655e-24
+ uc = -1.046491178e-10 luc = -2.033642163e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.297654578e+04 lvsat = -2.571566868e-1
+ a0 = 1.627231194e+00 la0 = -3.274119030e-6
+ ags = 1.127413528e-01 lags = 1.100485920e-8
+ a1 = 0.0
+ a2 = 1.084157408e+00 la2 = -2.289788703e-6
+ b0 = 1.075896438e-07 lb0 = -2.043146133e-12 wb0 = -3.308722450e-29 pb0 = 2.117582368e-34
+ b1 = 5.694535280e-08 lb1 = -4.266644107e-13
+ keta = 3.426055353e-02 lketa = -2.186199026e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.958323949e-02 lpclm = 1.696584997e-06 ppclm = -2.220446049e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 1.912368050e-03 lpdiblc2 = -1.274113513e-08 ppdiblc2 = 1.387778781e-29
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 8.855588799e-09 lpscbe2 = 2.417082098e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.715141667e-11 lalpha0 = 1.346934531e-15
+ alpha1 = -6.715141667e-11 lalpha1 = 1.346934531e-15
+ beta0 = 4.813088250e+01 lbeta0 = -3.636723234e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.815887098e-09 lagidl = -1.836585614e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.444180322e-01 lkt1 = 1.237194387e-7
+ kt2 = -6.525229044e-02 lkt2 = 1.345159137e-7
+ at = 7.718690531e+04 lat = -1.242985802e-1
+ ute = 5.651519091e-01 lute = -1.300034001e-05 wute = -2.220446049e-22 pute = -5.329070518e-27
+ ua1 = 3.782821288e-09 lua1 = -3.395088554e-14
+ ub1 = -2.655052084e-18 lub1 = 2.860600094e-23
+ uc1 = -9.472964564e-11 luc1 = 1.302590510e-15 puc1 = 8.271806126e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.146 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 6.4e-07 wmax = 7.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.150668308e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.366938589e-8
+ k1 = 4.604697380e-01 lk1 = -5.606969765e-8
+ k2 = 1.430285893e-02 lk2 = 2.773918708e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.322146530e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.316562590e-7
+ nfactor = {8.355552889e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.341463636e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 9.316969502e-03 lu0 = 7.143773174e-9
+ ua = -9.431379082e-10 lua = 1.405598021e-15
+ ub = 1.281825696e-18 lub = -6.018346318e-25
+ uc = -1.070056741e-10 luc = -1.346889891e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.346148460e+04 lvsat = -1.931930625e-2
+ a0 = 1.168757490e+00 la0 = 4.203400132e-7
+ ags = 4.417072978e-02 lags = 5.635585964e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = -1.140830747e-07 lb0 = -2.568696835e-13
+ b1 = 9.055190034e-09 lb1 = -4.075733774e-14
+ keta = 7.543931899e-03 lketa = -3.332823646e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -4.156864620e-01 lpclm = 4.485543601e-06 wpclm = -2.220446049e-22
+ pdiblc1 = 0.39
+ pdiblc2 = 2.310096564e-04 lpdiblc2 = 8.075366429e-10
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.465883797e-08 lpscbe2 = -2.259274738e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.014542500e-10 lalpha0 = -8.175355937e-16
+ alpha1 = 2.014542500e-10 lalpha1 = -8.175355937e-16
+ beta0 = -2.439264750e+01 lbeta0 = 2.207346103e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.959945019e-10 lagidl = -1.283401221e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.136586484e-01 lkt1 = -1.241449055e-7
+ kt2 = -3.842712868e-02 lkt2 = -8.164580001e-8
+ at = 2.196300907e+04 lat = 3.207049638e-1
+ ute = -1.925921477e+00 lute = 7.073152815e-6
+ ua1 = -2.987663864e-09 lua1 = 2.060683480e-14 pua1 = -6.617444900e-36
+ ub1 = 2.948102001e-18 lub1 = -1.654516721e-23
+ uc1 = 5.590315313e-10 luc1 = -3.965528193e-15 wuc1 = 2.067951531e-31 puc1 = -8.271806126e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.147 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 6.4e-07 wmax = 7.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.155676044e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.334714119e-8
+ k1 = 3.842913476e-01 lk1 = 2.530751608e-7
+ k2 = 4.432685200e-02 lk2 = -9.410328086e-08 wk2 = 2.775557562e-23
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.687254897e-01 ldsub = -1.252860521e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.037637994e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.619785835e-8
+ nfactor = {2.243457684e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.720436259e-7
+ eta0 = 1.618122575e-01 leta0 = -3.320080490e-7
+ etab = -1.415214075e-01 letab = 2.902460303e-7
+ u0 = 1.216753903e-02 lu0 = -4.424322556e-9
+ ua = -2.772390642e-10 lua = -1.296732691e-15
+ ub = 8.233204951e-19 lub = 1.258857421e-24
+ uc = -1.342621486e-10 luc = 1.092645171e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.432087493e+04 lvsat = -1.039702583e-1
+ a0 = 1.402964339e+00 la0 = -5.301111964e-7
+ ags = -4.821423619e-02 lags = 9.384724937e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = -2.208073870e-07 lb0 = 1.762357191e-13
+ b1 = -1.625453795e-09 lb1 = 2.586530631e-15
+ keta = 2.308642681e-02 lketa = -6.640691024e-08 pketa = -2.775557562e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.045581146e-01 lpclm = 3.452176679e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 4.183469811e-04 lpdiblc2 = 4.728993188e-11
+ pdiblcb = -4.308170000e-01 lpdiblcb = 8.352403749e-07 wpdiblcb = 4.440892099e-22
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 8.705986359e-09 lpscbe2 = 1.564936435e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.029085000e-10 lalpha0 = 4.176201874e-16
+ alpha1 = -1.029085000e-10 lalpha1 = 4.176201874e-16
+ beta0 = 5.514271247e+01 lbeta0 = -1.020334014e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -8.125329299e-11 lagidl = 1.870802463e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.353792873e-01 lkt1 = -3.599886016e-8
+ kt2 = -6.329111094e-02 lkt2 = 1.925646684e-8
+ at = 1.637106726e+05 lat = -2.545311518e-1
+ ute = -8.998158855e-02 lute = -3.774033634e-7
+ ua1 = 2.900604438e-09 lua1 = -3.288758976e-15
+ ub1 = -1.918105287e-18 lub1 = 3.202729218e-24
+ uc1 = -8.850008756e-10 luc1 = 1.894600800e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.148 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 6.4e-07 wmax = 7.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.166873031e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.698160864e-9
+ k1 = 5.064385921e-01 lk1 = 1.675366545e-9
+ k2 = -1.550530049e-03 lk2 = 3.201705484e-10
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.600000206e-01 ldsub = -2.177893776e-14
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.008592856e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.021987531e-8
+ nfactor = {2.582745438e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.070355502e-6
+ eta0 = -5.174742150e-01 leta0 = 1.066078990e-06 weta0 = -6.765421556e-23 peta0 = -9.627715292e-29
+ etab = 2.904247369e-04 letab = -1.626828481e-09 petab = 8.673617380e-31
+ u0 = 1.299481844e-02 lu0 = -6.127004236e-9
+ ua = -2.335251343e-10 lua = -1.386703390e-15
+ ub = 1.100219537e-18 lub = 6.889521208e-25
+ uc = -1.209494201e-10 luc = 8.186465865e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.474998785e+04 lvsat = 3.921845435e-2
+ a0 = 1.027063579e+00 la0 = 2.435564714e-7
+ ags = 2.421456228e-01 lags = 3.408625427e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = -3.571202000e-08 lb0 = -2.047220124e-13
+ b1 = -8.958356404e-10 lb1 = 1.084852434e-15 pb1 = -8.271806126e-37
+ keta = -1.779393475e-02 lketa = 1.773182353e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.249152049e-01 lpclm = -3.141316846e-7
+ pdiblc1 = 3.959901522e-01 lpdiblc1 = -1.232875161e-8
+ pdiblc2 = 4.533060379e-04 lpdiblc2 = -2.466175011e-11
+ pdiblcb = 1.866340000e-01 lpdiblcb = -4.355787498e-07 wpdiblcb = 5.551115123e-23 ppdiblcb = -5.551115123e-29
+ drout = 3.733753506e-01 ldrout = 3.841052546e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 9.779790288e-09 lpscbe2 = -6.451345974e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.611938067e+00 lbeta0 = 1.967522498e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 3.976755324e-10 lagidl = 8.850855221e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.251515120e-01 lkt1 = -5.704936050e-8
+ kt2 = -5.962353039e-02 lkt2 = 1.170796260e-8
+ at = 2.764051955e+04 lat = 2.552435502e-2
+ ute = 5.465304861e-01 lute = -1.687453420e-06 pute = 4.440892099e-28
+ ua1 = 3.136618649e-09 lua1 = -3.774516346e-15 pua1 = 3.308722450e-36
+ ub1 = -1.649671782e-18 lub1 = 2.650247432e-24 wub1 = 7.703719778e-40 pub1 = -7.703719778e-46
+ uc1 = 2.307099871e-12 luc1 = 6.837014368e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.149 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 6.4e-07 wmax = 7.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.701718888e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.756560016e-07 wvth0 = 2.867896520e-07 pvth0 = -3.034722060e-13
+ k1 = -2.689738389e-01 lk1 = 8.221935387e-07 wk1 = 4.781577466e-07 pk1 = -5.059721828e-13
+ k2 = 4.441753006e-01 lk2 = -4.713335317e-07 wk2 = -2.709646065e-07 pk2 = 2.867266176e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 7.242244383e+00 ldsub = -7.388401539e-06 wdsub = -4.348634092e-06 pdsub = 4.601594137e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {3.148845983e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.355248304e-07 wvoff = -3.007483831e-07 pvoff = 3.182429166e-13
+ nfactor = {-1.904042172e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 2.181063129e-05 wnfactor = 1.236592880e-05 pnfactor = -1.308525487e-11
+ eta0 = -4.073855518e+00 leta0 = 4.829334993e-06 weta0 = 2.841271814e-06 peta0 = -3.006548596e-12
+ etab = -5.493259536e-03 letab = 4.493292706e-09 wetab = 2.211302724e-09 petab = -2.339934204e-15
+ u0 = 1.723166120e-02 lu0 = -1.061030413e-08 wu0 = -5.610287385e-09 pu0 = 5.936637802e-15
+ ua = 5.028599774e-09 lua = -6.954926104e-15 wua = -4.291270995e-15 pua = 4.540894228e-21
+ ub = -9.048668152e-18 lub = 1.142820061e-23 wub = 7.017503617e-24 pub = -7.425711802e-30
+ uc = -2.352634358e-10 luc = 2.028283207e-16 wuc = 1.097014761e-16 puc = -1.160828109e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -5.672224092e+05 lvsat = 6.550441858e-01 wvsat = 3.154854222e-01 pvsat = -3.338372092e-7
+ a0 = 5.628911146e+00 la0 = -4.625980569e-06 wa0 = -2.345822367e-06 pa0 = 2.482278854e-12
+ ags = -2.012374466e-01 lags = 8.100372052e-07 wags = -3.776055024e-16 pags = 3.995701547e-22
+ a1 = 0.0
+ a2 = -4.128599006e+00 la2 = 5.215295610e-06 wa2 = 2.936236215e-06 pa2 = -3.107037076e-12
+ b0 = -1.333206905e-06 lb0 = 1.168248150e-12 wb0 = 5.232634338e-13 pb0 = -5.537016678e-19
+ b1 = -3.028966319e-08 lb1 = 3.218851893e-14 wb1 = 1.885528028e-14 pb1 = -1.995209194e-20
+ keta = -1.514859230e-02 lketa = 1.493260150e-08 wketa = 3.427833748e-08 pketa = -3.627230837e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.131002325e+00 lpclm = -4.764886892e-06 wpclm = -2.386218545e-06 ppclm = 2.525024878e-12
+ pdiblc1 = 1.358743952e+00 lpdiblc1 = -1.031085940e-06 wpdiblc1 = -3.471589477e-07 ppdiblc1 = 3.673531836e-13
+ pdiblc2 = 8.096992318e-03 lpdiblc2 = -8.112981261e-09 wpdiblc2 = -4.502208017e-09 ppdiblc2 = 4.764101457e-15
+ pdiblcb = -2.400581086e+00 lpdiblcb = 2.302134638e-06 wpdiblcb = 1.211628970e-06 ppdiblcb = -1.282109427e-12
+ drout = -4.180479008e+00 ldrout = 5.202857321e-06 wdrout = 2.877805594e-06 pdrout = -3.045207546e-12
+ pscbe1 = -5.467721479e+09 lpscbe1 = 6.632314837e+03 wpscbe1 = 3.902029831e+03 ppscbe1 = -4.129010906e-3
+ pscbe2 = 6.611049608e-07 lpscbe2 = -6.898578903e-13 wpscbe2 = -4.059780867e-13 ppscbe2 = 4.295938320e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.946226562e-01 lbeta0 = 5.795257146e-06 wbeta0 = 1.824796389e-06 pbeta0 = -1.930944795e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.207631967e-08 lagidl = -1.147290534e-14 wagidl = -5.838878003e-15 pagidl = 6.178525537e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 1.000891385e-01 lkt1 = -6.128432597e-07 wkt1 = -3.195498203e-07 pkt1 = 3.381380334e-13
+ kt2 = -3.208985282e-01 lkt2 = 2.881813270e-07 wkt2 = 1.585011930e-07 pkt2 = -1.677212074e-13
+ at = 4.957469138e+05 lat = -4.698117882e-01 wat = -2.648212376e-01 pat = 2.802258890e-7
+ ute = -2.375964054e+00 lute = 1.405042627e-06 wute = 2.361684920e-07 pute = -2.499064131e-13
+ ua1 = -1.230923051e-08 lua1 = 1.256981786e-14 wua1 = 5.312464159e-15 pua1 = -5.621490200e-21
+ ub1 = 1.942292642e-17 lub1 = -1.964814381e-23 wub1 = -9.270777740e-24 pub1 = 9.810058881e-30
+ uc1 = 1.571904803e-09 luc1 = -1.592531058e-15 wuc1 = -7.546836241e-16 puc1 = 7.985835705e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.150 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 6.4e-07 wmax = 7.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.685326626e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -2.801225540e-07 wvth0 = -5.735793039e-07 pvth0 = 1.767599341e-13
+ k1 = 1.975920369e+00 lk1 = -4.308390611e-07 wk1 = -9.563154933e-07 pk1 = 2.947077456e-13
+ k2 = -8.466172075e-01 lk2 = 2.491481226e-07 wk2 = 5.419292130e-07 pk2 = -1.670063256e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -1.435114142e+01 ldsub = 4.664378613e-06 wdsub = 8.697268185e-06 pdsub = -2.680237136e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.223317462e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.230534135e-07 wvoff = 6.014967663e-07 pvoff = -1.853632585e-13
+ nfactor = {4.303901536e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.284024811e-05 wnfactor = -2.473185759e-05 pnfactor = 7.621616554e-12
+ eta0 = 9.617711034e+00 leta0 = -2.812886709e-06 weta0 = -5.682543628e-06 peta0 = 1.751189470e-12
+ etab = 5.796992128e-03 letab = -1.808587065e-09 wetab = -4.422605448e-09 petab = 1.362914321e-15
+ u0 = -1.055921488e-02 lu0 = 4.901729168e-09 wu0 = 1.122057477e-08 pu0 = -3.457844527e-15
+ ua = -1.586312114e-08 lua = 4.706205758e-15 wua = 8.582541989e-15 pua = -2.644881965e-21
+ ub = 2.538109179e-17 lub = -7.789458499e-24 wub = -1.403500723e-23 pub = 4.325168179e-30
+ uc = 2.872654212e-10 luc = -8.883161144e-17 wuc = -2.194029521e-16 puc = 6.761340776e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.140706181e+06 lvsat = -2.982703154e-01 wvsat = -6.309708443e-01 pvsat = 1.944462851e-7
+ a0 = -6.693927312e+00 la0 = 2.252258173e-06 wa0 = 4.691644735e-06 pa0 = -1.445824158e-12
+ ags = 9.336688743e-01 lags = 1.765665441e-07 wags = 7.552092285e-16 pags = -2.327329440e-22
+ a1 = 0.0
+ a2 = 1.066210169e+01 la2 = -3.040429795e-06 wa2 = -5.872472431e-06 pa2 = 1.809719829e-12
+ b0 = 1.696368207e-06 lb0 = -5.227697899e-13 wb0 = -1.046526868e-12 pb0 = 3.225081848e-19
+ b1 = 6.112695052e-08 lb1 = -1.883749234e-14 wb1 = -3.771056057e-14 pb1 = 1.162126345e-20
+ keta = 6.503788185e-02 lketa = -2.982508278e-08 wketa = -6.855667496e-08 pketa = 2.112711052e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -8.389126474e+00 lpclm = 2.781643399e-06 wpclm = 4.772437090e-06 ppclm = -1.470721938e-12
+ pdiblc1 = -1.589482375e+00 lpdiblc1 = 6.145255490e-07 wpdiblc1 = 6.943178953e-07 ppdiblc1 = -2.139679458e-13
+ pdiblc2 = -2.494602682e-02 lpdiblc2 = 1.033064073e-08 wpdiblc2 = 9.004416034e-09 ppdiblc2 = -2.774890889e-15
+ pdiblcb = 4.203845483e+00 lpdiblcb = -1.384258140e-06 wpdiblcb = -2.423257939e-06 ppdiblcb = 7.467753991e-13
+ drout = 1.082606268e+01 ldrout = -3.173344054e-06 wdrout = -5.755611189e-06 pdrout = 1.773706700e-12
+ pscbe1 = 1.333547588e+10 lpscbe1 = -3.863065830e+03 wpscbe1 = -7.804059662e+03 ppscbe1 = 2.404977066e-3
+ pscbe2 = -1.294298445e-06 lpscbe2 = 4.015896288e-13 wpscbe2 = 8.119561734e-13 ppscbe2 = -2.502205340e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.441859009e+01 lbeta0 = -1.697598759e-06 wbeta0 = -3.649592778e-06 pbeta0 = 1.124695007e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.892680226e-08 lagidl = 5.832107221e-15 wagidl = 1.167775601e-14 pagidl = -3.598734069e-21
+ bgidl = 7.033052157e+08 lbgidl = 1.656061277e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.00081386752815302
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207367379934e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.583655948e+00 lkt1 = 3.269727351e-07 wkt1 = 6.390996406e-07 pkt1 = -1.969513363e-13
+ kt2 = 5.013633405e-01 lkt2 = -1.707805802e-07 wkt2 = -3.170023861e-07 pkt2 = 9.769062531e-14
+ at = -8.560867386e+05 lat = 2.847412016e-01 wat = 5.296424753e-01 pat = -1.632199216e-7
+ ute = 1.344183633e+00 lute = -6.714322068e-07 wute = -4.723369839e-07 pute = 1.455600883e-13
+ ua1 = 2.243301344e-08 lua1 = -6.822260444e-15 wua1 = -1.062492832e-14 pua1 = 3.274284160e-21
+ ub1 = -3.501867671e-17 lub1 = 1.073952581e-23 wub1 = 1.854155548e-23 pub1 = -5.713951152e-30
+ uc1 = -2.739901682e-09 luc1 = 8.141899675e-16 wuc1 = 1.509367248e-15 puc1 = -4.651417049e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.151 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.4e-07 wmax = 7.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.239991813e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.006901243e-8
+ k1 = -1.102372845e+00 lk1 = 5.177985587e-7
+ k2 = 4.847969085e-01 lk2 = -1.611537656e-07 wk2 = 1.110223025e-22 pk2 = -2.775557562e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.977511515e+00 ldsub = -3.676223612e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-3.638620714e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.819504583e-8
+ nfactor = {2.927995871e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.792352313e-7
+ eta0 = 4.900000008e-01 leta0 = -9.356160291e-17
+ etab = 2.581819860e-03 letab = -8.177674270e-10 wetab = -8.673617380e-25 petab = -4.336808690e-31
+ u0 = 1.290521855e-02 lu0 = -2.329305283e-9
+ ua = 2.912788267e-09 lua = -1.079966243e-15
+ ub = -2.678685290e-18 lub = 8.577230029e-25 wub = 3.851859889e-40 pub = -1.925929944e-46
+ uc = 4.100502134e-11 luc = -1.294154402e-17 wuc = 2.584939414e-32 puc = -6.462348536e-39
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.107233529e+05 lvsat = -1.041285073e-1
+ a0 = -2.787929715e-01 la0 = 2.753062236e-7
+ ags = 2.379753986e+00 lags = -2.690735049e-7
+ a1 = 0.0
+ a2 = 9.570523633e-01 la2 = -4.962474518e-8
+ b0 = -4.369331260e-14 lb0 = 1.383167812e-20 wb0 = -2.524354897e-35 pb0 = 6.310887242e-42
+ b1 = -1.379167911e-17 lb1 = 3.284876207e-24
+ keta = -9.702710173e-02 lketa = 2.011848322e-08 wketa = -1.110223025e-22
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.931004364e-01 lpclm = -1.722646764e-8
+ pdiblc1 = 5.732445572e-01 lpdiblc1 = -5.196200978e-8
+ pdiblc2 = 3.354825457e-02 lpdiblc2 = -7.695541966e-9
+ pdiblcb = 2.607591983e+00 lpdiblcb = -8.923406993e-07 wpdiblcb = -8.881784197e-22
+ drout = -1.074947477e+00 ldrout = 4.941902469e-7
+ pscbe1 = 7.998824354e+08 lpscbe1 = 2.800036250e-2
+ pscbe2 = 2.140020980e-08 lpscbe2 = -3.869225705e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.080169809e+01 lbeta0 = -5.829811493e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -3.530736764e-09 lagidl = 1.087501718e-15 wagidl = -5.428372770e-31 pagidl = -3.505824081e-37
+ bgidl = 2.059624081e+09 lbgidl = -2.523706570e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.00081386752815302
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207367379934e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.047221533e-01 lkt1 = -6.715629230e-8
+ kt2 = -5.971042874e-02 lkt2 = 2.125523229e-9
+ at = 2.366743202e+05 lat = -5.201497393e-02 pat = -5.820766091e-23
+ ute = -2.029992490e+00 lute = 3.683876490e-7
+ ua1 = 1.080932106e-10 lua1 = 5.761022195e-17
+ ub1 = -3.579906755e-19 lub1 = 5.814219486e-26
+ uc1 = -3.312416379e-10 luc1 = 7.191320187e-17 wuc1 = 4.135903063e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.152 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.4e-07 wmax = 7.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -3.7585e-8
+ vth0 = {3.059119475e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.043361410e-06 wvth0 = -2.277191254e-06 pvth0 = 5.810708922e-13
+ k1 = -1.724570507e-02 lk1 = 2.778658782e-07 wk1 = 6.064567129e-07 pk1 = -1.547495594e-13
+ k2 = 3.580484714e+00 lk2 = -9.625831898e-07 wk2 = -2.100888619e-06 pk2 = 5.360837488e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 3.901209382e+00 ldsub = -8.847323429e-07 wdsub = -1.930975199e-06 pdsub = 4.927269416e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {2.231141376e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.998181619e-07 wvoff = -1.309134824e-06 pvoff = 3.340519330e-13
+ nfactor = {-2.569123910e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.789328303e-06 wnfactor = 1.481806762e-05 pnfactor = -3.781126315e-12
+ eta0 = 8.174365791e+00 leta0 = -1.960819619e-06 weta0 = -4.279592363e-06 peta0 = 1.092023583e-12
+ etab = 7.392235300e-01 letab = -1.888450029e-07 wetab = -4.121642335e-07 petab = 1.051719475e-13
+ u0 = -5.059688435e-02 lu0 = 1.370826612e-08 wu0 = 2.991900338e-08 pu0 = -7.634432094e-15
+ ua = -2.184387129e-08 lua = 5.160105190e-15 wua = 1.126220189e-14 pua = -2.873776057e-21
+ ub = 8.905281889e-18 lub = -2.036935704e-24 wub = -4.445719689e-24 pub = 1.134414293e-30
+ uc = -3.878321234e-10 luc = 9.556109401e-17 wuc = 2.085671400e-16 puc = -5.322007711e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.754288622e+07 lvsat = 4.495178605e+00 wvsat = 9.810964703e+00 pvsat = -2.503463863e-6
+ a0 = -6.399638652e+00 la0 = 1.856813110e-06 wa0 = 4.052593536e-06 pa0 = -1.034100293e-12
+ ags = 1.250000072e+00 lags = -1.619899592e-14 wags = 4.646167895e-16 pags = -1.185558318e-22
+ a1 = 0.0
+ a2 = 3.636999024e+00 la2 = -7.370088291e-07 wa2 = -1.608560655e-06 pa2 = 4.104564224e-13
+ b0 = 8.333196256e-06 lb0 = -2.126381685e-12 wb0 = -4.640940257e-12 pb0 = 1.184228725e-18
+ b1 = -1.394394178e-13 lb1 = 3.558075637e-20 wb1 = 7.765688169e-20 pb1 = -1.981570650e-26
+ keta = -3.912113512e-01 lketa = 9.662148694e-08 wketa = 2.108815137e-07 pketa = -5.381063585e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 5.843522881e-01 lpclm = 9.293213645e-09 wpclm = 2.028294385e-08 ppclm = -5.175598783e-15
+ pdiblc1 = 5.583746724e+00 lpdiblc1 = -1.334200771e-06 wpdiblc1 = -2.911963379e-06 ppdiblc1 = 7.430456954e-13
+ pdiblc2 = -7.194035094e-02 lpdiblc2 = 1.867269628e-08 wpdiblc2 = 4.075414114e-08 ppdiblc2 = -1.039923419e-14
+ pdiblcb = -2.233303216e+01 lpdiblcb = 5.408065236e-06 wpdiblcb = 1.180338795e-05 ppdiblcb = -3.011870503e-12
+ drout = 1.000000254e+00 ldrout = -5.808437109e-14 wdrout = -1.852413334e-14 pdrout = 4.726803837e-21
+ pscbe1 = 8.000000019e+08 lpscbe1 = -4.826679230e-07 wpscbe1 = -8.151931763e-07 ppscbe1 = 2.080135345e-13
+ pscbe2 = -5.690684101e-08 lpscbe2 = 1.583620845e-14 wpscbe2 = 3.456335862e-14 ppscbe2 = -8.819532220e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 8.423401005e+00 lbeta0 = -1.772287036e-08 wbeta0 = -3.868170173e-08 pbeta0 = 9.870409829e-15
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 8.133594101e-08 lagidl = -2.049030520e-14 wagidl = -4.472117438e-14 pagidl = 1.141150207e-20
+ bgidl = 1.000000350e+09 lbgidl = -7.814711380e-05 wbgidl = 1.182498932e-05 pbgidl = -3.017381668e-12
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -2.8385e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.018922143e+00 lkt1 = 3.654626648e-07 wkt1 = 7.976413853e-07 pkt1 = -2.035341523e-13
+ kt2 = 1.218353969e+00 lkt2 = -3.238464545e-07 wkt2 = -7.068121285e-07 pkt2 = 1.803572508e-13
+ at = -6.230581952e+05 lat = 1.636502687e-01 wat = 3.571753766e-01 pat = -9.114044086e-8
+ ute = -1.257515134e+01 lute = 3.085490454e-06 wute = 6.734245681e-06 pute = -1.718377470e-12
+ ua1 = -1.063529764e-08 lua1 = 2.803113345e-15 wua1 = 6.117943697e-15 pua1 = -1.561115693e-21
+ ub1 = 9.898195170e-18 lub1 = -2.554778698e-24 wub1 = -5.575939884e-24 pub1 = 1.422812580e-30
+ uc1 = -2.347726057e-10 luc1 = 5.243018976e-17 wuc1 = 1.144316601e-16 puc1 = -2.919952671e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.153 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 6.3e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.143603+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43165561
+ k2 = 0.046387026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
+ voff = {-0.16725342+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.5720692+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.00827017
+ ua = -7.4124916e-10
+ ub = 6.3364395e-19
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = 5.7286e-9
+ b1 = 3.5674e-8
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.154 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 6.3e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.136052763e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.514439310e-07 wvth0 = -7.105427358e-21
+ k1 = 4.169789897e-01 lk1 = 2.943861458e-7
+ k2 = 6.562039979e-02 lk2 = -3.857862811e-7
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.172472591e-06 lcit = 1.303205335e-10 wcit = 1.355252716e-26 pcit = -1.626303259e-31
+ voff = {-1.346023867e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.549199771e-7
+ nfactor = {1.621526756e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -9.920280577e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 6.971914874e-03 lu0 = 2.604062203e-8
+ ua = -7.228111739e-10 lua = -3.698322591e-16
+ ub = 2.485336107e-19 lub = 7.724608655e-24
+ uc = -1.046491178e-10 luc = -2.033642163e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.297654578e+04 lvsat = -2.571566868e-01 wvsat = -4.656612873e-16
+ a0 = 1.627231194e+00 la0 = -3.274119030e-6
+ ags = 1.127413528e-01 lags = 1.100485920e-8
+ a1 = 0.0
+ a2 = 1.084157408e+00 la2 = -2.289788703e-6
+ b0 = 1.075896438e-07 lb0 = -2.043146133e-12 wb0 = -1.588186776e-28 pb0 = -5.082197684e-33
+ b1 = 5.694535280e-08 lb1 = -4.266644107e-13
+ keta = 3.426055353e-02 lketa = -2.186199026e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.958323949e-02 lpclm = 1.696584997e-06 wpclm = 2.220446049e-22 ppclm = -1.776356839e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 1.912368050e-03 lpdiblc2 = -1.274113513e-8
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 8.855588799e-09 lpscbe2 = 2.417082098e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.715141667e-11 lalpha0 = 1.346934531e-15
+ alpha1 = -6.715141667e-11 lalpha1 = 1.346934531e-15
+ beta0 = 4.813088250e+01 lbeta0 = -3.636723234e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.815887098e-09 lagidl = -1.836585614e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.444180322e-01 lkt1 = 1.237194387e-7
+ kt2 = -6.525229044e-02 lkt2 = 1.345159137e-7
+ at = 7.718690531e+04 lat = -1.242985802e-01 wat = -4.656612873e-16
+ ute = 5.651519091e-01 lute = -1.300034001e-05 wute = 8.881784197e-22 pute = 2.131628207e-26
+ ua1 = 3.782821288e-09 lua1 = -3.395088554e-14 pua1 = -1.058791184e-34
+ ub1 = -2.655052084e-18 lub1 = 2.860600094e-23
+ uc1 = -9.472964564e-11 luc1 = 1.302590510e-15 wuc1 = -2.067951531e-31 puc1 = -3.308722450e-36
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.155 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 6.3e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.150668308e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.366938589e-8
+ k1 = 4.604697380e-01 lk1 = -5.606969765e-8
+ k2 = 1.430285893e-02 lk2 = 2.773918708e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.322146530e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.316562590e-7
+ nfactor = {8.355552889e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.341463636e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 9.316969502e-03 lu0 = 7.143773174e-9
+ ua = -9.431379082e-10 lua = 1.405598021e-15
+ ub = 1.281825696e-18 lub = -6.018346318e-25
+ uc = -1.070056741e-10 luc = -1.346889891e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.346148460e+04 lvsat = -1.931930625e-2
+ a0 = 1.168757490e+00 la0 = 4.203400132e-7
+ ags = 4.417072978e-02 lags = 5.635585964e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = -1.140830746e-07 lb0 = -2.568696835e-13
+ b1 = 9.055190034e-09 lb1 = -4.075733774e-14
+ keta = 7.543931899e-03 lketa = -3.332823646e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -4.156864620e-01 lpclm = 4.485543601e-06 ppclm = 1.421085472e-26
+ pdiblc1 = 0.39
+ pdiblc2 = 2.310096564e-04 lpdiblc2 = 8.075366429e-10
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.465883797e-08 lpscbe2 = -2.259274738e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.014542500e-10 lalpha0 = -8.175355937e-16
+ alpha1 = 2.014542500e-10 lalpha1 = -8.175355937e-16
+ beta0 = -2.439264750e+01 lbeta0 = 2.207346103e-04 pbeta0 = 1.136868377e-25
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.959945019e-10 lagidl = -1.283401221e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.136586484e-01 lkt1 = -1.241449055e-7
+ kt2 = -3.842712868e-02 lkt2 = -8.164580001e-8
+ at = 2.196300907e+04 lat = 3.207049638e-1
+ ute = -1.925921477e+00 lute = 7.073152815e-6
+ ua1 = -2.987663864e-09 lua1 = 2.060683480e-14 wua1 = 3.308722450e-30 pua1 = 3.970466940e-35
+ ub1 = 2.948102001e-18 lub1 = -1.654516721e-23 wub1 = 6.162975822e-39 pub1 = -4.930380658e-44
+ uc1 = 5.590315313e-10 luc1 = -3.965528193e-15 wuc1 = 8.271806126e-31 puc1 = -6.617444900e-36
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.156 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 6.3e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.155676044e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.334714119e-8
+ k1 = 3.842913476e-01 lk1 = 2.530751608e-7
+ k2 = 4.432685200e-02 lk2 = -9.410328086e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.687254897e-01 ldsub = -1.252860521e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.037637994e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.619785835e-8
+ nfactor = {2.243457684e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.720436259e-7
+ eta0 = 1.618122575e-01 leta0 = -3.320080490e-7
+ etab = -1.415214075e-01 letab = 2.902460303e-7
+ u0 = 1.216753903e-02 lu0 = -4.424322556e-9
+ ua = -2.772390642e-10 lua = -1.296732691e-15
+ ub = 8.233204951e-19 lub = 1.258857421e-24
+ uc = -1.342621486e-10 luc = 1.092645171e-16 wuc = -8.271806126e-31
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.432087493e+04 lvsat = -1.039702583e-01 wvsat = 4.656612873e-16
+ a0 = 1.402964339e+00 la0 = -5.301111964e-7
+ ags = -4.821423619e-02 lags = 9.384724937e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = -2.208073870e-07 lb0 = 1.762357191e-13
+ b1 = -1.625453795e-09 lb1 = 2.586530631e-15
+ keta = 2.308642681e-02 lketa = -6.640691024e-08 pketa = 1.110223025e-28
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.045581146e-01 lpclm = 3.452176679e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 4.183469811e-04 lpdiblc2 = 4.728993188e-11
+ pdiblcb = -4.308170000e-01 lpdiblcb = 8.352403749e-7
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 8.705986359e-09 lpscbe2 = 1.564936435e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.029085000e-10 lalpha0 = 4.176201874e-16
+ alpha1 = -1.029085000e-10 lalpha1 = 4.176201874e-16
+ beta0 = 5.514271247e+01 lbeta0 = -1.020334014e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -8.125329299e-11 lagidl = 1.870802463e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.353792873e-01 lkt1 = -3.599886016e-8
+ kt2 = -6.329111093e-02 lkt2 = 1.925646684e-8
+ at = 1.637106726e+05 lat = -2.545311518e-1
+ ute = -8.998158855e-02 lute = -3.774033634e-7
+ ua1 = 2.900604437e-09 lua1 = -3.288758976e-15
+ ub1 = -1.918105286e-18 lub1 = 3.202729218e-24
+ uc1 = -8.850008756e-10 luc1 = 1.894600800e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.157 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 6.3e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.166873031e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.698160864e-9
+ k1 = 5.064385921e-01 lk1 = 1.675366545e-9
+ k2 = -1.550530049e-03 lk2 = 3.201705484e-10
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.600000206e-01 ldsub = -2.177893421e-14
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.008592856e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.021987531e-8
+ nfactor = {2.582745438e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.070355502e-6
+ eta0 = -5.174742150e-01 leta0 = 1.066078990e-06 weta0 = 7.077671782e-22 peta0 = -5.342948306e-28
+ etab = 2.904247369e-04 letab = -1.626828481e-9
+ u0 = 1.299481844e-02 lu0 = -6.127004236e-9
+ ua = -2.335251343e-10 lua = -1.386703390e-15
+ ub = 1.100219537e-18 lub = 6.889521208e-25
+ uc = -1.209494201e-10 luc = 8.186465865e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.474998785e+04 lvsat = 3.921845435e-2
+ a0 = 1.027063579e+00 la0 = 2.435564714e-7
+ ags = 2.421456228e-01 lags = 3.408625427e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = -3.571202000e-08 lb0 = -2.047220124e-13
+ b1 = -8.958356404e-10 lb1 = 1.084852434e-15
+ keta = -1.779393475e-02 lketa = 1.773182353e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.249152049e-01 lpclm = -3.141316846e-7
+ pdiblc1 = 3.959901522e-01 lpdiblc1 = -1.232875161e-8
+ pdiblc2 = 4.533060379e-04 lpdiblc2 = -2.466175011e-11
+ pdiblcb = 1.866340000e-01 lpdiblcb = -4.355787498e-07 wpdiblcb = 2.220446049e-22
+ drout = 3.733753506e-01 ldrout = 3.841052546e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 9.779790288e-09 lpscbe2 = -6.451345974e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.611938067e+00 lbeta0 = 1.967522498e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 3.976755324e-10 lagidl = 8.850855221e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.251515120e-01 lkt1 = -5.704936050e-8
+ kt2 = -5.962353039e-02 lkt2 = 1.170796260e-8
+ at = 2.764051955e+04 lat = 2.552435502e-2
+ ute = 5.465304861e-01 lute = -1.687453420e-06 pute = 3.552713679e-27
+ ua1 = 3.136618649e-09 lua1 = -3.774516346e-15
+ ub1 = -1.649671782e-18 lub1 = 2.650247432e-24 wub1 = -3.081487911e-39 pub1 = 3.081487911e-45
+ uc1 = 2.307099871e-12 luc1 = 6.837014368e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.158 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 6.3e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.186764098e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.074629071e-8
+ k1 = 5.895983608e-01 lk1 = -8.632180590e-8
+ k2 = -4.236429828e-02 lk2 = 4.350807568e-08 wk2 = 5.551115123e-23 pk2 = -6.245004514e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -5.660916000e-01 ldsub = 8.741453484e-07 pdsub = 1.776356839e-27
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.251342609e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.590692590e-8
+ nfactor = {3.163637012e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.685037539e-6
+ eta0 = 1.027885506e+00 leta0 = -5.691743056e-7
+ etab = -1.522680668e-03 letab = 2.917452658e-10
+ u0 = 7.157921276e-03 lu0 = 4.942524115e-11
+ ua = -2.676735973e-09 lua = 1.198629023e-15
+ ub = 3.551846133e-18 lub = -1.905285595e-24
+ uc = -3.828526639e-11 luc = -5.608068851e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -7.419646049e+02 lvsat = 5.561157368e-2
+ a0 = 1.416791016e+00 la0 = -1.688414103e-7
+ ags = -2.012374473e-01 lags = 8.100372059e-7
+ a1 = 0.0
+ a2 = 1.143658537e+00 la2 = -3.636491546e-7
+ b0 = -3.936436742e-07 lb0 = 1.740305261e-13
+ b1 = 3.566568533e-09 lb1 = -3.637129790e-15 wb1 = -4.963083675e-30 pb1 = -3.308722450e-36
+ keta = 4.640102772e-02 lketa = -5.019735991e-08 wketa = 4.163336342e-23 pketa = -5.551115123e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 8.463474809e-01 lpclm = -2.309936761e-7
+ pdiblc1 = 7.353910455e-01 lpdiblc1 = -3.714725948e-7
+ pdiblc2 = 1.290151741e-05 lpdiblc2 = 4.413611013e-10
+ pdiblcb = -0.225
+ drout = 9.868614715e-01 ldrout = -2.650673539e-7
+ pscbe1 = 1.538699225e+09 lpscbe1 = -7.816693584e+02 ppscbe1 = -3.814697266e-18
+ pscbe2 = -6.786262656e-08 lpscbe2 = 8.151374164e-14 wpscbe2 = -1.058791184e-28 ppscbe2 = -5.293955920e-35
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.271197094e+00 lbeta0 = 2.328084373e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.592126185e-09 lagidl = -3.788463250e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.736892727e-01 lkt1 = -5.688158284e-9
+ kt2 = -3.629638816e-02 lkt2 = -1.297611950e-8
+ at = 2.023824718e+04 lat = 3.335721757e-2
+ ute = -1.951903787e+00 lute = 9.563147749e-7
+ ua1 = -2.770257084e-09 lua1 = 2.475962349e-15 wua1 = 3.308722450e-30 pua1 = -6.617444900e-36
+ ub1 = 2.776470114e-18 lub1 = -2.033363139e-24 pub1 = -6.162975822e-45
+ uc1 = 2.168072778e-10 luc1 = -1.586075096e-16 puc1 = 4.135903063e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.159 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 6.3e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.198442244e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.726468175e-8
+ k1 = 2.587759691e-01 lk1 = 9.833332850e-8
+ k2 = 1.264619903e-01 lk2 = -5.072569381e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.265530550e+00 ldsub = -1.482111871e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.432797432e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -9.781810251e-9
+ nfactor = {-1.369102099e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.450014502e-07 pnfactor = 1.776356839e-27
+ eta0 = -5.857710121e-01 leta0 = 3.315203530e-07 weta0 = -1.221245327e-21 peta0 = 8.049116929e-28
+ etab = -2.144165608e-03 letab = 6.386395146e-10
+ u0 = 9.588264965e-03 lu0 = -1.307119696e-09 wu0 = 5.551115123e-23
+ ua = -4.524496467e-10 lua = -4.290087548e-17
+ ub = 1.800632172e-19 lub = -2.325752460e-26
+ uc = -1.066909176e-10 luc = 3.257391349e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.745291629e+03 lvsat = 5.087424187e-2
+ a0 = 1.730312949e+00 la0 = -3.438399480e-7
+ ags = 9.336688757e-01 lags = 1.765665437e-7
+ a1 = 0.0
+ a2 = 1.175865985e-01 la2 = 2.090734196e-7
+ b0 = -1.827582555e-07 lb0 = 5.632061198e-14
+ b1 = -6.585512924e-09 lb1 = 2.029457517e-15
+ keta = -5.806135818e-02 lketa = 8.110410026e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.801832138e-01 lpclm = 1.408392328e-7
+ pdiblc1 = -3.427765615e-01 lpdiblc1 = 2.303282184e-07 ppdiblc1 = 2.220446049e-28
+ pdiblc2 = -8.777845214e-03 lpdiblc2 = 5.348092205e-09 wpdiblc2 = 2.775557562e-23 ppdiblc2 = 3.469446952e-30
+ pdiblcb = -1.473166890e-01 lpdiblcb = -4.336049373e-8
+ drout = 4.913817236e-01 ldrout = 1.149457697e-8
+ pscbe1 = -6.773655310e+08 lpscbe1 = 4.552715062e+02 wpscbe1 = -1.907348633e-12 ppscbe1 = 4.768371582e-19
+ pscbe2 = 1.636367297e-07 lpscbe2 = -4.770225404e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.865441218e+00 lbeta0 = 3.218851306e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.041584712e-09 lagidl = -6.297205910e-16
+ bgidl = 7.033052157e+08 lbgidl = 1.656061277e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.00081386752815302
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207367379934e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.360991252e-01 lkt1 = -2.666985086e-8
+ kt2 = -6.784093954e-02 lkt2 = 4.631102743e-9
+ at = 9.493059464e+04 lat = -8.333810011e-3
+ ute = 4.960630988e-01 lute = -4.100669019e-07 pute = 8.881784197e-28
+ ua1 = 3.355066581e-09 lua1 = -9.430095617e-16
+ ub1 = -1.725764093e-18 lub1 = 4.796489289e-25
+ uc1 = -2.970663052e-11 luc1 = -2.101084137e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.160 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.3e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.239991813e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.006901243e-8
+ k1 = -1.102372845e+00 lk1 = 5.177985587e-7
+ k2 = 4.847969085e-01 lk2 = -1.611537656e-07 pk2 = 2.220446049e-28
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.977511515e+00 ldsub = -3.676223612e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-3.638620714e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.819504583e-8
+ nfactor = {2.927995871e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.792352313e-7
+ eta0 = 4.900000008e-01 leta0 = -9.356071473e-17
+ etab = 2.581819860e-03 letab = -8.177674270e-10 wetab = -1.734723476e-24
+ u0 = 1.290521855e-02 lu0 = -2.329305283e-9
+ ua = 2.912788267e-09 lua = -1.079966243e-15
+ ub = -2.678685290e-18 lub = 8.577230029e-25 wub = 6.162975822e-39 pub = -1.540743956e-45
+ uc = 4.100502134e-11 luc = -1.294154402e-17 wuc = 2.584939414e-32 puc = 2.584939414e-38
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.107233529e+05 lvsat = -1.041285073e-1
+ a0 = -2.787929715e-01 la0 = 2.753062236e-7
+ ags = 2.379753986e+00 lags = -2.690735049e-7
+ a1 = 0.0
+ a2 = 9.570523633e-01 la2 = -4.962474518e-8
+ b0 = -4.369331260e-14 lb0 = 1.383167812e-20 wb0 = -7.573064690e-35 pb0 = -6.310887242e-42
+ b1 = -1.379167911e-17 lb1 = 3.284876207e-24
+ keta = -9.702710173e-02 lketa = 2.011848322e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.931004364e-01 lpclm = -1.722646764e-8
+ pdiblc1 = 5.732445572e-01 lpdiblc1 = -5.196200978e-8
+ pdiblc2 = 3.354825457e-02 lpdiblc2 = -7.695541966e-9
+ pdiblcb = 2.607591983e+00 lpdiblcb = -8.923406993e-7
+ drout = -1.074947477e+00 ldrout = 4.941902469e-7
+ pscbe1 = 7.998824354e+08 lpscbe1 = 2.800036250e-2
+ pscbe2 = 2.140020980e-08 lpscbe2 = -3.869225705e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.080169809e+01 lbeta0 = -5.829811493e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -3.530736764e-09 lagidl = 1.087501718e-15 wagidl = -1.861156378e-30 pagidl = -2.352294867e-36
+ bgidl = 2.059624081e+09 lbgidl = -2.523706570e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.00081386752815302
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207367379934e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.047221533e-01 lkt1 = -6.715629230e-8
+ kt2 = -5.971042874e-02 lkt2 = 2.125523229e-9
+ at = 2.366743202e+05 lat = -5.201497393e-2
+ ute = -2.029992490e+00 lute = 3.683876490e-7
+ ua1 = 1.080932106e-10 lua1 = 5.761022195e-17
+ ub1 = -3.579906755e-19 lub1 = 5.814219486e-26
+ uc1 = -3.312416379e-10 luc1 = 7.191320187e-17 puc1 = -4.135903063e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.161 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.3e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -3.7585e-8
+ vth0 = {-2.810850035e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.909680141e-06 wvth0 = 1.508074191e-05 pvth0 = -3.848152914e-12
+ k1 = 2.203721088e-01 lk1 = 2.172329406e-07 wk1 = 4.741221247e-07 pk1 = -1.209817426e-13
+ k2 = -1.856359089e+01 lk2 = 4.687920581e-06 wk2 = 1.023163425e-05 pk2 = -2.610806112e-12
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -5.476699010e+00 ldsub = 1.508228541e-06 wdsub = 3.291788298e-06 pdsub = -8.399656200e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-7.218421820e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.838874914e-05 wvoff = 4.013441606e-05 pvoff = -1.024109895e-11
+ nfactor = {5.412193772e+02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.378692537e-04 wnfactor = -3.009069266e-04 pnfactor = 7.678242046e-11
+ eta0 = -1.159313922e+01 leta0 = 3.083254636e-06 weta0 = 6.729366065e-06 peta0 = -1.717132339e-12
+ etab = -6.869665587e-01 letab = 1.750759221e-07 wetab = 3.821124031e-07 petab = -9.750362190e-14
+ u0 = -1.872561060e-01 lu0 = 4.857959972e-08 wu0 = 1.060275304e-07 pu0 = -2.705504494e-14
+ ua = -3.031727040e-07 lua = 7.694678343e-14 wua = 1.679404180e-13 pua = -4.285335647e-20
+ ub = 4.613163166e-16 lub = -1.174786594e-22 wub = -2.564033780e-22 pub = 6.542644996e-29
+ uc = 5.159472478e-10 luc = -1.350562881e-16 wuc = -2.947674749e-16 puc = 7.521581658e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.564931368e+07 lvsat = -1.928467504e+01 wvsat = -4.208982165e+01 pvsat = 1.074005979e-5
+ a0 = 6.271206215e+00 la0 = -1.376406375e-06 wa0 = -3.004078729e-06 pa0 = 7.665507692e-13
+ ags = 1.250000077e+00 lags = -1.754415280e-14 wags = -2.471324478e-15 pags = 6.306066780e-22
+ a1 = 0.0
+ a2 = 8.995225520e+00 la2 = -2.104267484e-06 wa2 = -4.592674872e-06 pa2 = 1.171912847e-12
+ b0 = -3.741268902e-05 lb0 = 9.546595861e-12 wb0 = 2.083594966e-11 pb0 = -5.316709275e-18
+ b1 = 3.999568671e-21 lb1 = -9.005828797e-28 wb1 = -3.808420539e-35 pb1 = 9.717947591e-42
+ keta = 2.111861687e+00 lketa = -5.420876601e-07 wketa = -1.183134929e-06 pketa = 3.019005397e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.657719152e-01 lpclm = -1.148263258e-08 wpclm = -2.506143767e-08 ppclm = 6.394927049e-15
+ pdiblc1 = -6.902533407e+00 lpdiblc1 = 1.851923331e-06 wpdiblc1 = 4.041920725e-06 ppdiblc1 = -1.031376911e-12
+ pdiblc2 = 3.614446410e-02 lpdiblc2 = -8.907305972e-09 wpdiblc2 = -1.944067023e-08 ppdiblc2 = 4.960675822e-15
+ pdiblcb = 4.104240453e+01 lpdiblcb = -1.076344494e-05 wpdiblcb = -2.349178700e-05 ppdiblcb = 5.994399290e-12
+ drout = 1.000000075e+00 ldrout = -1.245808789e-14 wdrout = 8.105763527e-14 pdrout = -2.068347982e-20
+ pscbe1 = 3.716511143e+07 lpscbe1 = 1.946525785e+02 wpscbe1 = 4.248395321e+02 ppscbe1 = -1.084063034e-4
+ pscbe2 = 1.648999131e-07 lpscbe2 = -4.076222098e-14 wpscbe2 = -8.896570247e-14 ppscbe2 = 2.270137830e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -5.978599455e+00 lbeta0 = 3.657235587e-06 wbeta0 = 7.982109199e-06 pbeta0 = -2.036794804e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -4.239719767e-07 lagidl = 1.084491162e-13 wagidl = 2.366959218e-13 pagidl = -6.039769836e-20
+ bgidl = 1.000000484e+09 lbgidl = -1.123832397e-04 wbgidl = -6.289721680e-05 pbgidl = 1.604947662e-11
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -2.8385e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.346826027e-02 lkt1 = -1.462690023e-07 wkt1 = -3.192400017e-07 pkt1 = 8.146047123e-14
+ kt2 = -1.730770971e+00 lkt2 = 4.286817564e-07 wkt2 = 9.356204315e-07 pkt2 = -2.387422655e-13
+ at = 1.503860742e+06 lat = -3.790756365e-01 wat = -8.273525717e-01 pat = 2.111155557e-7
+ ute = 1.220414244e+01 lute = -3.237441940e-06 wute = -7.065888171e-06 pute = 1.803002684e-12
+ ua1 = 1.595303410e-08 lua1 = -3.981431265e-15 wua1 = -8.689683193e-15 pua1 = 2.217346460e-21
+ ub1 = -2.126402367e-17 lub1 = 5.396884685e-24 wub1 = 1.177898536e-23 pub1 = -3.005643694e-30
+ uc1 = -5.086906146e-10 luc1 = 1.223258481e-16 wuc1 = 2.669826255e-16 puc1 = -6.812595654e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.162 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.5e-07 wmax = 6.3e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.143603+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43165561
+ k2 = 0.046387026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
+ voff = {-0.16725342+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.5720692+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.00827017
+ ua = -7.4124916e-10
+ ub = 6.3364395e-19
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = 5.7286e-9
+ b1 = 3.5674e-8
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.163 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.5e-07 wmax = 6.3e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.136052763e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.514439310e-7
+ k1 = 4.169789897e-01 lk1 = 2.943861458e-7
+ k2 = 6.562039979e-02 lk2 = -3.857862811e-07 wk2 = 2.775557562e-23
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.172472591e-06 lcit = 1.303205335e-10 wcit = 1.694065895e-27 pcit = 8.470329473e-33
+ voff = {-1.346023867e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.549199771e-7
+ nfactor = {1.621526756e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -9.920280577e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 6.971914874e-03 lu0 = 2.604062203e-8
+ ua = -7.228111739e-10 lua = -3.698322591e-16
+ ub = 2.485336107e-19 lub = 7.724608655e-24
+ uc = -1.046491178e-10 luc = -2.033642163e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.297654578e+04 lvsat = -2.571566868e-01 wvsat = -5.820766091e-17
+ a0 = 1.627231194e+00 la0 = -3.274119030e-06 wa0 = -8.881784197e-22
+ ags = 1.127413528e-01 lags = 1.100485920e-8
+ a1 = 0.0
+ a2 = 1.084157408e+00 la2 = -2.289788703e-6
+ b0 = 1.075896438e-07 lb0 = -2.043146133e-12 wb0 = -1.985233470e-29 pb0 = -1.588186776e-34
+ b1 = 5.694535280e-08 lb1 = -4.266644107e-13
+ keta = 3.426055353e-02 lketa = -2.186199026e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.958323949e-02 lpclm = 1.696584997e-06 ppclm = 1.110223025e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 1.912368050e-03 lpdiblc2 = -1.274113513e-8
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 8.855588799e-09 lpscbe2 = 2.417082098e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.715141667e-11 lalpha0 = 1.346934531e-15
+ alpha1 = -6.715141667e-11 lalpha1 = 1.346934531e-15
+ beta0 = 4.813088250e+01 lbeta0 = -3.636723234e-04 pbeta0 = -2.273736754e-25
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.815887098e-09 lagidl = -1.836585614e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.444180322e-01 lkt1 = 1.237194387e-7
+ kt2 = -6.525229044e-02 lkt2 = 1.345159137e-7
+ at = 7.718690531e+04 lat = -1.242985802e-1
+ ute = 5.651519091e-01 lute = -1.300034001e-05 pute = -8.881784197e-28
+ ua1 = 3.782821288e-09 lua1 = -3.395088554e-14
+ ub1 = -2.655052084e-18 lub1 = 2.860600094e-23
+ uc1 = -9.472964564e-11 luc1 = 1.302590510e-15 puc1 = 2.067951531e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.164 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.5e-07 wmax = 6.3e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.150668308e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.366938589e-8
+ k1 = 4.604697380e-01 lk1 = -5.606969765e-8
+ k2 = 1.430285893e-02 lk2 = 2.773918708e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.322146530e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.316562590e-7
+ nfactor = {8.355552889e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.341463636e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 9.316969502e-03 lu0 = 7.143773174e-9
+ ua = -9.431379082e-10 lua = 1.405598021e-15
+ ub = 1.281825696e-18 lub = -6.018346318e-25
+ uc = -1.070056741e-10 luc = -1.346889891e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.346148460e+04 lvsat = -1.931930625e-2
+ a0 = 1.168757490e+00 la0 = 4.203400132e-7
+ ags = 4.417072978e-02 lags = 5.635585964e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = -1.140830747e-07 lb0 = -2.568696835e-13
+ b1 = 9.055190034e-09 lb1 = -4.075733774e-14
+ keta = 7.543931899e-03 lketa = -3.332823646e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -4.156864620e-01 lpclm = 4.485543601e-06 wpclm = -1.110223025e-22 ppclm = -4.440892099e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 2.310096564e-04 lpdiblc2 = 8.075366429e-10
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.465883797e-08 lpscbe2 = -2.259274738e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.014542500e-10 lalpha0 = -8.175355937e-16
+ alpha1 = 2.014542500e-10 lalpha1 = -8.175355937e-16
+ beta0 = -2.439264750e+01 lbeta0 = 2.207346103e-04 pbeta0 = 4.263256415e-26
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.959945019e-10 lagidl = -1.283401221e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.136586484e-01 lkt1 = -1.241449055e-7
+ kt2 = -3.842712868e-02 lkt2 = -8.164580001e-8
+ at = 2.196300907e+04 lat = 3.207049638e-1
+ ute = -1.925921477e+00 lute = 7.073152815e-06 pute = 3.552713679e-27
+ ua1 = -2.987663864e-09 lua1 = 2.060683480e-14 wua1 = -4.135903063e-31 pua1 = 3.308722450e-36
+ ub1 = 2.948102001e-18 lub1 = -1.654516721e-23
+ uc1 = 5.590315313e-10 luc1 = -3.965528193e-15 wuc1 = 1.033975766e-31 puc1 = -6.203854594e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.165 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.5e-07 wmax = 6.3e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.155676044e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.334714119e-8
+ k1 = 3.842913476e-01 lk1 = 2.530751608e-7
+ k2 = 4.432685200e-02 lk2 = -9.410328086e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.687254897e-01 ldsub = -1.252860521e-06 wdsub = 4.440892099e-22
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.037637994e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.619785835e-8
+ nfactor = {2.243457684e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.720436259e-7
+ eta0 = 1.618122575e-01 leta0 = -3.320080490e-7
+ etab = -1.415214075e-01 letab = 2.902460303e-7
+ u0 = 1.216753903e-02 lu0 = -4.424322556e-9
+ ua = -2.772390642e-10 lua = -1.296732691e-15
+ ub = 8.233204951e-19 lub = 1.258857421e-24
+ uc = -1.342621486e-10 luc = 1.092645171e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.432087493e+04 lvsat = -1.039702583e-1
+ a0 = 1.402964339e+00 la0 = -5.301111964e-7
+ ags = -4.821423619e-02 lags = 9.384724937e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = -2.208073870e-07 lb0 = 1.762357191e-13
+ b1 = -1.625453795e-09 lb1 = 2.586530631e-15 wb1 = 8.271806126e-31
+ keta = 2.308642681e-02 lketa = -6.640691024e-08 wketa = 6.938893904e-24 pketa = 1.387778781e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.045581146e-01 lpclm = 3.452176679e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 4.183469811e-04 lpdiblc2 = 4.728993188e-11
+ pdiblcb = -4.308170000e-01 lpdiblcb = 8.352403749e-7
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 8.705986359e-09 lpscbe2 = 1.564936435e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.029085000e-10 lalpha0 = 4.176201874e-16
+ alpha1 = -1.029085000e-10 lalpha1 = 4.176201874e-16
+ beta0 = 5.514271247e+01 lbeta0 = -1.020334014e-04 pbeta0 = -5.684341886e-26
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -8.125329299e-11 lagidl = 1.870802463e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.353792873e-01 lkt1 = -3.599886016e-8
+ kt2 = -6.329111093e-02 lkt2 = 1.925646684e-8
+ at = 1.637106726e+05 lat = -2.545311518e-1
+ ute = -8.998158855e-02 lute = -3.774033634e-7
+ ua1 = 2.900604438e-09 lua1 = -3.288758976e-15
+ ub1 = -1.918105286e-18 lub1 = 3.202729218e-24
+ uc1 = -8.850008756e-10 luc1 = 1.894600800e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.166 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.5e-07 wmax = 6.3e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.166873031e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.698160864e-9
+ k1 = 5.064385921e-01 lk1 = 1.675366545e-9
+ k2 = -1.550530049e-03 lk2 = 3.201705484e-10
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.600000206e-01 ldsub = -2.177893732e-14
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.008592856e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.021987531e-8
+ nfactor = {2.582745438e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.070355502e-06 wnfactor = 1.776356839e-21
+ eta0 = -5.174742150e-01 leta0 = 1.066078990e-06 weta0 = -5.507747036e-23 peta0 = -2.077331362e-28
+ etab = 2.904247369e-04 letab = -1.626828481e-09 petab = -4.336808690e-31
+ u0 = 1.299481844e-02 lu0 = -6.127004236e-9
+ ua = -2.335251343e-10 lua = -1.386703390e-15
+ ub = 1.100219537e-18 lub = 6.889521208e-25
+ uc = -1.209494201e-10 luc = 8.186465865e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.474998785e+04 lvsat = 3.921845435e-2
+ a0 = 1.027063579e+00 la0 = 2.435564714e-7
+ ags = 2.421456228e-01 lags = 3.408625427e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = -3.571202000e-08 lb0 = -2.047220124e-13
+ b1 = -8.958356404e-10 lb1 = 1.084852434e-15 wb1 = 4.135903063e-31
+ keta = -1.779393475e-02 lketa = 1.773182353e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.249152049e-01 lpclm = -3.141316846e-7
+ pdiblc1 = 3.959901522e-01 lpdiblc1 = -1.232875161e-8
+ pdiblc2 = 4.533060379e-04 lpdiblc2 = -2.466175011e-11
+ pdiblcb = 1.866340000e-01 lpdiblcb = -4.355787498e-07 ppdiblcb = -5.551115123e-29
+ drout = 3.733753506e-01 ldrout = 3.841052546e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 9.779790288e-09 lpscbe2 = -6.451345974e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.611938067e+00 lbeta0 = 1.967522498e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 3.976755324e-10 lagidl = 8.850855221e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.251515120e-01 lkt1 = -5.704936050e-8
+ kt2 = -5.962353039e-02 lkt2 = 1.170796260e-8
+ at = 2.764051955e+04 lat = 2.552435502e-2
+ ute = 5.465304861e-01 lute = -1.687453420e-06 pute = -2.220446049e-28
+ ua1 = 3.136618649e-09 lua1 = -3.774516346e-15
+ ub1 = -1.649671782e-18 lub1 = 2.650247432e-24 pub1 = 3.851859889e-46
+ uc1 = 2.307099871e-12 luc1 = 6.837014368e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.167 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.5e-07 wmax = 6.3e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.186764098e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.074629071e-8
+ k1 = 5.895983608e-01 lk1 = -8.632180590e-8
+ k2 = -4.236429828e-02 lk2 = 4.350807568e-08 wk2 = 1.734723476e-24 pk2 = 8.673617380e-31
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -5.660916000e-01 ldsub = 8.741453484e-07 pdsub = -2.220446049e-28
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.251342609e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.590692590e-8
+ nfactor = {3.163637012e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.685037539e-6
+ eta0 = 1.027885506e+00 leta0 = -5.691743056e-7
+ etab = -1.522680668e-03 letab = 2.917452658e-10
+ u0 = 7.157921276e-03 lu0 = 4.942524115e-11
+ ua = -2.676735973e-09 lua = 1.198629023e-15 pua = 8.271806126e-37
+ ub = 3.551846133e-18 lub = -1.905285595e-24
+ uc = -3.828526639e-11 luc = -5.608068851e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -7.419646049e+02 lvsat = 5.561157368e-2
+ a0 = 1.416791016e+00 la0 = -1.688414103e-7
+ ags = -2.012374473e-01 lags = 8.100372059e-7
+ a1 = 0.0
+ a2 = 1.143658537e+00 la2 = -3.636491546e-7
+ b0 = -3.936436742e-07 lb0 = 1.740305261e-13 pb0 = -1.058791184e-34
+ b1 = 3.566568533e-09 lb1 = -3.637129790e-15 wb1 = 3.101927297e-31 pb1 = 6.203854594e-37
+ keta = 4.640102772e-02 lketa = -5.019735991e-08 wketa = 8.673617380e-25 pketa = -1.214306433e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 8.463474809e-01 lpclm = -2.309936761e-7
+ pdiblc1 = 7.353910455e-01 lpdiblc1 = -3.714725948e-07 ppdiblc1 = 2.220446049e-28
+ pdiblc2 = 1.290151741e-05 lpdiblc2 = 4.413611013e-10
+ pdiblcb = -0.225
+ drout = 9.868614715e-01 ldrout = -2.650673539e-7
+ pscbe1 = 1.538699225e+09 lpscbe1 = -7.816693584e+2
+ pscbe2 = -6.786262656e-08 lpscbe2 = 8.151374164e-14 wpscbe2 = -1.323488980e-29 ppscbe2 = -1.323488980e-35
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.271197094e+00 lbeta0 = 2.328084373e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.592126185e-09 lagidl = -3.788463250e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.736892727e-01 lkt1 = -5.688158284e-9
+ kt2 = -3.629638816e-02 lkt2 = -1.297611950e-8
+ at = 2.023824718e+04 lat = 3.335721757e-2
+ ute = -1.951903787e+00 lute = 9.563147749e-7
+ ua1 = -2.770257084e-09 lua1 = 2.475962349e-15 wua1 = 4.135903063e-31 pua1 = 4.135903063e-37
+ ub1 = 2.776470114e-18 lub1 = -2.033363139e-24 wub1 = -7.703719778e-40 pub1 = -3.851859889e-46
+ uc1 = 2.168072778e-10 luc1 = -1.586075096e-16 wuc1 = 5.169878828e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.168 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.5e-07 wmax = 6.3e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.198442244e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.726468175e-8
+ k1 = 2.587759691e-01 lk1 = 9.833332850e-8
+ k2 = 1.264619903e-01 lk2 = -5.072569381e-08 pk2 = 1.387778781e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.265530550e+00 ldsub = -1.482111871e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.432797432e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -9.781810251e-9
+ nfactor = {-1.369102099e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.450014502e-07 wnfactor = 2.220446049e-22
+ eta0 = -5.857710121e-01 leta0 = 3.315203530e-07 weta0 = -1.040834086e-22 peta0 = 1.040834086e-29
+ etab = -2.144165608e-03 letab = 6.386395146e-10
+ u0 = 9.588264965e-03 lu0 = -1.307119696e-9
+ ua = -4.524496467e-10 lua = -4.290087548e-17
+ ub = 1.800632172e-19 lub = -2.325752460e-26
+ uc = -1.066909176e-10 luc = 3.257391349e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.745291629e+03 lvsat = 5.087424187e-2
+ a0 = 1.730312949e+00 la0 = -3.438399480e-7
+ ags = 9.336688757e-01 lags = 1.765665437e-7
+ a1 = 0.0
+ a2 = 1.175865985e-01 la2 = 2.090734196e-7
+ b0 = -1.827582555e-07 lb0 = 5.632061198e-14
+ b1 = -6.585512924e-09 lb1 = 2.029457517e-15
+ keta = -5.806135818e-02 lketa = 8.110410026e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.801832138e-01 lpclm = 1.408392328e-7
+ pdiblc1 = -3.427765615e-01 lpdiblc1 = 2.303282184e-7
+ pdiblc2 = -8.777845214e-03 lpdiblc2 = 5.348092205e-09 wpdiblc2 = 8.673617380e-25 ppdiblc2 = -1.301042607e-30
+ pdiblcb = -1.473166890e-01 lpdiblcb = -4.336049373e-8
+ drout = 4.913817236e-01 ldrout = 1.149457697e-8
+ pscbe1 = -6.773655310e+08 lpscbe1 = 4.552715062e+02 ppscbe1 = -5.960464478e-20
+ pscbe2 = 1.636367297e-07 lpscbe2 = -4.770225404e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.865441218e+00 lbeta0 = 3.218851306e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.041584712e-09 lagidl = -6.297205910e-16
+ bgidl = 7.033052157e+08 lbgidl = 1.656061277e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.00081386752815302
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207367379934e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.360991252e-01 lkt1 = -2.666985086e-8
+ kt2 = -6.784093954e-02 lkt2 = 4.631102743e-9
+ at = 9.493059464e+04 lat = -8.333810011e-3
+ ute = 4.960630988e-01 lute = -4.100669019e-07 pute = -1.110223025e-28
+ ua1 = 3.355066581e-09 lua1 = -9.430095617e-16 pua1 = 4.135903063e-37
+ ub1 = -1.725764093e-18 lub1 = 4.796489289e-25
+ uc1 = -2.970663052e-11 luc1 = -2.101084137e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.169 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.5e-07 wmax = 6.3e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.239991813e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.006901243e-8
+ k1 = -1.102372845e+00 lk1 = 5.177985587e-7
+ k2 = 4.847969085e-01 lk2 = -1.611537656e-07 pk2 = -2.775557562e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.977511515e+00 ldsub = -3.676223612e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-3.638620714e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.819504583e-8
+ nfactor = {2.927995871e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.792352313e-7
+ eta0 = 4.900000008e-01 leta0 = -9.356115882e-17
+ etab = 2.581819860e-03 letab = -8.177674270e-10 wetab = 4.336808690e-25 petab = -2.710505431e-32
+ u0 = 1.290521855e-02 lu0 = -2.329305283e-9
+ ua = 2.912788267e-09 lua = -1.079966243e-15
+ ub = -2.678685290e-18 lub = 8.577230029e-25 wub = -3.851859889e-40
+ uc = 4.100502134e-11 luc = -1.294154402e-17 wuc = 8.077935669e-33 puc = -4.038967835e-40
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.107233529e+05 lvsat = -1.041285073e-1
+ a0 = -2.787929715e-01 la0 = 2.753062236e-7
+ ags = 2.379753986e+00 lags = -2.690735049e-7
+ a1 = 0.0
+ a2 = 9.570523633e-01 la2 = -4.962474518e-8
+ b0 = -4.369331260e-14 lb0 = 1.383167812e-20 wb0 = -6.310887242e-36 pb0 = 1.577721810e-42
+ b1 = -1.379167911e-17 lb1 = 3.284876207e-24
+ keta = -9.702710173e-02 lketa = 2.011848322e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.931004364e-01 lpclm = -1.722646764e-8
+ pdiblc1 = 5.732445572e-01 lpdiblc1 = -5.196200978e-8
+ pdiblc2 = 3.354825457e-02 lpdiblc2 = -7.695541966e-9
+ pdiblcb = 2.607591983e+00 lpdiblcb = -8.923406993e-07 wpdiblcb = 8.881784197e-22
+ drout = -1.074947477e+00 ldrout = 4.941902469e-7
+ pscbe1 = 7.998824354e+08 lpscbe1 = 2.800036250e-2
+ pscbe2 = 2.140020980e-08 lpscbe2 = -3.869225705e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.080169809e+01 lbeta0 = -5.829811493e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -3.530736764e-09 lagidl = 1.087501718e-15 wagidl = 4.652890946e-31 pagidl = -9.208846663e-38
+ bgidl = 2.059624081e+09 lbgidl = -2.523706570e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.00081386752815302
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207367379934e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.047221533e-01 lkt1 = -6.715629230e-8
+ kt2 = -5.971042874e-02 lkt2 = 2.125523229e-9
+ at = 2.366743202e+05 lat = -5.201497393e-2
+ ute = -2.029992490e+00 lute = 3.683876490e-7
+ ua1 = 1.080932106e-10 lua1 = 5.761022195e-17
+ ub1 = -3.579906755e-19 lub1 = 5.814219486e-26
+ uc1 = -3.312416379e-10 luc1 = 7.191320187e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.170 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.5e-07 wmax = 6.3e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -3.7585e-8
+ vth0 = {4.855709437e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.501797270e-06 wvth0 = -2.948109631e-06 pvth0 = 7.522691344e-13
+ k1 = 2.373406629e-01 lk1 = 2.129030746e-07 wk1 = 4.648416492e-07 pk1 = -1.186136436e-13
+ k2 = 3.149838409e+00 lk2 = -8.526951723e-07 wk2 = -1.643917924e-06 pk2 = 4.194785368e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -5.358887946e+00 ldsub = 1.478166692e-06 wdsub = 3.227354836e-06 pdsub = -8.235241334e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {1.055589365e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -2.724045199e-06 wvoff = -5.117971391e-06 pvoff = 1.305952760e-12
+ nfactor = {-3.289670969e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.627948231e-06 wnfactor = 1.308979184e-05 pnfactor = -3.340122184e-12
+ eta0 = -1.135230044e+01 leta0 = 3.021799803e-06 weta0 = 6.597646034e-06 peta0 = -1.683521339e-12
+ etab = -6.732909212e-01 letab = 1.715863097e-07 wetab = 3.746328961e-07 petab = -9.559507609e-14
+ u0 = -5.486089861e-02 lu0 = 1.479631464e-08 wu0 = 3.361767881e-08 pu0 = -8.578223102e-15
+ ua = -6.078191387e-09 lua = 1.137176650e-15 wua = 5.452893038e-15 pua = -1.391414716e-21
+ ub = -9.442467106e-18 lub = 2.644859408e-24 wub = 1.064957539e-24 pub = -2.717452153e-31
+ uc = 5.053976959e-10 luc = -1.323643590e-16 wuc = -2.889976929e-16 puc = 7.374354129e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -6.691101680e+06 lvsat = 1.726128745e+00 wvsat = 2.943963002e+00 pvsat = -7.512110391e-7
+ a0 = 6.163692469e+00 la0 = -1.348972092e-06 wa0 = -2.945277096e-06 pa0 = 7.515463565e-13
+ ags = 1.250000072e+00 lags = -1.627033441e-14 wags = 2.589999326e-16 pags = -6.608846803e-23
+ a1 = 0.0
+ a2 = 8.830856808e+00 la2 = -2.062325520e-06 wa2 = -4.502778008e-06 pa2 = 1.148973864e-12
+ b0 = 4.676586265e-06 lb0 = -1.193324514e-12 wb0 = -2.183600955e-12 pb0 = 5.571894557e-19
+ b1 = 3.999568594e-21 lb1 = -9.005828601e-28 wb1 = 3.991212957e-36 pb1 = -1.018437773e-42
+ keta = 2.069517876e+00 lketa = -5.312827901e-07 wketa = -1.159976167e-06 pketa = 2.959911186e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.648749876e-01 lpclm = -1.125376359e-08 wpclm = -2.457088828e-08 ppclm = 6.269753561e-15
+ pdiblc1 = -6.757875588e+00 lpdiblc1 = 1.815010995e-06 wpdiblc1 = 3.962804181e-06 ppdiblc1 = -1.011188743e-12
+ pdiblc2 = 3.544868813e-02 lpdiblc2 = -8.729764817e-09 wpdiblc2 = -1.906013504e-08 ppdiblc2 = 4.863574658e-15
+ pdiblcb = 4.020165187e+01 lpdiblcb = -1.054891009e-05 wpdiblcb = -2.303196088e-05 ppdiblcb = 5.877065457e-12
+ drout = 1.000000238e+00 ldrout = -5.423936678e-14 wdrout = -8.494815518e-15 pdrout = 2.167621638e-21
+ pscbe1 = 5.236991324e+07 lpscbe1 = 1.907727693e+02 wpscbe1 = 4.165236915e+02 ppscbe1 = -1.062843504e-4
+ pscbe2 = 1.617158566e-07 lpscbe2 = -3.994974529e-14 wpscbe2 = -8.722427193e-14 ppscbe2 = 2.225701747e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = -5.692925215e+00 lbeta0 = 3.584340091e-06 wbeta0 = 7.825867672e-06 pbeta0 = -1.996926654e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 5.567352337e-08 lagidl = -1.394202609e-14 wagidl = -2.563275443e-14 pagidl = 6.540709947e-21
+ bgidl = 1.000000357e+09 lbgidl = -7.996280289e-05 wbgidl = 6.591606140e-06 pbgidl = -1.681980133e-12
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -2.8385e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.489374835e-02 lkt1 = -1.433535605e-07 wkt1 = -3.129911509e-07 pkt1 = 7.986595197e-14
+ kt2 = -1.697285524e+00 lkt2 = 4.201372749e-07 wkt2 = 9.173065039e-07 pkt2 = -2.340691006e-13
+ at = 1.474250203e+06 lat = -3.715199153e-01 wat = -8.111579164e-01 pat = 2.069831655e-7
+ ute = 1.195125946e+01 lute = -3.172913790e-06 wute = -6.927580906e-06 pute = 1.767710820e-12
+ ua1 = 1.564203964e-08 lua1 = -3.902074811e-15 wua1 = -8.519593484e-15 pua1 = 2.173944669e-21
+ ub1 = -2.084245651e-17 lub1 = 5.289313391e-24 wub1 = 1.154842100e-23 pub1 = -2.946810587e-30
+ uc1 = -4.991354789e-10 luc1 = 1.198876641e-16 wuc1 = 2.617567115e-16 puc1 = -6.679246007e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.171 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.143603+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43165561
+ k2 = 0.046387026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
+ voff = {-0.16725342+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.5720692+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.00827017
+ ua = -7.4124916e-10
+ ub = 6.3364395e-19
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = 5.7286e-9
+ b1 = 3.5674e-8
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.172 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.136052763e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.514439310e-7
+ k1 = 4.169789897e-01 lk1 = 2.943861458e-7
+ k2 = 6.562039979e-02 lk2 = -3.857862811e-7
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.172472591e-06 lcit = 1.303205335e-10 wcit = 1.355252716e-26 pcit = -8.131516294e-32
+ voff = {-1.346023867e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.549199771e-7
+ nfactor = {1.621526756e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -9.920280577e-07 wnfactor = 7.105427358e-21
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 6.971914874e-03 lu0 = 2.604062203e-8
+ ua = -7.228111739e-10 lua = -3.698322591e-16
+ ub = 2.485336107e-19 lub = 7.724608655e-24
+ uc = -1.046491178e-10 luc = -2.033642163e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.297654578e+04 lvsat = -2.571566868e-1
+ a0 = 1.627231194e+00 la0 = -3.274119030e-6
+ ags = 1.127413528e-01 lags = 1.100485920e-8
+ a1 = 0.0
+ a2 = 1.084157408e+00 la2 = -2.289788703e-6
+ b0 = 1.075896438e-07 lb0 = -2.043146133e-12 wb0 = -7.940933881e-29 pb0 = 1.905824131e-33
+ b1 = 5.694535280e-08 lb1 = -4.266644107e-13
+ keta = 3.426055353e-02 lketa = -2.186199026e-7
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -6.958323949e-02 lpclm = 1.696584997e-06 ppclm = -1.776356839e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 1.912368050e-03 lpdiblc2 = -1.274113513e-08 ppdiblc2 = 5.551115123e-29
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 8.855588799e-09 lpscbe2 = 2.417082098e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.715141667e-11 lalpha0 = 1.346934531e-15
+ alpha1 = -6.715141667e-11 lalpha1 = 1.346934531e-15
+ beta0 = 4.813088250e+01 lbeta0 = -3.636723234e-04 wbeta0 = 2.273736754e-19
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.815887098e-09 lagidl = -1.836585614e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.444180322e-01 lkt1 = 1.237194387e-7
+ kt2 = -6.525229044e-02 lkt2 = 1.345159137e-7
+ at = 7.718690531e+04 lat = -1.242985802e-1
+ ute = 5.651519091e-01 lute = -1.300034001e-05 wute = 8.881784197e-22 pute = 7.105427358e-27
+ ua1 = 3.782821288e-09 lua1 = -3.395088554e-14 pua1 = -1.058791184e-34
+ ub1 = -2.655052084e-18 lub1 = 2.860600094e-23 wub1 = -6.162975822e-39 pub1 = -4.930380658e-44
+ uc1 = -9.472964564e-11 luc1 = 1.302590510e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.173 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.150668308e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.366938589e-8
+ k1 = 4.604697380e-01 lk1 = -5.606969765e-8
+ k2 = 1.430285893e-02 lk2 = 2.773918708e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.322146530e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.316562590e-7
+ nfactor = {8.355552889e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.341463636e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 9.316969502e-03 lu0 = 7.143773174e-9
+ ua = -9.431379082e-10 lua = 1.405598021e-15
+ ub = 1.281825696e-18 lub = -6.018346318e-25
+ uc = -1.070056741e-10 luc = -1.346889891e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.346148460e+04 lvsat = -1.931930625e-2
+ a0 = 1.168757490e+00 la0 = 4.203400132e-7
+ ags = 4.417072978e-02 lags = 5.635585964e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = -1.140830747e-07 lb0 = -2.568696835e-13
+ b1 = 9.055190034e-09 lb1 = -4.075733774e-14 pb1 = 1.058791184e-34
+ keta = 7.543931899e-03 lketa = -3.332823646e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -4.156864620e-01 lpclm = 4.485543601e-06 wpclm = -8.881784197e-22
+ pdiblc1 = 0.39
+ pdiblc2 = 2.310096564e-04 lpdiblc2 = 8.075366429e-10
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.465883797e-08 lpscbe2 = -2.259274738e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.014542500e-10 lalpha0 = -8.175355937e-16
+ alpha1 = 2.014542500e-10 lalpha1 = -8.175355937e-16
+ beta0 = -2.439264750e+01 lbeta0 = 2.207346103e-04 wbeta0 = -2.842170943e-20 pbeta0 = 2.273736754e-25
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 6.959945019e-10 lagidl = -1.283401221e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.136586484e-01 lkt1 = -1.241449055e-7
+ kt2 = -3.842712868e-02 lkt2 = -8.164580001e-8
+ at = 2.196300907e+04 lat = 3.207049638e-1
+ ute = -1.925921477e+00 lute = 7.073152815e-6
+ ua1 = -2.987663864e-09 lua1 = 2.060683480e-14 wua1 = 6.617444900e-30 pua1 = -2.646977960e-35
+ ub1 = 2.948102001e-18 lub1 = -1.654516721e-23
+ uc1 = 5.590315313e-10 luc1 = -3.965528193e-15 wuc1 = -4.135903063e-31 puc1 = 1.654361225e-36
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.174 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.155676044e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -1.334714119e-8
+ k1 = 3.842913476e-01 lk1 = 2.530751608e-7
+ k2 = 4.432685200e-02 lk2 = -9.410328086e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.687254897e-01 ldsub = -1.252860521e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.037637994e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.619785835e-8
+ nfactor = {2.243457684e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.720436259e-7
+ eta0 = 1.618122575e-01 leta0 = -3.320080490e-7
+ etab = -1.415214075e-01 letab = 2.902460303e-7
+ u0 = 1.216753903e-02 lu0 = -4.424322556e-09 wu0 = -5.551115123e-23
+ ua = -2.772390642e-10 lua = -1.296732691e-15
+ ub = 8.233204951e-19 lub = 1.258857421e-24
+ uc = -1.342621486e-10 luc = 1.092645171e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.432087493e+04 lvsat = -1.039702583e-1
+ a0 = 1.402964339e+00 la0 = -5.301111964e-7
+ ags = -4.821423619e-02 lags = 9.384724937e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = -2.208073870e-07 lb0 = 1.762357191e-13
+ b1 = -1.625453795e-09 lb1 = 2.586530631e-15
+ keta = 2.308642681e-02 lketa = -6.640691024e-08 pketa = 1.110223025e-28
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.045581146e-01 lpclm = 3.452176679e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 4.183469811e-04 lpdiblc2 = 4.728993188e-11
+ pdiblcb = -4.308170000e-01 lpdiblcb = 8.352403749e-7
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 8.705986359e-09 lpscbe2 = 1.564936435e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.029085000e-10 lalpha0 = 4.176201874e-16
+ alpha1 = -1.029085000e-10 lalpha1 = 4.176201874e-16
+ beta0 = 5.514271247e+01 lbeta0 = -1.020334014e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -8.125329299e-11 lagidl = 1.870802463e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.353792873e-01 lkt1 = -3.599886016e-8
+ kt2 = -6.329111093e-02 lkt2 = 1.925646684e-8
+ at = 1.637106726e+05 lat = -2.545311518e-1
+ ute = -8.998158855e-02 lute = -3.774033634e-7
+ ua1 = 2.900604437e-09 lua1 = -3.288758976e-15
+ ub1 = -1.918105286e-18 lub1 = 3.202729218e-24 pub1 = 1.232595164e-44
+ uc1 = -8.850008756e-10 luc1 = 1.894600800e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.175 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.166873031e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 9.698160864e-9
+ k1 = 5.064385921e-01 lk1 = 1.675366545e-9
+ k2 = -1.550530049e-03 lk2 = 3.201705484e-10
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.600000206e-01 ldsub = -2.177893776e-14
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.008592856e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.021987531e-8
+ nfactor = {2.582745438e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.070355502e-6
+ eta0 = -5.174742150e-01 leta0 = 1.066078990e-06 weta0 = 1.457167720e-22 peta0 = 7.910339050e-28
+ etab = 2.904247369e-04 letab = -1.626828481e-9
+ u0 = 1.299481844e-02 lu0 = -6.127004236e-9
+ ua = -2.335251343e-10 lua = -1.386703390e-15
+ ub = 1.100219537e-18 lub = 6.889521208e-25
+ uc = -1.209494201e-10 luc = 8.186465865e-17 wuc = 4.135903063e-31
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.474998785e+04 lvsat = 3.921845435e-2
+ a0 = 1.027063579e+00 la0 = 2.435564714e-7
+ ags = 2.421456228e-01 lags = 3.408625427e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = -3.571202000e-08 lb0 = -2.047220124e-13
+ b1 = -8.958356404e-10 lb1 = 1.084852434e-15 wb1 = -3.308722450e-30
+ keta = -1.779393475e-02 lketa = 1.773182353e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.249152049e-01 lpclm = -3.141316846e-7
+ pdiblc1 = 3.959901522e-01 lpdiblc1 = -1.232875161e-8
+ pdiblc2 = 4.533060379e-04 lpdiblc2 = -2.466175011e-11
+ pdiblcb = 1.866340000e-01 lpdiblcb = -4.355787498e-07 wpdiblcb = -2.220446049e-22 ppdiblcb = -6.661338148e-28
+ drout = 3.733753506e-01 ldrout = 3.841052546e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 9.779790288e-09 lpscbe2 = -6.451345974e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.611938067e+00 lbeta0 = 1.967522498e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 3.976755324e-10 lagidl = 8.850855221e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.251515120e-01 lkt1 = -5.704936050e-8
+ kt2 = -5.962353039e-02 lkt2 = 1.170796260e-8
+ at = 2.764051955e+04 lat = 2.552435502e-2
+ ute = 5.465304861e-01 lute = -1.687453420e-06 pute = 1.776356839e-27
+ ua1 = 3.136618649e-09 lua1 = -3.774516346e-15 wua1 = -6.617444900e-30
+ ub1 = -1.649671782e-18 lub1 = 2.650247432e-24 wub1 = 3.081487911e-39
+ uc1 = 2.307099871e-12 luc1 = 6.837014368e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.176 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.186764098e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.074629071e-8
+ k1 = 5.895983608e-01 lk1 = -8.632180590e-8
+ k2 = -4.236429828e-02 lk2 = 4.350807568e-08 wk2 = -4.163336342e-23 pk2 = 4.163336342e-29
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -5.660916000e-01 ldsub = 8.741453484e-07 pdsub = -8.881784197e-28
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.251342609e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 3.590692590e-8
+ nfactor = {3.163637012e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.685037539e-6
+ eta0 = 1.027885506e+00 leta0 = -5.691743056e-7
+ etab = -1.522680668e-03 letab = 2.917452658e-10
+ u0 = 7.157921276e-03 lu0 = 4.942524115e-11
+ ua = -2.676735973e-09 lua = 1.198629023e-15
+ ub = 3.551846133e-18 lub = -1.905285595e-24
+ uc = -3.828526639e-11 luc = -5.608068851e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -7.419646049e+02 lvsat = 5.561157368e-2
+ a0 = 1.416791016e+00 la0 = -1.688414103e-7
+ ags = -2.012374473e-01 lags = 8.100372059e-07 pags = -1.776356839e-27
+ a1 = 0.0
+ a2 = 1.143658537e+00 la2 = -3.636491546e-7
+ b0 = -3.936436742e-07 lb0 = 1.740305261e-13
+ b1 = 3.566568533e-09 lb1 = -3.637129790e-15 pb1 = 3.308722450e-36
+ keta = 4.640102772e-02 lketa = -5.019735991e-08 wketa = -2.775557562e-23 pketa = 8.673617380e-29
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 8.463474809e-01 lpclm = -2.309936761e-7
+ pdiblc1 = 7.353910455e-01 lpdiblc1 = -3.714725948e-7
+ pdiblc2 = 1.290151741e-05 lpdiblc2 = 4.413611013e-10
+ pdiblcb = -0.225
+ drout = 9.868614715e-01 ldrout = -2.650673539e-7
+ pscbe1 = 1.538699225e+09 lpscbe1 = -7.816693584e+2
+ pscbe2 = -6.786262656e-08 lpscbe2 = 8.151374164e-14 wpscbe2 = 1.058791184e-28 ppscbe2 = -2.646977960e-35
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 4.271197094e+00 lbeta0 = 2.328084373e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.592126185e-09 lagidl = -3.788463250e-16
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.736892727e-01 lkt1 = -5.688158284e-9
+ kt2 = -3.629638816e-02 lkt2 = -1.297611950e-8
+ at = 2.023824718e+04 lat = 3.335721757e-2
+ ute = -1.951903787e+00 lute = 9.563147749e-7
+ ua1 = -2.770257084e-09 lua1 = 2.475962349e-15 wua1 = -3.308722450e-30 pua1 = 3.308722450e-36
+ ub1 = 2.776470114e-18 lub1 = -2.033363139e-24 wub1 = 6.162975822e-39
+ uc1 = 2.168072778e-10 luc1 = -1.586075096e-16 wuc1 = 4.135903063e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.177 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.198442244e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.726468175e-8
+ k1 = 2.587759691e-01 lk1 = 9.833332850e-8
+ k2 = 1.264619903e-01 lk2 = -5.072569381e-08 wk2 = 2.220446049e-22 pk2 = -1.110223025e-28
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.265530550e+00 ldsub = -1.482111871e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.432797432e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -9.781810251e-9
+ nfactor = {-1.369102099e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 8.450014502e-07 wnfactor = 8.881784197e-22 pnfactor = 1.776356839e-27
+ eta0 = -5.857710121e-01 leta0 = 3.315203530e-07 weta0 = 3.885780586e-22 peta0 = -3.747002708e-28
+ etab = -2.144165608e-03 letab = 6.386395146e-10
+ u0 = 9.588264965e-03 lu0 = -1.307119696e-9
+ ua = -4.524496467e-10 lua = -4.290087548e-17
+ ub = 1.800632172e-19 lub = -2.325752460e-26
+ uc = -1.066909176e-10 luc = 3.257391349e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.745291629e+03 lvsat = 5.087424187e-2
+ a0 = 1.730312949e+00 la0 = -3.438399480e-7
+ ags = 9.336688757e-01 lags = 1.765665437e-7
+ a1 = 0.0
+ a2 = 1.175865985e-01 la2 = 2.090734196e-7
+ b0 = -1.827582555e-07 lb0 = 5.632061198e-14
+ b1 = -6.585512924e-09 lb1 = 2.029457517e-15
+ keta = -5.806135818e-02 lketa = 8.110410026e-9
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.801832138e-01 lpclm = 1.408392328e-7
+ pdiblc1 = -3.427765615e-01 lpdiblc1 = 2.303282184e-7
+ pdiblc2 = -8.777845214e-03 lpdiblc2 = 5.348092205e-09 wpdiblc2 = 6.938893904e-24 ppdiblc2 = -3.469446952e-30
+ pdiblcb = -1.473166890e-01 lpdiblcb = -4.336049373e-8
+ drout = 4.913817236e-01 ldrout = 1.149457697e-8
+ pscbe1 = -6.773655310e+08 lpscbe1 = 4.552715062e+02 wpscbe1 = 9.536743164e-13 ppscbe1 = -2.384185791e-19
+ pscbe2 = 1.636367297e-07 lpscbe2 = -4.770225404e-14
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.865441218e+00 lbeta0 = 3.218851306e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.041584712e-09 lagidl = -6.297205910e-16
+ bgidl = 7.033052157e+08 lbgidl = 1.656061277e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.00081386752815302
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207367379934e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.360991252e-01 lkt1 = -2.666985086e-8
+ kt2 = -6.784093954e-02 lkt2 = 4.631102743e-9
+ at = 9.493059464e+04 lat = -8.333810011e-3
+ ute = 4.960630988e-01 lute = -4.100669019e-07 pute = 4.440892099e-28
+ ua1 = 3.355066581e-09 lua1 = -9.430095617e-16
+ ub1 = -1.725764093e-18 lub1 = 4.796489289e-25
+ uc1 = -2.970663052e-11 luc1 = -2.101084137e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.178 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.239991813e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 5.006901243e-8
+ k1 = -1.102372845e+00 lk1 = 5.177985587e-7
+ k2 = 4.847969085e-01 lk2 = -1.611537656e-07 wk2 = 4.440892099e-22 pk2 = 1.110223025e-28
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.977511515e+00 ldsub = -3.676223612e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-3.638620714e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 5.819504583e-8
+ nfactor = {2.927995871e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -4.792352313e-7
+ eta0 = 4.900000008e-01 leta0 = -9.356071473e-17
+ etab = 2.581819860e-03 letab = -8.177674270e-10 wetab = -1.734723476e-24 petab = -1.734723476e-30
+ u0 = 1.290521855e-02 lu0 = -2.329305283e-9
+ ua = 2.912788267e-09 lua = -1.079966243e-15
+ ub = -2.678685290e-18 lub = 8.577230029e-25 pub = -1.155557967e-45
+ uc = 4.100502134e-11 luc = -1.294154402e-17 puc = 2.261821987e-38
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.107233529e+05 lvsat = -1.041285073e-1
+ a0 = -2.787929715e-01 la0 = 2.753062236e-7
+ ags = 2.379753986e+00 lags = -2.690735049e-7
+ a1 = 0.0
+ a2 = 9.570523633e-01 la2 = -4.962474518e-8
+ b0 = -4.369331260e-14 lb0 = 1.383167812e-20 wb0 = -2.524354897e-35 pb0 = -1.893266173e-41
+ b1 = -1.379167911e-17 lb1 = 3.284876207e-24
+ keta = -9.702710173e-02 lketa = 2.011848322e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.931004364e-01 lpclm = -1.722646764e-8
+ pdiblc1 = 5.732445572e-01 lpdiblc1 = -5.196200978e-8
+ pdiblc2 = 3.354825457e-02 lpdiblc2 = -7.695541966e-9
+ pdiblcb = 2.607591983e+00 lpdiblcb = -8.923406993e-07 ppdiblcb = 8.881784197e-28
+ drout = -1.074947477e+00 ldrout = 4.941902469e-7
+ pscbe1 = 7.998824354e+08 lpscbe1 = 2.800036250e-2
+ pscbe2 = 2.140020980e-08 lpscbe2 = -3.869225705e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.080169809e+01 lbeta0 = -5.829811493e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -3.530736764e-09 lagidl = 1.087501718e-15 wagidl = -1.137373342e-30 pagidl = -7.754818243e-37
+ bgidl = 2.059624081e+09 lbgidl = -2.523706570e+2
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.00081386752815302
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207367379934e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.047221533e-01 lkt1 = -6.715629230e-8
+ kt2 = -5.971042874e-02 lkt2 = 2.125523229e-9
+ at = 2.366743202e+05 lat = -5.201497393e-02 wat = 9.313225746e-16
+ ute = -2.029992490e+00 lute = 3.683876490e-7
+ ua1 = 1.080932106e-10 lua1 = 5.761022195e-17
+ ub1 = -3.579906755e-19 lub1 = 5.814219486e-26
+ uc1 = -3.312416379e-10 luc1 = 7.191320187e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.179 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -3.7585e-8
+ vth0 = {-5.047112983e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.261595230e-05 wvth0 = 2.288520881e-05 pvth0 = -5.839618733e-12
+ k1 = -3.554095183e-01 lk1 = 3.641551384e-07 wk1 = 7.416097493e-07 pk1 = -1.892365597e-13
+ k2 = -2.492928582e+01 lk2 = 6.312254958e-06 wk2 = 1.146684292e-05 pk2 = -2.925994308e-12
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 5.655408957e+00 ldsub = -1.332351449e-06 wdsub = -1.915462703e-06 pdsub = 4.887686180e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-7.392059876e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.883182137e-05 wvoff = 3.432596140e-05 pvoff = -8.758955570e-12
+ nfactor = {2.321454864e+02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -5.900286895e-05 wnfactor = -1.106642405e-04 pnfactor = 2.823819424e-11
+ eta0 = 8.967739560e+00 leta0 = -2.163264803e-06 weta0 = -2.890227681e-06 peta0 = 7.374993975e-13
+ etab = 4.851421498e-01 letab = -1.240110571e-07 wetab = -1.662649903e-07 petab = 4.242583758e-14
+ u0 = 6.759426426e-01 lu0 = -1.716828250e-07 wu0 = -3.076105723e-07 pu0 = 7.849298973e-14
+ ua = 1.430032198e-07 lua = -3.690392705e-14 wua = -6.415649765e-14 pua = 1.637081351e-20
+ ub = -1.302410537e-17 lub = 3.558786044e-24 wub = 2.737303243e-24 pub = -6.984776685e-31
+ uc = -5.030527678e-10 luc = 1.249619459e-16 wuc = 1.818700145e-16 puc = -4.640777160e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.114750179e+07 lvsat = -1.558424770e+01 wvsat = -2.873137341e+01 pvsat = 7.331384553e-6
+ a0 = -3.111422112e-01 la0 = 3.032114732e-07 wa0 = 7.796566293e-08 pa0 = -1.989449821e-14
+ ags = 1.249999929e+00 lags = 2.020171053e-14 wags = 6.699724509e-14 pags = -1.709568664e-20
+ a1 = 0.0
+ a2 = -7.363872496e+00 la2 = 2.070083557e-06 wa2 = 3.058897389e-06 pa2 = -7.805388467e-13
+ b0 = -4.992672238e-05 lb0 = 1.273980175e-11 wb0 = 2.331188512e-11 pb0 = -5.948493727e-18
+ b1 = 3.999570915e-21 lb1 = -9.005834523e-28 wb1 = -1.079595847e-33 pb1 = 2.754804722e-40
+ keta = -1.598144941e+00 lketa = 4.045947310e-07 wketa = 5.525362907e-07 pketa = -1.409906853e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 6.663560035e-01 lpclm = -1.163167441e-08 wpclm = -2.526240718e-08 ppclm = 6.446208440e-15
+ pdiblc1 = 1.551553496e+00 lpdiblc1 = -3.053060247e-07 wpdiblc1 = 8.294893393e-08 ppdiblc1 = -2.116607947e-14
+ pdiblc2 = 2.687923105e-02 lpdiblc2 = -6.543096453e-09 wpdiblc2 = -1.505886700e-08 ppdiblc2 = 3.842571092e-15
+ pdiblcb = -1.788329392e+01 lpdiblcb = 4.272625531e-06 wpdiblcb = 4.089178185e-06 ppdiblcb = -1.043435598e-12
+ drout = 1.000000074e+00 ldrout = -1.220824686e-14 wdrout = 6.841568734e-14 pdrout = -1.745763001e-20
+ pscbe1 = 1.335209438e+09 lpscbe1 = -1.365693924e+02 wpscbe1 = -1.824623053e+02 ppscbe1 = 4.655890645e-5
+ pscbe2 = -1.925410871e-08 lpscbe2 = 6.228360753e-15 wpscbe2 = -2.725413796e-15 ppscbe2 = 6.954438383e-22
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.897858558e+01 lbeta0 = -2.711089319e-06 wbeta0 = -3.693803493e-06 pbeta0 = 9.425478374e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -3.661321268e-07 lagidl = 9.369012167e-14 wagidl = 1.713175834e-13 pagidl = -4.371510775e-20
+ bgidl = 1.000000471e+09 lbgidl = -1.090464325e-04 wbgidl = -4.662698364e-05 pbgidl = 1.189780426e-11
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -2.8385e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 3.219943884e-01 lkt1 = -2.318690064e-07 wkt1 = -4.749608535e-07 pkt1 = 1.211957610e-13
+ kt2 = 1.168718090e+00 lkt2 = -3.111808672e-07 wkt2 = -4.208936354e-07 pkt2 = 1.073994290e-13
+ at = -6.408211581e+05 lat = 1.681828439e-01 wat = 1.764154336e-01 pat = -4.501592619e-8
+ ute = -2.885438840e+00 lute = 6.129665157e-07 wute = -6.072284009e-14 pute = 1.549464557e-20
+ ua1 = -5.692061196e-10 lua1 = 2.345487707e-16 wua1 = -9.502061899e-16 pua1 = 2.424641135e-22
+ ub1 = 4.254339820e-18 lub1 = -1.114636128e-24 wub1 = -1.698253339e-25 pub1 = 4.333433045e-32
+ uc1 = -7.791755265e-10 luc1 = 1.913454831e-16 wuc1 = 3.925135706e-16 puc1 = -1.001576878e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.180 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 4.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.143603+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43165561
+ k2 = 0.046387026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
+ voff = {-0.16725342+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.5720692+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.00827017
+ ua = -7.4124916e-10
+ ub = 6.3364395e-19
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = 5.7286e-9
+ b1 = 3.5674e-8
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.181 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 4.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.209193806e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.315631539e-06 wvth0 = 3.341975154e-08 pvth0 = -6.703390577e-13
+ k1 = 3.754552419e-01 lk1 = 1.127276537e-06 wk1 = 1.897311385e-08 pk1 = -3.805659431e-13
+ k2 = 8.667148822e-02 lk2 = -8.080325915e-07 wk2 = -9.618705427e-09 pk2 = 1.929336286e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.172472591e-06 lcit = 1.303205335e-10 wcit = -8.470329473e-28 pcit = -5.929230631e-33
+ voff = {-1.288670968e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -7.699593968e-07 wvoff = -2.620580129e-09 pvoff = 5.256404174e-14
+ nfactor = {1.985534167e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -8.293350606e-06 wnfactor = -1.663229946e-07 pnfactor = 3.336134902e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.038204571e-02 lu0 = -4.236036209e-08 wu0 = -1.558163804e-09 pu0 = 3.125391447e-14
+ ua = -7.876854956e-10 lua = 9.314279145e-16 wua = 2.964250483e-17 pua = -5.945744011e-22
+ ub = 8.645053103e-19 lub = -4.630656411e-24 wub = -2.814510209e-25 pub = 5.645392425e-30
+ uc = -1.098054016e-10 luc = 8.308919582e-17 wuc = 2.356019516e-18 puc = -4.725743998e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.289725785e+05 lvsat = -9.791712305e-01 wvsat = -1.644737926e-02 pvsat = 3.299043293e-7
+ a0 = 1.957702634e+00 la0 = -9.902771362e-06 wa0 = -1.509996715e-07 pa0 = 3.028777081e-12
+ ags = 1.345421664e-01 lags = -4.262795666e-07 wags = -9.961271362e-09 pags = 1.998048744e-13
+ a1 = 0.0
+ a2 = 1.404675261e+00 la2 = -8.718790282e-06 wa2 = -1.464516583e-07 pa2 = 2.937552259e-12
+ b0 = -4.048960415e-08 lb0 = 9.270525959e-13 wb0 = 6.766066614e-14 pb0 = -1.357149144e-18
+ b1 = 3.136852434e-07 lb1 = -5.576396783e-12 wb1 = -1.173101043e-13 pb1 = 2.353026015e-18
+ keta = 6.678954219e-02 lketa = -8.710918870e-07 wketa = -1.486321056e-08 pketa = 2.981288041e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -3.025368140e-01 lpclm = 6.369207396e-06 wpclm = 1.064416132e-07 ppclm = -2.135023972e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 7.107520204e-03 lpdiblc2 = -1.169463802e-07 wpdiblc2 = -2.373779312e-09 ppdiblc2 = 4.761366899e-14
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 5.361370337e+08 lpscbe1 = 5.292608234e+03 wpscbe1 = 1.205647943e+02 ppscbe1 = -2.418309140e-3
+ pscbe2 = 4.807968877e-09 lpscbe2 = 1.053586695e-13 wpscbe2 = 1.849446590e-15 ppscbe2 = -3.709651410e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -2.556913301e-10 lalpha0 = 5.128700166e-15 walpha0 = 8.614803430e-17 palpha0 = -1.727971917e-21
+ alpha1 = -2.556913301e-10 lalpha1 = 5.128700166e-15 walpha1 = 8.614803430e-17 palpha1 = -1.727971917e-21
+ beta0 = 9.903665911e+01 lbeta0 = -1.384749045e-03 wbeta0 = -2.325996926e-05 pbeta0 = 4.665524177e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 3.218243378e-09 lagidl = -2.643638680e-14 wagidl = -1.838454359e-16 pagidl = 3.687603007e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.895471207e-01 lkt1 = 3.034743368e-06 wkt1 = 6.631267339e-08 pkt1 = -1.330110876e-12
+ kt2 = -7.217324940e-02 lkt2 = 2.733376851e-07 wkt2 = 3.162338411e-09 pkt2 = -6.343072145e-14
+ at = -2.040464011e+04 lat = 1.833209228e+00 wat = 4.459172412e-02 pat = -8.944283829e-7
+ ute = 5.882665254e-01 lute = -1.346397692e-05 wute = -1.056157671e-08 pute = 2.118459011e-13
+ ua1 = 5.510005249e-09 lua1 = -6.859503505e-14 wua1 = -7.891883500e-16 pua1 = 1.582967409e-20
+ ub1 = -4.855417607e-18 lub1 = 7.274130667e-23 wub1 = 1.005395416e-24 pub1 = -2.016639216e-29
+ uc1 = -1.225897776e-10 luc1 = 1.861413774e-15 wuc1 = 1.272990723e-17 puc1 = -2.553386432e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.182 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 4.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.046333694e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 3.277067664e-09 wvth0 = -4.767278067e-08 pvth0 = -1.688164745e-14
+ k1 = 5.142563750e-01 lk1 = 8.793409904e-09 wk1 = -2.457629777e-08 pk1 = -2.963738083e-14
+ k2 = -1.182757966e-02 lk2 = -1.431035765e-08 wk2 = 1.193957227e-08 pk2 = 1.921336208e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.510046953e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.142461354e-07 wvoff = 8.585583708e-09 pvoff = -3.773713151e-14
+ nfactor = {-9.594631276e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.543793825e-05 wnfactor = 8.201834049e-07 pnfactor = -4.613301372e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 5.096172851e-03 lu0 = 2.341000404e-10 wu0 = 1.928574847e-09 pu0 = 3.157181668e-15
+ ua = -1.867734404e-09 lua = 9.634645630e-15 wua = 4.224684803e-16 pua = -3.760032892e-21
+ ub = 2.144848073e-18 lub = -1.494787605e-23 wub = -3.943339105e-25 pub = 6.555021939e-30
+ uc = -9.090883925e-11 luc = -6.918251592e-17 wuc = -7.354997985e-18 puc = 3.099558992e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -5.560395780e+04 lvsat = 5.081778771e-01 wvsat = 5.440362007e-02 pvsat = -2.410250680e-7
+ a0 = 1.405933495e-01 la0 = 4.739804161e-06 wa0 = 4.697908155e-07 pa0 = -1.973658197e-12
+ ags = 7.385913981e-03 lags = 5.983671320e-07 wags = 1.680779160e-08 pags = -1.590478572e-14
+ a1 = 0.0
+ a2 = -1.615535583e-01 la2 = 3.902147804e-06 wa2 = 4.393549749e-07 pa2 = -1.782977179e-12
+ b0 = 3.650489666e-07 lb0 = -2.340846149e-12 wb0 = -2.189259706e-13 pb0 = 9.522146944e-19
+ b1 = -7.301510286e-07 lb1 = 2.835013349e-12 wb1 = 3.377595838e-13 pb1 = -1.314002894e-18
+ keta = -7.032600481e-02 lketa = 2.338085004e-07 wketa = 3.558048722e-08 pketa = -1.083550881e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -7.040557399e-01 lpclm = 9.604715160e-06 wpclm = 1.317622672e-07 ppclm = -2.339062107e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -1.493130810e-02 lpdiblc2 = 6.064624489e-08 wpdiblc2 = 6.927996555e-09 ppdiblc2 = -2.734162225e-14
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 1.591588899e+09 lpscbe1 = -3.212402321e+03 wpscbe1 = -3.616943828e+02 ppscbe1 = 1.467817294e-3
+ pscbe2 = 2.811198116e-08 lpscbe2 = -8.242902320e-14 wpscbe2 = -6.147037094e-15 ppscbe2 = 2.734051082e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.670739902e-10 lalpha0 = -3.112916655e-15 walpha0 = -2.584441029e-16 palpha0 = 1.048810105e-21
+ alpha1 = 7.670739902e-10 lalpha1 = -3.112916655e-15 walpha1 = -2.584441029e-16 palpha1 = 1.048810105e-21
+ beta0 = -1.771099773e+02 lbeta0 = 8.404874967e-04 wbeta0 = 6.977990779e-05 pbeta0 = -2.831787284e-10
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.606115054e-09 lagidl = -2.150375270e-14 wagidl = -8.727761029e-16 pagidl = 9.239123440e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 9.578998301e-02 lkt1 = -2.487819521e-06 wkt1 = -2.327782875e-07 pkt1 = 1.080014933e-12
+ kt2 = -1.766425180e-02 lkt2 = -1.659050841e-07 wkt2 = -9.487015234e-09 pkt2 = 3.849992061e-14
+ at = 2.292822233e+05 lat = -1.788099636e-01 wat = -9.472871000e-02 pat = 2.282393596e-7
+ ute = -1.824354482e+00 lute = 5.977333305e-06 wute = -4.640819458e-08 pute = 5.007040418e-13
+ ua1 = -8.169215747e-09 lua1 = 4.163445320e-14 wua1 = 2.367565050e-15 pua1 = -9.607981458e-21
+ ub1 = 9.549198571e-18 lub1 = -4.333353928e-23 wub1 = -3.016186247e-24 pub1 = 1.224019654e-29
+ uc1 = 1.748835214e-09 luc1 = -1.321884695e-14 wuc1 = -5.436474784e-16 puc1 = 4.228044914e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.183 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 4.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-9.168434063e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -5.222165322e-07 wvth0 = -1.091278866e-07 pvth0 = 2.325136199e-13
+ k1 = 4.235316687e-01 lk1 = 3.769696913e-07 wk1 = -1.792976601e-08 pk1 = -5.661013664e-14
+ k2 = 6.986078642e-02 lk2 = -3.458156343e-07 wk2 = -1.166701638e-08 pk2 = 1.150129119e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.687254608e-01 ldsub = -1.252860403e-06 wdsub = 1.320205212e-14 pdsub = -5.357617150e-20
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-5.310124969e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -5.888796904e-07 wvoff = -6.884103352e-08 pvoff = 2.764732437e-13
+ nfactor = {3.475899239e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -2.561516247e-06 wnfactor = -5.631296601e-07 pnfactor = 1.000418209e-12
+ eta0 = 1.618122575e-01 leta0 = -3.320080490e-7
+ etab = -1.415214075e-01 letab = 2.902460303e-7
+ u0 = -6.352854481e-03 lu0 = 4.669619929e-08 wu0 = 8.462375242e-09 pu0 = -2.335809108e-14
+ ua = 2.152606094e-09 lua = -6.680579572e-15 wua = -1.110249710e-15 pua = 2.459998085e-21
+ ub = -6.913737733e-18 lub = 2.181340511e-23 wub = 3.535232120e-24 pub = -9.391825038e-30
+ uc = -1.005085977e-10 luc = -3.022506433e-17 wuc = -1.542274000e-17 puc = 6.373585854e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.551965825e+05 lvsat = -3.472865516e-01 wvsat = -3.238467005e-02 pvsat = 1.111765673e-7
+ a0 = 1.719945020e+00 la0 = -1.669473406e-06 wa0 = -1.448354464e-07 pa0 = 5.205996596e-13
+ ags = -4.751785709e-01 lags = 2.556695848e-06 wags = 1.950893977e-07 pags = -7.394018513e-13
+ a1 = 0.0
+ a2 = 0.8
+ b0 = -1.545714070e-07 lb0 = -2.321383371e-13 wb0 = -3.026467644e-14 pb0 = 1.865950905e-19
+ b1 = -7.028213537e-08 lb1 = 1.571532030e-13 wb1 = 3.137074826e-14 pb1 = -7.062491306e-20
+ keta = 7.074275049e-03 lketa = -8.029499335e-08 wketa = 7.316304409e-09 pketa = 6.345770713e-15
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.181890474e+00 lpclm = -2.106945188e-06 wpclm = -7.207178564e-07 ppclm = 1.120447156e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -4.606484131e-04 lpdiblc2 = 1.921847856e-09 wpdiblc2 = 4.016323335e-10 ppdiblc2 = -8.565267560e-16
+ pdiblcb = -1.008685961e+00 lpdiblcb = 3.180330855e-06 wpdiblcb = 2.640410412e-07 ppdiblcb = -1.071523432e-12
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 5.830584491e-09 lpscbe2 = 7.992672319e-15 wpscbe2 = 1.313834372e-15 ppscbe2 = -2.936973936e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.029085000e-10 lalpha0 = 4.176201874e-16
+ alpha1 = -1.029085000e-10 lalpha1 = 4.176201874e-16
+ beta0 = 5.239738070e+01 lbeta0 = -9.089237842e-05 wbeta0 = 1.254402482e-06 pbeta0 = -5.090578521e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -3.047933694e-09 lagidl = 1.441338304e-15 wagidl = 1.355541542e-15 pagidl = 1.962316222e-22
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -8.238088261e-01 lkt1 = 1.244068778e-06 wkt1 = 1.774820017e-07 pkt1 = -5.848910655e-13
+ kt2 = -5.836477805e-02 lkt2 = -7.354294981e-10 wkt2 = -2.250949876e-09 pkt2 = 9.134737260e-15
+ at = 2.478198201e+05 lat = -2.540386828e-01 wat = -3.843131990e-02 pat = -2.250199208e-10
+ ute = -2.721753500e+00 lute = 9.619131080e-06 wute = 1.202514486e-06 pute = -4.567636511e-12
+ ua1 = 4.532716024e-10 lua1 = 6.642933715e-15 wua1 = 1.118240214e-15 pua1 = -4.538008888e-21
+ ub1 = -1.658555443e-18 lub1 = 2.149431828e-24 wub1 = -1.185940337e-25 pub1 = 4.812747496e-31
+ uc1 = -3.049438096e-09 luc1 = 6.253361847e-15 wuc1 = 9.889789837e-16 puc1 = -1.991613815e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.184 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 4.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.193281473e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 4.674000278e-08 wvth0 = 1.206659798e-08 pvth0 = -1.692523249e-14
+ k1 = 6.300045407e-01 lk1 = -4.798657961e-08 wk1 = -5.646000034e-08 pk1 = 2.269163576e-14
+ k2 = -9.922083548e-02 lk2 = 2.183087494e-09 wk2 = 4.462771130e-08 pk2 = -8.512077366e-16
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 2.458544720e+00 ldsub = -4.524978709e-06 wdsub = -1.004563441e-06 pdsub = 2.067562312e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-3.787229918e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 8.130521048e-08 wvoff = 8.126984034e-08 pvoff = -3.248045351e-14
+ nfactor = {-1.041266780e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 6.735579338e-06 wnfactor = 1.655890911e-06 pnfactor = -3.566703359e-12
+ eta0 = -1.319645909e+00 leta0 = 2.717084705e-06 weta0 = 3.665298946e-07 peta0 = -7.543808332e-13
+ etab = -2.510562138e+00 letab = 5.166134591e-06 wetab = 1.147263775e-06 petab = -2.361263883e-12
+ u0 = 2.457874415e-02 lu0 = -1.696628907e-08 wu0 = -5.292950502e-09 pu0 = 4.952707706e-15
+ ua = 1.095700303e-09 lua = -4.505287779e-15 wua = -6.073523451e-16 pua = 1.424949816e-21
+ ub = 2.510825216e-18 lub = 2.416052383e-24 wub = -6.445367681e-25 pub = -7.891501061e-31
+ uc = -2.218434558e-10 luc = 2.195027007e-16 wuc = 4.610070460e-17 puc = -6.288984945e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -1.165181303e+05 lvsat = 2.119485189e-01 wvsat = 5.997929109e-02 pvsat = -7.892416656e-8
+ a0 = 1.609084003e-01 la0 = 1.539288993e-06 wa0 = 3.957653566e-07 pa0 = -5.920486951e-13
+ ags = 1.691525206e+00 lags = -1.902748865e-06 wags = -6.622534179e-07 pags = 1.025155412e-12
+ a1 = 0.0
+ a2 = 0.8
+ b0 = -6.731763162e-08 lb0 = -4.117214400e-13 wb0 = 1.444129927e-14 pb0 = 9.458259246e-20
+ b1 = 2.695973342e-08 lb1 = -4.298709412e-14 wb1 = -1.272782233e-14 pb1 = 2.013744196e-20
+ keta = -1.028067094e-01 lketa = 1.458587525e-07 wketa = 3.884420703e-08 pketa = -5.854401262e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.047353926e+00 lpclm = 2.281238986e-07 wpclm = -5.594494554e-08 ppclm = -2.477685056e-13
+ pdiblc1 = 4.087959914e-01 lpdiblc1 = -3.868534569e-08 wpdiblc1 = -5.851269662e-09 ppdiblc1 = 1.204290768e-14
+ pdiblc2 = 5.187420120e-04 lpdiblc2 = -9.390413486e-11 wpdiblc2 = -2.989913617e-11 ppdiblc2 = 3.163836892e-17
+ pdiblcb = 1.342371921e+00 lpdiblcb = -1.658545946e-06 wpdiblcb = -5.280820824e-07 ppdiblcb = 5.588006172e-13
+ drout = 6.954239038e-01 ldrout = -2.787254161e-07 wdrout = -1.471510690e-07 pdrout = 3.028619157e-13
+ pscbe1 = 800000000.0
+ pscbe2 = 1.006754100e-08 lpscbe2 = -7.277044506e-16 wpscbe2 = -1.314796290e-16 ppscbe2 = 3.772798247e-23
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.135167652e-11 lalpha0 = 1.412899199e-16 walpha0 = 3.136692926e-17 palpha0 = -6.455847279e-23
+ alpha1 = -4.942012546e-10 lalpha1 = 1.222967196e-15 walpha1 = 2.715036256e-16 palpha1 = -5.588006172e-22
+ beta0 = 9.477026225e+00 lbeta0 = -2.554992460e-06 wbeta0 = -2.222965811e-06 pbeta0 = 2.066436580e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -6.554718001e-09 lagidl = 8.658896561e-15 wagidl = 3.176701558e-15 pagidl = -3.552025287e-21
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 1.031014157e-01 lkt1 = -6.636700741e-07 wkt1 = -2.413703842e-07 pkt1 = 2.771783497e-13
+ kt2 = -7.787172214e-02 lkt2 = 3.941317764e-08 wkt2 = 8.338000272e-09 pkt2 = -1.265912227e-14
+ at = 1.655955720e+05 lat = -8.480720209e-02 wat = -6.303469847e-02 pat = 5.041291574e-8
+ ute = 5.240992341e+00 lute = -6.769553529e-06 wute = -2.145002900e-06 pute = 2.322123346e-12
+ ua1 = 7.503912850e-09 lua1 = -7.868484582e-15 wua1 = -1.995512801e-15 pua1 = 1.870624154e-21
+ ub1 = -1.266433934e-18 lub1 = 1.342379102e-24 wub1 = -1.751098043e-25 pub1 = 5.975938133e-31
+ uc1 = 2.572646423e-11 luc1 = -7.584959596e-17 wuc1 = -1.070082280e-17 puc1 = 6.589717187e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.185 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 4.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.206918173e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.116994999e-08 wvth0 = 9.208840485e-09 pvth0 = -1.390123924e-14
+ k1 = 9.560985435e-01 lk1 = -3.930494705e-07 wk1 = -1.674619964e-07 pk1 = 1.401506180e-13
+ k2 = -2.983106602e-01 lk2 = 2.128539673e-07 wk2 = 1.169475236e-07 pk2 = -7.737786349e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -7.282584501e+00 ldsub = 5.782791999e-06 wdsub = 3.068913369e-06 pdsub = -2.242868645e-12
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-4.321243112e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.378128847e-07 wvoff = 9.457830778e-08 pvoff = -4.656307451e-14
+ nfactor = {1.284595305e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -7.959460065e-06 wnfactor = -4.424063207e-06 pnfactor = 2.866921689e-12
+ eta0 = 4.142441063e+00 leta0 = -3.062731866e-06 weta0 = -1.423108954e-06 peta0 = 1.139361307e-12
+ etab = 5.023297182e+00 letab = -2.805969325e-06 wetab = -2.295950741e-06 petab = 1.282242421e-12
+ u0 = 3.356618409e-03 lu0 = 5.490327725e-09 wu0 = 1.736898909e-09 pu0 = -2.486068045e-15
+ ua = -8.598411362e-09 lua = 5.752730362e-15 wua = 2.705743762e-15 pua = -2.080869092e-21
+ ub = 1.224438622e-17 lub = -7.883709862e-24 wub = -3.971812800e-24 pub = 2.731673573e-30
+ uc = 1.199763002e-10 luc = -1.422007106e-16 wuc = -7.231319154e-17 puc = 6.241218304e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.613515306e+04 lvsat = 8.088594048e-03 wvsat = -3.512684636e-02 pvsat = 2.171429490e-8
+ a0 = 1.322629914e+00 la0 = 3.099901387e-07 wa0 = 4.302427900e-08 pa0 = -2.187886690e-13
+ ags = -1.621080275e+00 lags = 1.602550877e-06 wags = 6.487574248e-07 pags = -3.621169318e-13
+ a1 = 0.0
+ a2 = 2.641378852e+00 la2 = -1.948491859e-06 wa2 = -6.843413614e-07 pa2 = 7.241494984e-13
+ b0 = -8.555962667e-07 lb0 = 4.224113633e-13 wb0 = 2.110763025e-13 pb0 = -1.134906689e-19
+ b1 = -8.327733484e-09 lb1 = -5.646955262e-15 wb1 = 5.434768266e-15 pb1 = 9.183334740e-22
+ keta = 1.677497041e-01 lketa = -1.404359276e-07 wketa = -5.544687991e-08 pketa = 4.123198684e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 9.563645027e-01 lpclm = 3.244061771e-07 wpclm = -5.026919765e-08 ppclm = -2.537744117e-13
+ pdiblc1 = 5.316336387e-01 lpdiblc1 = -1.686684589e-07 wpdiblc1 = 9.310124184e-08 ppdiblc1 = -9.266567141e-14
+ pdiblc2 = -2.421705404e-03 lpdiblc2 = 3.017589108e-09 wpdiblc2 = 1.112425464e-09 ppdiblc2 = -1.177135253e-15
+ pdiblcb = 1.664964306e-01 lpdiblcb = -4.142697779e-07 wpdiblcb = -1.788833320e-07 ppdiblcb = 1.892889755e-13
+ drout = 1.872395222e+00 ldrout = -1.524161156e-06 wdrout = -4.046198525e-07 pdrout = 5.753076583e-13
+ pscbe1 = 3.612732726e+09 lpscbe1 = -2.976349388e+03 wpscbe1 = -9.476715353e+02 ppscbe1 = 1.002797589e-3
+ pscbe2 = -2.837714525e-07 lpscbe2 = 3.102039033e-13 wpscbe2 = 9.865349257e-14 ppscbe2 = -1.044935661e-19
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.372966470e-10 lalpha0 = -7.663486943e-17 walpha0 = -6.273385852e-17 palpha0 = 3.501615781e-23
+ alpha1 = 1.288402509e-09 lalpha1 = -6.633306285e-16 walpha1 = -5.430072513e-16 palpha1 = 3.030903574e-22
+ beta0 = 4.657246032e+00 lbeta0 = 2.545154346e-06 wbeta0 = -1.763942528e-07 pbeta0 = -9.918404630e-14
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.696375984e-09 lagidl = -1.130333561e-15 wagidl = -5.045560266e-16 pagidl = 3.433710508e-22
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -6.316544831e-01 lkt1 = 1.138265754e-07 wkt1 = 7.217777991e-08 pkt1 = -5.460891114e-14
+ kt2 = -1.950533621e-02 lkt2 = -2.234838097e-08 wkt2 = -7.672201039e-09 pkt2 = 4.282392454e-15
+ at = 9.153492862e+04 lat = -6.438451107e-03 wat = -3.257702228e-02 pat = 1.818351652e-8
+ ute = -1.961623558e+00 lute = 8.520385367e-07 wute = 4.441176974e-09 pute = 4.764610728e-14
+ ua1 = -2.792783096e-09 lua1 = 3.027170168e-15 wua1 = 1.029263042e-17 pua1 = -2.518589792e-22
+ ub1 = 1.186277190e-18 lub1 = -1.253006228e-24 wub1 = 7.265941313e-25 pub1 = -3.565622403e-31
+ uc1 = -2.206886395e-11 luc1 = -2.527401354e-17 wuc1 = 1.091477644e-16 puc1 = -6.092300767e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.186 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 4.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.014085485e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.646347151e-08 wvth0 = -8.423665907e-08 pvth0 = 3.825723524e-14
+ k1 = 7.976885510e-01 lk1 = -3.046297650e-07 wk1 = -2.462410148e-07 pk1 = 1.841227026e-13
+ k2 = -7.941673422e-02 lk2 = 9.067394465e-08 wk2 = 9.407051856e-08 pk2 = -6.460860560e-14
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 5.480523523e+00 ldsub = -1.341192006e-06 wdsub = -1.925923019e-06 pdsub = 5.450991818e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {9.620922656e-02+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.570870461e-07 wvoff = -1.094277790e-07 pvoff = 6.730700297e-14
+ nfactor = {3.335962107e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -9.754378502e-07 wnfactor = -7.780003171e-07 pnfactor = 8.317987660e-13
+ eta0 = -3.606195353e+00 leta0 = 1.262324523e-06 weta0 = 1.380098331e-06 peta0 = -4.253049028e-13
+ etab = -8.146755628e-03 letab = 2.431737036e-09 wetab = 2.742715437e-09 petab = -8.193057055e-16
+ u0 = 1.020588157e-02 lu0 = 1.667274509e-09 wu0 = -2.822026123e-10 pu0 = -1.359066149e-15
+ ua = -2.127039694e-09 lua = 2.140604838e-15 wua = 7.651570335e-16 pua = -9.976917975e-22
+ ub = 2.144234583e-18 lub = -2.246108224e-24 wub = -8.974731088e-25 pub = 1.015669387e-30
+ uc = -2.953953041e-10 luc = 8.964725785e-17 wuc = 8.622318571e-17 puc = -2.607806665e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.651318611e+04 lvsat = 2.295887341e-03 wvsat = -3.599078388e-02 pvsat = 2.219651891e-8
+ a0 = 5.344999447e+00 la0 = -1.935175864e-06 wa0 = -1.651629784e-06 pa0 = 7.271163893e-13
+ ags = 4.551125016e-02 lags = 6.723094855e-07 wags = 4.058187586e-07 pags = -2.265158565e-13
+ a1 = 0.0
+ a2 = -4.066788929e+00 la2 = 1.795806151e-06 wa2 = 1.911933235e-06 pa2 = -7.250130929e-13
+ b0 = -2.206272252e-07 lb0 = 6.799069339e-14 wb0 = 1.730316536e-14 pb0 = -5.332316938e-21
+ b1 = -4.118098503e-08 lb1 = 1.269074415e-14 wb1 = 1.580743230e-14 pb1 = -4.871376412e-21
+ keta = -1.358841569e-01 lketa = 2.904338454e-08 wketa = 3.555894882e-08 pketa = -9.564736582e-15
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 3.303125265e+00 lpclm = -9.854852774e-07 wpclm = -1.426940928e-06 ppclm = 5.146424479e-13
+ pdiblc1 = -7.370382191e-01 lpdiblc1 = 5.394661120e-07 wpdiblc1 = 1.801468251e-07 ppdiblc1 = -1.412519046e-13
+ pdiblc2 = -1.042254405e-02 lpdiblc2 = 7.483417215e-09 wpdiblc2 = 7.514990819e-10 ppdiblc2 = -9.756769745e-16
+ pdiblcb = -7.121994124e-01 lpdiblcb = 7.619188073e-08 wpdiblcb = 2.581073438e-07 ppdiblcb = -5.462611004e-14
+ drout = -9.432183044e-01 ldrout = 4.742984606e-08 wdrout = 6.555003140e-07 pdrout = -1.641961502e-14
+ pscbe1 = -4.825448957e+09 lpscbe1 = 1.733590482e+03 wpscbe1 = 1.895350575e+03 ppscbe1 = -5.840920629e-4
+ pscbe2 = 5.979782820e-07 lpscbe2 = -1.819623460e-13 wpscbe2 = -1.984602108e-13 ppscbe2 = 6.134638975e-20
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.020224373e+01 lbeta0 = -5.498970205e-07 wbeta0 = -1.067736479e-06 pbeta0 = 3.983364441e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.163518314e-08 lagidl = -6.119707551e-15 wagidl = -4.383526180e-15 pagidl = 2.508495822e-21
+ bgidl = -1.297197852e+08 lbgidl = 6.305756925e+02 wbgidl = 3.806274495e+02 pbgidl = -2.124548235e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.746786053e-01 lkt1 = -2.960965036e-08 wkt1 = -2.806438682e-08 pkt1 = 1.343259067e-15
+ kt2 = -3.156927611e-02 lkt2 = -1.561465164e-08 wkt2 = -1.657332100e-08 pkt2 = 9.250730582e-15
+ at = 2.235172536e+05 lat = -8.010702546e-02 wat = -5.875407340e-02 pat = 3.279476115e-8
+ ute = 1.474728761e+00 lute = -1.066030237e-06 wute = -4.471738717e-07 pute = 2.997240790e-13
+ ua1 = 5.503699356e-09 lua1 = -1.603677442e-15 wua1 = -9.817575847e-16 pua1 = 3.018736894e-22
+ ub1 = -1.379831809e-18 lub1 = 1.793188322e-25 wub1 = -1.580640708e-25 pub1 = 1.372274284e-31
+ uc1 = 1.071784524e-10 luc1 = -9.741598810e-17 wuc1 = -6.254580585e-17 puc1 = 3.491119245e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.187 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 4.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.783499820e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.906469442e-07 wvth0 = 2.483407656e-07 pvth0 = -6.423314972e-14
+ k1 = -6.588632983e+00 lk1 = 1.971612942e-06 wk1 = 2.506792954e-06 pk1 = -6.642797756e-13
+ k2 = 2.205998627e+00 lk2 = -6.136225072e-07 wk2 = -7.864549316e-07 pk2 = 2.067429224e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 5.670670297e+00 ldsub = -1.399789538e-06 wdsub = -1.687485497e-06 pdsub = 4.716198906e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.132577976e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.215883061e-07 wvoff = 3.512432085e-07 pvoff = -7.465797527e-14
+ nfactor = {3.089666409e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.824776003e-06 wnfactor = -7.387082528e-08 pnfactor = 6.148071805e-13
+ eta0 = 4.900000032e-01 leta0 = -3.562510287e-16 weta0 = -1.075423306e-15 peta0 = 1.200287647e-22
+ etab = 9.848300470e-03 letab = -3.113799402e-09 wetab = -3.320214854e-09 petab = 1.049107522e-15
+ u0 = 4.439652769e-02 lu0 = -8.869256906e-09 wu0 = -1.438907195e-08 pu0 = 2.988247775e-15
+ ua = 1.816297654e-08 lua = -4.112169466e-15 wua = -6.968146527e-15 pua = 1.385480361e-21
+ ub = -1.574214568e-17 lub = 3.265937583e-24 wub = 5.968982450e-24 pub = -1.100366222e-30
+ uc = 1.554096389e-10 luc = -4.927730146e-17 wuc = -5.227398668e-17 puc = 1.660260696e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.380553063e+06 lvsat = -3.964883816e-01 wvsat = -3.974443310e-01 pvsat = 1.335856585e-7
+ a0 = -4.336198538e+00 la0 = 1.048278919e-06 wa0 = 1.853917866e-06 pa0 = -3.531882301e-13
+ ags = 5.551745424e+00 lags = -1.024546700e-06 wags = -1.449352672e-06 pags = 3.451923232e-13
+ a1 = 0.0
+ a2 = 2.373686996e+00 la2 = -1.889553151e-07 wa2 = -6.472915295e-07 pa2 = 6.366320268e-14
+ b0 = -1.663702982e-13 lb0 = 5.266665024e-20 wb0 = 5.605381359e-20 pb0 = -1.774455313e-26
+ b1 = -5.251434669e-17 lb1 = 1.250776839e-23 wb1 = 1.769323872e-23 pb1 = -4.214142340e-30
+ keta = -2.902191950e-01 lketa = 7.660481324e-08 wketa = 8.827371763e-08 pketa = -2.580984689e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 3.181093848e-01 lpclm = -6.559293371e-08 wpclm = 1.713416613e-07 ppclm = 2.209970241e-14
+ pdiblc1 = 1.655540522e+00 lpdiblc1 = -1.978548786e-07 wpdiblc1 = -4.945248368e-07 ppdiblc1 = 6.666166141e-14
+ pdiblc2 = 1.089453506e-01 lpdiblc2 = -2.930218689e-08 wpdiblc2 = -3.445059192e-08 ppdiblc2 = 9.872551410e-15
+ pdiblcb = 1.056061329e+01 lpdiblcb = -3.397750808e-06 wpdiblcb = -3.633910399e-06 ppdiblcb = 1.144776998e-12
+ drout = -6.895420402e+00 ldrout = 1.881719966e-06 wdrout = 2.659502130e-06 pdrout = -6.339928545e-13
+ pscbe1 = 7.996406531e+08 lpscbe1 = 1.066165136e-01 wpscbe1 = 1.104756920e-01 ppscbe1 = -3.592144900e-8
+ pscbe2 = 5.532468244e-08 lpscbe2 = -1.473278623e-14 wpscbe2 = -1.550083788e-14 ppscbe2 = 4.963799802e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.562104045e+01 lbeta0 = -2.219807606e-06 wbeta0 = -2.202063552e-06 pbeta0 = 7.479020182e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -2.165997771e-08 lagidl = 4.140862167e-15 wagidl = 8.283649030e-15 pagidl = -1.395147563e-21
+ bgidl = 5.034712953e+09 lbgidl = -9.609475445e+02 wbgidl = -1.359383558e+03 pbgidl = 3.237643686e-4
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 3.590081408e-01 lkt1 = -2.557098949e-07 wkt1 = -3.032729735e-07 pkt1 = 8.615428921e-14
+ kt2 = -1.085007458e-01 lkt2 = 8.093319375e-09 wkt2 = 2.229336925e-08 pkt2 = -2.726817351e-15
+ at = 6.062589996e+05 lat = -1.980565493e-01 wat = -1.688713709e-01 pat = 6.672960871e-8
+ ute = -6.536218925e+00 lute = 1.402703511e-06 wute = 2.058993995e-06 pute = -4.726016724e-13
+ ua1 = -4.119930358e-10 lua1 = 2.193614819e-16 wua1 = 2.376388479e-16 pua1 = -7.390770922e-23
+ ub1 = -1.516341639e-18 lub1 = 2.213870663e-25 wub1 = 5.292760388e-25 pub1 = -7.459017317e-32
+ uc1 = -1.097477057e-09 luc1 = 2.738227002e-16 wuc1 = 3.501098201e-16 puc1 = -9.225689179e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.188 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 4.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -3.7585e-8
+ vth0 = {1.339839766e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -5.927276991e-07 wvth0 = -7.883630360e-07 pvth0 = 1.957177521e-13
+ k1 = 4.972229255e+00 lk1 = -8.376433001e-07 wk1 = -1.692705614e-06 pk1 = 3.598915864e-13
+ k2 = -7.144369606e-02 lk2 = -7.628644380e-08 wk2 = 1.087479801e-07 pk2 = -6.929193578e-15
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.965541803e-02 ldsub = -5.773367104e-08 wdsub = 6.596370753e-07 pdsub = -9.363228619e-14
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {4.705032907e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.252178424e-06 wvoff = -1.599819475e-06 pvoff = 4.178657834e-13
+ nfactor = {-7.540355062e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.807409008e-05 wnfactor = 2.986168065e-05 pnfactor = -6.979964037e-12
+ eta0 = 8.685316948e+00 leta0 = -2.091199025e-06 weta0 = -2.761182577e-06 peta0 = 7.045709579e-13
+ etab = 4.487043903e-01 letab = -1.153189633e-07 wetab = -1.496157764e-07 petab = 3.845422872e-14
+ u0 = 3.638856988e-02 lu0 = -7.458932472e-09 wu0 = -1.538424624e-08 pu0 = 3.455480317e-15
+ ua = 3.728320601e-08 lua = -9.284595155e-15 wua = -1.585069750e-14 pua = 3.750933137e-21
+ ub = -5.587170849e-17 lub = 1.373891287e-23 wub = 2.231531575e-23 pub = -5.350001577e-30
+ uc = -8.098373510e-10 luc = 1.935074781e-16 wuc = 3.220466398e-16 puc = -7.772773327e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -9.099999229e+06 lvsat = 2.249533763e+00 wvsat = 3.366255253e+00 pvsat = -8.172625422e-7
+ a0 = -7.209609720e+00 la0 = 1.856310871e-06 wa0 = 3.230027234e-06 pa0 = -7.295397812e-13
+ ags = 1.250000289e+00 lags = -6.554234844e-14 wags = -9.753430241e-14 pags = 2.208265926e-20
+ a1 = 0.0
+ a2 = 8.598455755e-03 la2 = 4.010571531e-07 wa2 = -3.097467835e-07 pa2 = -1.792396435e-14
+ b0 = 4.160560674e-06 lb0 = -1.061650253e-12 wb0 = -1.401784424e-12 pb0 = 3.576933266e-19
+ b1 = 1.522909052e-20 lb1 = -3.429134306e-27 wb1 = -5.131015635e-27 pb1 = 1.155350789e-33
+ keta = -1.170107609e+00 lketa = 3.065938067e-07 wketa = 3.569566172e-07 pketa = -9.621190696e-14
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -4.252953167e+00 lpclm = 1.096123232e-06 wpclm = 2.222478178e-06 ppclm = -4.997113791e-13
+ pdiblc1 = 5.555095881e+00 lpdiblc1 = -1.207026823e-06 wpdiblc1 = -1.746357660e-06 ppdiblc1 = 3.908499914e-13
+ pdiblc2 = -1.049188729e-01 lpdiblc2 = 2.317802763e-08 wpdiblc2 = 4.516258627e-08 ppdiblc2 = -9.737664368e-15
+ pdiblcb = -3.931263837e+01 lpdiblcb = 9.085883561e-06 wpdiblcb = 1.388071711e-05 ppdiblcb = -3.242719083e-12
+ drout = 1.045272477e+00 ldrout = -1.019400399e-08 wdrout = -2.068588858e-08 pdrout = 4.657841654e-15
+ pscbe1 = 1.318130850e+09 lpscbe1 = -1.321889171e+02 wpscbe1 = -1.746587227e+02 ppscbe1 = 4.455737091e-5
+ pscbe2 = -1.189360255e-07 lpscbe2 = 2.868172788e-14 wpscbe2 = 4.282144700e-14 ppscbe2 = -9.563993577e-21
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 1.154054742e+00 lbeta0 = 1.313288627e-06 wbeta0 = 4.450616788e-06 pbeta0 = -8.962789824e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 5.088526994e-08 lagidl = -1.407494392e-14 wagidl = -1.922683959e-14 pagidl = 5.525121551e-21
+ bgidl = 1.000001405e+09 lbgidl = -3.160658941e-04 wbgidl = -4.733031311e-04 pbgidl = 1.064895535e-10
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -2.8385e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -8.126851427e-01 lkt1 = 2.501912487e-08 wkt1 = 4.349918723e-08 pkt1 = 3.817922281e-15
+ kt2 = 9.257212280e-01 lkt2 = -2.552314201e-07 wkt2 = -3.098630233e-07 pkt2 = 8.183489569e-14
+ at = -2.695540674e+06 lat = 6.303268747e-01 wat = 1.115261984e+00 pat = -2.561797010e-7
+ ute = -4.275804516e+00 lute = 9.260351592e-07 wute = 6.352886048e-07 pute = -1.430479352e-13
+ ua1 = 6.908188662e-10 lua1 = -4.638553775e-17 wua1 = -1.525939327e-15 pua1 = 3.708291796e-22
+ ub1 = 2.150944155e-19 lub1 = -2.046213969e-25 wub1 = 1.675794755e-24 pub1 = -3.724714206e-31
+ uc1 = -4.745326686e-11 luc1 = 2.543293342e-17 wuc1 = 5.817357230e-17 puc1 = -2.434859381e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.189 pmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 3.6e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.143603+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.43165561
+ k2 = 0.046387026
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 3.2465718e-7
+ voff = {-0.16725342+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {1.5720692+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.00827017
+ ua = -7.4124916e-10
+ ub = 6.3364395e-19
+ uc = -1.0566299e-10
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.464
+ ags = 0.11329
+ a1 = 0.0
+ a2 = 0.97
+ b0 = 5.7286e-9
+ b1 = 3.5674e-8
+ keta = 0.023361259
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.015
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0012771588
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0060625e-8
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.9002574e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.43825
+ kt2 = -0.058546
+ at = 70990.0
+ ute = -0.08298
+ ua1 = 2.0902e-9
+ ub1 = -1.2289e-18
+ uc1 = -2.9789e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.190 pmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 3.6e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.110002446e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -6.739656314e-7
+ k1 = 4.317683169e-01 lk1 = -2.260694917e-9
+ k2 = 5.812272789e-02 lk2 = -2.353967036e-7
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = -6.172472591e-06 lcit = 1.303205335e-10 wcit = -7.411538288e-28 pcit = -8.470329473e-33
+ voff = {-1.366450992e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -6.139469022e-7
+ nfactor = {1.491879866e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.608451299e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 5.757343843e-03 lu0 = 5.040269424e-8
+ ua = -6.997051773e-10 lua = -8.332962681e-16
+ ub = 2.914572873e-20 lub = 1.212512809e-23 pub = 1.540743956e-45
+ uc = -1.028126272e-10 luc = -5.717306066e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80156.0
+ a0 = 1.509528661e+00 la0 = -9.132216122e-07 wa0 = -4.440892099e-22
+ ags = 1.049766546e-01 lags = 1.667504950e-7
+ a1 = 0.0
+ a2 = 0.97
+ b0 = 1.603303665e-07 lb0 = -3.101028514e-12 wb0 = 9.926167351e-30 pb0 = 7.940933881e-35
+ b1 = -3.449654436e-08 lb1 = 1.407492708e-12 pb1 = -2.117582368e-34
+ keta = 2.267484931e-02 lketa = 1.376812233e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 1.338679197e-02 lpclm = 3.235800090e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 6.203397145e-05 lpdiblc2 = 2.437318038e-8
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 8.939788911e+08 lpscbe1 = -1.885044574e+3
+ pscbe2 = 1.029721146e-08 lpscbe2 = -4.745491455e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.672581664e-09 lagidl = -1.549141138e-14
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.927280546e-01 lkt1 = -9.130869187e-7
+ kt2 = -6.278728348e-02 lkt2 = 8.507238499e-8
+ at = 1.119456490e+05 lat = -8.214953706e-1
+ ute = 5.569192797e-01 lute = -1.283520854e-05 wute = -2.775557562e-23 pute = -8.881784197e-28
+ ua1 = 3.167657911e-09 lua1 = -2.161183394e-14
+ ub1 = -1.871357749e-18 lub1 = 1.288652674e-23
+ uc1 = -8.480682719e-11 luc1 = 1.103556931e-15
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.191 pmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 3.6e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.187828701e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -4.682843881e-8
+ k1 = 4.413127923e-01 lk1 = -7.917170021e-8
+ k2 = 2.360962024e-02 lk2 = 4.271578513e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.56
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.255222878e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.022405926e-7
+ nfactor = {1.474878960e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.745447485e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.082027174e-02 lu0 = 9.604760513e-9
+ ua = -6.138285144e-10 lua = -1.525305016e-15
+ ub = 9.744468811e-19 lub = 4.507730700e-24
+ uc = -1.127388117e-10 luc = 2.281382126e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.058684900e+05 lvsat = -2.071956159e-01 wvsat = -2.910383046e-17
+ a0 = 1.534954108e+00 la0 = -1.118104190e-6
+ ags = 5.727221290e-02 lags = 5.511609961e-7
+ a1 = 0.0
+ a2 = 1.142472225e+00 la2 = -1.389810509e-6
+ b0 = -2.847333882e-07 lb0 = 4.853708820e-13
+ b1 = 2.723349587e-07 lb1 = -1.065007706e-12
+ keta = 3.527851856e-02 lketa = -8.779438710e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -3.129792676e-01 lpclm = 2.662271191e-06 wpclm = 1.387778781e-23 ppclm = -4.163336342e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 5.631304475e-03 lpdiblc2 = -2.050494811e-08 ppdiblc2 = 6.938893904e-30
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 5.180633267e+08 lpscbe1 = 1.144146950e+3
+ pscbe2 = 9.867292200e-09 lpscbe2 = -1.281128963e-15
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 0.0
+ alpha1 = 0.0
+ beta0 = 30.0
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.567541838e-11 lagidl = 5.918390819e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.951066861e-01 lkt1 = 7.177144977e-7
+ kt2 = -4.582214957e-02 lkt2 = -5.163554810e-8
+ at = -5.187694708e+04 lat = 4.986149586e-01 wat = -7.275957614e-18
+ ute = -1.962096139e+00 lute = 7.463445942e-6
+ ua1 = -1.142173732e-09 lua1 = 1.311752211e-14 pua1 = -8.271806126e-37
+ ub1 = 5.970189960e-19 lub1 = -7.004072692e-24 wub1 = -9.629649722e-41 pub1 = 3.851859889e-46
+ uc1 = 1.352644816e-10 luc1 = -6.698150873e-16 puc1 = -1.033975766e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.192 pmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 3.6e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.240739996e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.678945911e-7
+ k1 = 3.703152982e-01 lk1 = 2.089482007e-7
+ k2 = 3.523254492e-02 lk2 = -4.452019127e-9
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 8.687255000e-01 ldsub = -1.252860562e-6
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.574246050e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 2.317056194e-7
+ nfactor = {1.804504494e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 4.077710329e-7
+ eta0 = 1.618122575e-01 leta0 = -3.320080490e-7
+ etab = -1.415214075e-01 letab = 2.902460303e-7
+ u0 = 1.876386465e-02 lu0 = -2.263168990e-8
+ ua = -1.142666133e-09 lua = 6.208079441e-16
+ ub = 3.578993877e-18 lub = -6.061963785e-24
+ uc = -1.462839997e-10 luc = 1.589458967e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.907739155e+04 lvsat = -1.730938371e-2
+ a0 = 1.290066750e+00 la0 = -1.243096602e-7
+ ags = 1.038557390e-01 lags = 3.621171281e-7
+ a1 = 0.0
+ a2 = 0.8
+ b0 = -2.443983594e-07 lb0 = 3.216844780e-13
+ b1 = 2.282768904e-08 lb1 = -5.246478891e-14
+ keta = 2.878940321e-02 lketa = -6.146045387e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 4.276671144e-02 lpclm = 1.218593531e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 7.314148344e-04 lpdiblc2 = -6.203629698e-10
+ pdiblcb = -0.225
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 9.730105367e-09 lpscbe2 = -7.244014714e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.029085000e-10 lalpha0 = 4.176201874e-16
+ alpha1 = -1.029085000e-10 lalpha1 = 4.176201874e-16
+ beta0 = 5.612050499e+01 lbeta0 = -1.060014497e-4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 9.753759806e-10 lagidl = 2.023762789e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.970340779e-01 lkt1 = -4.919148188e-7
+ kt2 = -6.504570086e-02 lkt2 = 2.637689104e-8
+ at = 1.337538942e+05 lat = -2.547065523e-1
+ ute = 8.473648282e-01 lute = -3.937824271e-06 wute = 5.551115123e-23 pute = -2.220446049e-28
+ ua1 = 3.772260014e-09 lua1 = -6.826085488e-15
+ ub1 = -2.010547992e-18 lub1 = 3.577877432e-24
+ uc1 = -1.141029631e-10 luc1 = 3.421603958e-16 wuc1 = 1.292469707e-32 puc1 = -2.584939414e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.193 pmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 3.6e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.157467255e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = -3.494866099e-9
+ k1 = 4.624286616e-01 lk1 = 1.936323952e-8
+ k2 = 3.323626527e-02 lk2 = -3.433362379e-10
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -5.230458000e-01 ldsub = 1.611641374e-06 pdsub = -1.110223025e-28
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.375103659e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -1.509827019e-8
+ nfactor = {3.873493641e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -3.850560359e-6
+ eta0 = -2.317683150e-01 leta0 = 4.780476779e-07 weta0 = 2.818925648e-24 peta0 = -4.878909776e-29
+ etab = 8.945695385e-01 letab = -1.842205272e-06 wetab = 5.269222558e-23 petab = 4.878909776e-29
+ u0 = 8.869023499e-03 lu0 = -2.266424694e-9
+ ua = -7.069494059e-10 lua = -2.759711530e-16
+ ub = 5.978104287e-19 lub = 7.381855434e-26
+ uc = -8.501444316e-11 luc = 3.284273356e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.150316568e+04 lvsat = -2.230203925e-2
+ a0 = 1.335558190e+00 la0 = -2.179387784e-07 wa0 = 4.440892099e-22
+ ags = -2.740734130e-01 lags = 1.139959571e-06 pags = -1.110223025e-28
+ a1 = 0.0
+ a2 = 0.8
+ b0 = -2.445519084e-08 lb0 = -1.309959532e-13
+ b1 = -1.081702893e-08 lb1 = 1.678176028e-14
+ keta = 1.248468452e-02 lketa = -2.790257100e-08 wketa = -8.673617380e-25 pketa = -2.168404345e-30
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 8.813067537e-01 lpclm = -5.072644274e-7
+ pdiblc1 = 3.914291538e-01 lpdiblc1 = -2.941441518e-9
+ pdiblc2 = 0.00043
+ pdiblcb = -0.225
+ drout = 2.586727596e-01 ldrout = 6.201826865e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 9.677303407e-09 lpscbe2 = -6.157260625e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.244501660e-10 lalpha0 = -5.032259808e-17
+ alpha1 = 3.116340000e-10 lalpha1 = -4.355787498e-16
+ beta0 = 2.879161404e+00 lbeta0 = 3.578286399e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.873878404e-09 lagidl = -1.883677944e-15 wagidl = 8.271806126e-31
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -6.132969917e-01 lkt1 = 1.590080226e-7
+ kt2 = -5.312415365e-02 lkt2 = 1.840320218e-9
+ at = -2.149431371e+04 lat = 6.482065165e-02 wat = -3.637978807e-18
+ ute = -1.125474971e+00 lute = 1.226154181e-7
+ ua1 = 1.581139030e-09 lua1 = -2.316386012e-15 wua1 = -2.067951531e-31
+ ub1 = -1.786167891e-18 lub1 = 3.116065039e-24 pub1 = -1.925929944e-46
+ uc1 = -6.034070260e-12 luc1 = 1.197362425e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.194 pmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 3.6e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.179585911e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 1.991043223e-8
+ k1 = 4.590636320e-01 lk1 = 2.292401288e-8
+ k2 = 4.879497130e-02 lk2 = -1.680709220e-8
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 1.826091600e+00 ldsub = -8.741453484e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-1.514115416e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = -3.884631052e-10
+ nfactor = {-2.848701323e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 5.496954346e-7
+ eta0 = -8.141180000e-02 leta0 = 3.189449244e-7
+ etab = -1.791190270e+00 letab = 9.997851843e-7
+ u0 = 8.511814296e-03 lu0 = -1.888436632e-9
+ ua = -5.676393665e-10 lua = -4.233848574e-16
+ ub = 4.558630568e-19 lub = 2.240230049e-25
+ uc = -9.465257987e-11 luc = 4.304152068e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.812294335e+04 lvsat = 7.253762053e-2
+ a0 = 1.450327954e+00 la0 = -3.393846989e-7
+ ags = 3.044616148e-01 lags = 5.277711605e-7
+ a1 = 0.0
+ a2 = 6.102222000e-01 la2 = 2.008171746e-7
+ b0 = -2.291120879e-07 lb0 = 8.556583555e-14
+ b1 = 7.802908820e-09 lb1 = -2.921299252e-15
+ keta = 3.180813056e-03 lketa = -1.805749334e-8
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 8.071632109e-01 lpclm = -4.288079548e-7
+ pdiblc1 = 8.079624086e-01 lpdiblc1 = -4.437044358e-7
+ pdiblc2 = 8.800245625e-04 lpdiblc2 = -4.762024913e-10
+ pdiblcb = -3.644375305e-01 lpdiblcb = 1.475486117e-7
+ drout = 6.714648809e-01 ldrout = 1.833784474e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 9.036653136e-09 lpscbe2 = 6.219083455e-17
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 5.109966807e-11 lalpha0 = 2.729469827e-17
+ alpha1 = -3.232680000e-10 lalpha1 = 2.362554996e-16
+ beta0 = 4.133699773e+00 lbeta0 = 2.250771533e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 1.198830479e-09 lagidl = -1.111924814e-16 wagidl = 4.135903063e-31
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.174275110e-01 lkt1 = -4.825518579e-8
+ kt2 = -4.227678194e-02 lkt2 = -9.638043105e-9
+ at = -5.155172580e+03 lat = 4.753106268e-2
+ ute = -1.948441940e+00 lute = 9.934543756e-07 wute = 4.440892099e-22
+ ua1 = -2.762234095e-09 lua1 = 2.279641128e-15 wua1 = -4.135903063e-31
+ ub1 = 3.342842007e-18 lub1 = -2.311299365e-24
+ uc1 = 3.018867235e-10 luc1 = -2.060963038e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.195 pmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 3.6e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.264103765e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 6.708576316e-8
+ k1 = 6.683388805e-02 lk1 = 2.418548891e-7
+ k2 = 1.997888937e-01 lk2 = -1.010873698e-07 wk2 = 2.775557562e-23 pk2 = -3.469446952e-30
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = -2.357046223e-01 ldsub = 2.766874491e-7
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-2.285774571e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 4.268323597e-8
+ nfactor = {-1.975544531e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = 1.493379164e-06 pnfactor = -2.220446049e-28
+ eta0 = 0.49
+ etab = -6.25e-6
+ u0 = 9.368291226e-03 lu0 = -2.366496360e-9
+ ua = 1.439815915e-10 lua = -8.205903276e-16
+ ub = -5.195069026e-19 lub = 7.684452551e-25
+ uc = -3.948092127e-11 luc = 1.224635600e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.030911662e+04 lvsat = 6.817617687e-2
+ a0 = 4.428862462e-01 la0 = 2.229390391e-7
+ ags = 1.25
+ a1 = 0.0
+ a2 = 1.607916892e+00 la2 = -3.560660718e-7
+ b0 = -1.692706342e-07 lb0 = 5.216413134e-14
+ b1 = 5.736201456e-09 lb1 = -1.767725203e-15
+ keta = -3.034356046e-02 lketa = 6.548062299e-10
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = -9.321010719e-01 lpclm = 5.419971900e-07 wpclm = -8.326672685e-23 ppclm = 6.938893904e-30
+ pdiblc1 = -2.023541524e-01 lpdiblc1 = 1.202239591e-07 wpdiblc1 = -2.775557562e-23 ppdiblc1 = 3.469446952e-30
+ pdiblc2 = -8.192060195e-03 lpdiblc2 = 4.587563058e-09 wpdiblc2 = 5.014435048e-25 ppdiblc2 = -3.625301014e-31
+ pdiblcb = 5.387506110e-02 lpdiblcb = -8.594092758e-8
+ drout = 1.002336791e+00 ldrout = -1.304326898e-9
+ pscbe1 = 8.000387678e+08 lpscbe1 = -2.163901511e-2
+ pscbe2 = 8.939243981e-09 lpscbe2 = 1.165617027e-16
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 7.033152730e+00 lbeta0 = 6.323838756e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.375324279e-09 lagidl = 1.325623480e-15
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.579749968e-01 lkt1 = -2.562279564e-8
+ kt2 = -8.075965548e-02 lkt2 = 1.184194242e-08 wkt2 = -2.775557562e-23
+ at = 4.913246012e+04 lat = 1.722933473e-2
+ ute = 1.474961324e-01 lute = -1.764353782e-7
+ ua1 = 2.589797668e-09 lua1 = -7.077024411e-16
+ ub1 = -1.848973245e-18 lub1 = 5.866161545e-25 pub1 = 9.629649722e-47
+ uc1 = -7.846037752e-11 luc1 = 6.202037590e-18
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.196 pmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.6e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -2.9085e-8
+ vth0 = {-1.046413+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))}
+ k1 = 0.85164386
+ k2 = -0.1282358
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 0.66213569
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-0.09007197+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))}
+ nfactor = {2.8704144+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))}
+ eta0 = 0.49
+ etab = -6.25e-6
+ u0 = 0.0016891
+ ua = -2.518803e-9
+ ub = 1.9740689e-18
+ uc = 2.58041e-13
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 200920.0
+ a0 = 1.166315
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.45249595
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.028218739
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 0.82665932
+ pdiblc1 = 0.18776805
+ pdiblc2 = 0.0066944085
+ pdiblcb = -0.225
+ drout = 0.9981043
+ pscbe1 = 799968550.0
+ pscbe2 = 9.3174823e-9
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 9.0852145
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 2.9262738e-9
+ bgidl = 1000000000.0
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -1.9885e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.54112
+ kt2 = -0.042333
+ at = 105041.0
+ ute = -0.42503
+ ua1 = 2.9333e-10
+ ub1 = 5.4574e-20
+ uc1 = -5.8335e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__pfet_01v8_hvt__model.197 pmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.6e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.44996e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-9*1.052*(sky130_fd_pr__pfet_01v8_hvt__toxe_slope/sqrt(l*w*mult)))}
+ toxm = 4.23e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 4.1539e-8
+ lint = -3.7585e-8
+ vth0 = {-4.263958532e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__vth0_slope/sqrt(l*w*mult))} lvth0 = 8.210210934e-07 wvth0 = 1.099679894e-06 pvth0 = -2.806053186e-13
+ k1 = -1.998450892e+00 lk1 = 7.272586779e-07 wk1 = 6.558698822e-07 pk1 = -1.673583179e-13
+ k2 = -1.169590294e+00 lk2 = 2.657224262e-07 wk2 = 4.787377281e-07 pk2 = -1.221595061e-13
+ k3 = -13.778
+ k3b = 2.0
+ w0 = 0.0
+ dvt0 = 4.05
+ dvt1 = 0.3
+ dvt2 = 0.03
+ dvt0w = -4.254
+ dvt1w = 1147200.0
+ dvt2w = -0.00896
+ dsub = 7.005387830e+00 ldsub = -1.618607649e-06 wdsub = -1.694009861e-06 pdsub = 4.322604961e-13
+ minv = 0.0
+ voffl = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ cit = 1.0e-5
+ voff = {-5.439247112e+00+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__voff_slope/sqrt(l*w*mult))} lvoff = 1.364949021e-06 wvoff = 1.818011638e-06 pvoff = -4.639020297e-13
+ nfactor = {6.788592669e+01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_hvt__nfactor_slope/sqrt(l*w*mult))} lnfactor = -1.659000827e-05 wnfactor = -1.841569662e-05 pnfactor = 4.699133307e-12
+ eta0 = 8.076559862e+00 leta0 = -1.935862480e-06 weta0 = -2.556078922e-06 peta0 = 6.522346585e-13
+ etab = 4.410669612e-01 letab = -1.125486513e-07 wetab = -1.470425585e-07 petab = 3.752084965e-14
+ u0 = 3.849175305e-02 lu0 = -9.390932978e-09 wu0 = -1.609285492e-08 pu0 = 4.106413791e-15
+ ua = -2.530694941e-08 lua = 5.814851319e-15 wua = 5.237302848e-15 pua = -1.336402568e-21
+ ub = 4.347944645e-17 lub = -1.059092719e-23 wub = -1.115827407e-23 pub = 2.847256795e-30
+ uc = -3.313787141e-10 luc = 8.462375079e-17 wuc = 1.608433990e-16 puc = -4.104241011e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.128553123e+06 lvsat = -7.470441441e-01 wvsat = -7.538130629e-01 pvsat = 1.923504793e-7
+ a0 = 2.172606755e+00 la0 = -2.567754672e-07 wa0 = 6.895209465e-08 pa0 = -1.759450599e-14
+ ags = 1.249999986e+00 lags = 3.698335860e-15 wags = 4.883215610e-15 pags = -1.246050818e-21
+ a1 = 0.0
+ a2 = -8.940045776e+00 la2 = 2.396694872e-06 wa2 = 2.705248328e-06 pa2 = -6.902982160e-13
+ b0 = 0.0
+ b1 = 3.029193301e-28 lb1 = -7.729592547e-35 wb1 = -1.020601866e-34 pb1 = 2.604269780e-41
+ keta = -1.560996587e+00 lketa = 3.911189234e-07 wketa = 4.886557132e-07 pketa = -1.246902783e-13
+ dwg = -5.722e-9
+ dwb = -1.7864e-8
+ pclm = 2.409775491e+00 lpclm = -4.039637534e-07 wpclm = -2.234168728e-08 ppclm = 5.700928344e-15
+ pdiblc1 = 1.540931479e-01 lpdiblc1 = 8.592824768e-09 wpdiblc1 = 7.335898328e-08 ppdiblc1 = -1.871901176e-14
+ pdiblc2 = 6.865378525e-02 lpdiblc2 = -1.581017416e-08 wpdiblc2 = -1.331786087e-08 ppdiblc2 = 3.398318559e-15
+ pdiblcb = -8.847714611e+00 lpdiblcb = 2.200258087e-06 wpdiblcb = 3.616414065e-06 ppdiblcb = -9.228003771e-13
+ drout = 9.838757930e-01 ldrout = 3.630688140e-09 wdrout = 4.964615385e-15 pdrout = -1.266820870e-21
+ pscbe1 = 1.278681003e+09 lpscbe1 = -1.221530566e+02 wpscbe1 = -1.613672012e+02 ppscbe1 = 4.117606873e-5
+ pscbe2 = 1.531392544e-08 lpscbe2 = -1.530112395e-15 wpscbe2 = -2.410314978e-15 ppscbe2 = 6.150400730e-22
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 531.92
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = -0.32348
+ prwg = 0.02
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.0e-10
+ alpha1 = 1.0e-10
+ beta0 = 2.405955718e+01 lbeta0 = -3.821003023e-06 wbeta0 = -3.266750906e-06 pbeta0 = 8.335768286e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = -1.495839366e-07 lagidl = 3.891603038e-14 wagidl = 4.831564640e-14 pagidl = -1.232870349e-20
+ bgidl = 1.000000010e+09 lbgidl = -2.573869705e-06 wbgidl = -3.398494720e-06 pbgidl = 8.671936989e-13
+ cgidl = 300.0
+ egidl = 0.1
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.23e-9
+ dlcig = 0.0
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 1.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = -2.8385e-8
+ dwc = 3.2175e-8
+ xpart = 0.0
+ cgso = 7.2e-11
+ cgdo = 7.2e-11
+ cgbo = 0.0
+ cgdl = 9.12e-12
+ cgsl = 9.12e-12
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.2e-11
+ ckappas = 0.6
+ vfbcv = -0.1446893
+ acde = 0.552
+ moin = 14.504
+ noff = 4.0
+ voffcv = -0.1375
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.88
+ noia = 1.2e+41
+ noib = 2.0e+25
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -6.0e-8
+ af = 1.0
+ kf = 0.0
+ tnoia = 1.5
+ tnoib = 3.5
+ rnoia = 0.577
+ rnoib = 0.37
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 2.17e-5
+ jsws = 8.2e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 12.8
+ xjbvs = 1.0
+ pbs = 0.6587
+ cjs = 0.000813867531
+ mjs = 0.34629
+ pbsws = 0.7418
+ cjsws = 1.041095405e-10
+ mjsws = 0.26859
+ pbswgs = 1.3925
+ cjswgs = 2.78207363e-10
+ mjswgs = 0.70393
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 5.631474861e-01 lkt1 = -2.817759344e-07 wkt1 = -4.200490937e-07 pkt1 = 1.071839272e-13
+ kt2 = 1.110837488e+00 lkt2 = -2.942545135e-07 wkt2 = -3.722327639e-07 pkt2 = 9.498263437e-14
+ at = 1.515353355e+05 lat = -1.186395958e-02 wat = 1.560194409e-01 pat = -3.981148075e-8
+ ute = -2.390238694e+00 lute = 5.014623024e-07 wute = -3.199576604e-15 pute = 8.164360299e-22
+ ua1 = -1.344042497e-09 lua1 = 4.178083401e-16 wua1 = -8.403497662e-16 pua1 = 2.144320498e-22
+ ub1 = 5.634704891e-18 lub1 = -1.423881999e-24 wub1 = -1.501912456e-25 pub1 = 3.832430013e-32
+ uc1 = -9.051005315e-10 luc1 = 2.160691607e-16 wuc1 = 3.471338040e-16 puc1 = -8.857813276e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2556
+ tpb = 0.0019551
+ tcj = 0.0012407
+ tpbsw = 0.00014242
+ tcjsw = 0.0
+ tpbswg = 0.0
+ tcjswg = 2.0e-12
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 2.65e-8
+ lkvth0 = 0.0
+ wkvth0 = 2.5e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = 4.5e-8
+ lku0 = 0.0
+ wku0 = 2.5e-7
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.4
+ steta0 = 0.0
.ends sky130_fd_pr__pfet_01v8_hvt
* Well Proximity Effect Parameters
